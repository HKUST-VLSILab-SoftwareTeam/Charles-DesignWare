SITE  IOSite
    CLASS       PAD ;
    SYMMETRY    Y ;
    SIZE        0.005 BY 174.000 ;
END  IOSite

SITE  CornerSite
    CLASS	PAD ;
    SYMMETRY	R90 Y ;
    SIZE	174.000 BY 174.000 ;
END  CornerSite

MACRO PLVSSO
  CLASS  PAD ;
  FOREIGN PLVSSO 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN VSSO
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V6 ;
        RECT 4.310 173.515 4.670 173.875 ;
        RECT 5.020 173.515 5.380 173.875 ;
        RECT 5.730 173.515 6.090 173.875 ;
        RECT 6.440 173.515 6.800 173.875 ;
        RECT 7.150 173.515 7.510 173.875 ;
        RECT 7.860 173.515 8.220 173.875 ;
        RECT 8.570 173.515 8.930 173.875 ;
        RECT 9.280 173.515 9.640 173.875 ;
        RECT 9.990 173.515 10.350 173.875 ;
        RECT 10.700 173.515 11.060 173.875 ;
        RECT 11.410 173.515 11.770 173.875 ;
        RECT 12.120 173.515 12.480 173.875 ;
        RECT 12.830 173.515 13.190 173.875 ;
        RECT 13.540 173.515 13.900 173.875 ;
        RECT 14.250 173.515 14.610 173.875 ;
        RECT 14.960 173.515 15.320 173.875 ;
        RECT 15.670 173.515 16.030 173.875 ;
        RECT 16.380 173.515 16.740 173.875 ;
        RECT 17.090 173.515 17.450 173.875 ;
        RECT 17.800 173.515 18.160 173.875 ;
        RECT 18.510 173.515 18.870 173.875 ;
        RECT 19.220 173.515 19.580 173.875 ;
        RECT 19.930 173.515 20.290 173.875 ;
        RECT 20.640 173.515 21.000 173.875 ;
        RECT 21.350 173.515 21.710 173.875 ;
        RECT 22.060 173.515 22.420 173.875 ;
        RECT 22.770 173.515 23.130 173.875 ;
        RECT 23.480 173.515 23.840 173.875 ;
        RECT 24.190 173.515 24.550 173.875 ;
        RECT 24.900 173.515 25.260 173.875 ;
        RECT 25.610 173.515 25.970 173.875 ;
        RECT 26.320 173.515 26.680 173.875 ;
        RECT 27.030 173.515 27.390 173.875 ;
        RECT 27.740 173.515 28.100 173.875 ;
        RECT 28.450 173.515 28.810 173.875 ;
        RECT 29.160 173.515 29.520 173.875 ;
        RECT 29.870 173.515 30.230 173.875 ;
        RECT 30.580 173.515 30.940 173.875 ;
        RECT 31.290 173.515 31.650 173.875 ;
        RECT 32.000 173.515 32.360 173.875 ;
        RECT 32.710 173.515 33.070 173.875 ;
        RECT 33.420 173.515 33.780 173.875 ;
        RECT 34.130 173.515 34.490 173.875 ;
        RECT 34.840 173.515 35.200 173.875 ;
        RECT 35.550 173.515 35.910 173.875 ;
        RECT 36.260 173.515 36.620 173.875 ;
        RECT 36.970 173.515 37.330 173.875 ;
        RECT 37.680 173.515 38.040 173.875 ;
        RECT 38.390 173.515 38.750 173.875 ;
        RECT 39.100 173.515 39.460 173.875 ;
        RECT 39.810 173.515 40.170 173.875 ;
        RECT 40.520 173.515 40.880 173.875 ;
        RECT 41.230 173.515 41.590 173.875 ;
        RECT 41.940 173.515 42.300 173.875 ;
        RECT 42.650 173.515 43.010 173.875 ;
        RECT 43.360 173.515 43.720 173.875 ;
        RECT 44.070 173.515 44.430 173.875 ;
        RECT 44.780 173.515 45.140 173.875 ;
        RECT 45.490 173.515 45.850 173.875 ;
        RECT 46.200 173.515 46.560 173.875 ;
        RECT 46.910 173.515 47.270 173.875 ;
        RECT 47.620 173.515 47.980 173.875 ;
        RECT 48.330 173.515 48.690 173.875 ;
        RECT 49.040 173.515 49.400 173.875 ;
        RECT 49.750 173.515 50.110 173.875 ;
        RECT 50.460 173.515 50.820 173.875 ;
        RECT 51.170 173.515 51.530 173.875 ;
        RECT 51.880 173.515 52.240 173.875 ;
        RECT 52.590 173.515 52.950 173.875 ;
        RECT 53.300 173.515 53.660 173.875 ;
        RECT 54.010 173.515 54.370 173.875 ;
        RECT 54.720 173.515 55.080 173.875 ;
        RECT 55.430 173.515 55.790 173.875 ;
        RECT 56.140 173.515 56.500 173.875 ;
        RECT 56.850 173.515 57.210 173.875 ;
        RECT 57.560 173.515 57.920 173.875 ;
        RECT 58.270 173.515 58.630 173.875 ;
        RECT 58.980 173.515 59.340 173.875 ;
        RECT 59.690 173.515 60.050 173.875 ;
        RECT 60.400 173.515 60.760 173.875 ;
        RECT 61.110 173.515 61.470 173.875 ;
        RECT 61.820 173.515 62.180 173.875 ;
        RECT 62.530 173.515 62.890 173.875 ;
        RECT 63.240 173.515 63.600 173.875 ;
        RECT 63.950 173.515 64.310 173.875 ;
        RECT 64.660 173.515 65.020 173.875 ;
        RECT 65.370 173.515 65.730 173.875 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V3 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.300 66.490 174.000 ;
      LAYER V2 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.300 66.490 174.000 ;
      LAYER V1 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M1 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V5 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V4 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
    END
  END VSSO
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.600 0.700 113.895 ;
        RECT 0.190 92.280 0.700 100.280 ;
        RECT 0.205 81.280 0.700 89.280 ;
        RECT 0.205 70.000 0.700 79.520 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 110.465 69.415 113.895 ;
        RECT 69.420 150.320 69.675 151.785 ;
        RECT 69.300 152.430 69.685 154.220 ;
        RECT 69.300 81.365 69.740 89.280 ;
        RECT 69.300 70.000 69.740 77.985 ;
        RECT 69.300 115.135 69.780 118.565 ;
        RECT 69.300 105.320 69.780 108.750 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 162.720 69.845 170.465 ;
        RECT 69.300 92.360 69.850 100.195 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 118.565 ;
        RECT 69.420 150.320 70.000 151.785 ;
        RECT 69.560 115.135 70.000 154.220 ;
        RECT 69.300 152.430 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.600 0.700 113.895 ;
        RECT 0.190 92.280 0.700 100.280 ;
        RECT 0.205 81.280 0.700 89.280 ;
        RECT 0.205 70.000 0.700 79.520 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 110.465 69.415 113.895 ;
        RECT 69.420 150.320 69.675 151.785 ;
        RECT 69.300 152.430 69.685 154.220 ;
        RECT 69.300 81.365 69.740 89.280 ;
        RECT 69.300 70.000 69.740 77.985 ;
        RECT 69.300 115.135 69.780 118.565 ;
        RECT 69.300 105.320 69.780 108.750 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 162.720 69.845 170.465 ;
        RECT 69.300 92.360 69.850 100.195 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.600 0.700 113.895 ;
        RECT 0.190 92.280 0.700 100.280 ;
        RECT 0.205 81.280 0.700 89.280 ;
        RECT 0.205 70.000 0.700 79.520 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 110.465 69.415 113.895 ;
        RECT 69.420 150.320 69.675 151.785 ;
        RECT 69.300 152.430 69.685 154.220 ;
        RECT 69.300 81.365 69.740 89.280 ;
        RECT 69.300 70.000 69.740 77.985 ;
        RECT 69.300 115.135 69.780 118.565 ;
        RECT 69.300 105.320 69.780 108.750 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 162.720 69.845 170.465 ;
        RECT 69.300 92.360 69.850 100.195 ;
  END 
END PLVSSO

MACRO PLVSSH
  CLASS  PAD ;
  FOREIGN PLVSSH 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN VSSH
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V6 ;
        RECT 4.310 173.515 4.670 173.875 ;
        RECT 5.020 173.515 5.380 173.875 ;
        RECT 5.730 173.515 6.090 173.875 ;
        RECT 6.440 173.515 6.800 173.875 ;
        RECT 7.150 173.515 7.510 173.875 ;
        RECT 7.860 173.515 8.220 173.875 ;
        RECT 8.570 173.515 8.930 173.875 ;
        RECT 9.280 173.515 9.640 173.875 ;
        RECT 9.990 173.515 10.350 173.875 ;
        RECT 10.700 173.515 11.060 173.875 ;
        RECT 11.410 173.515 11.770 173.875 ;
        RECT 12.120 173.515 12.480 173.875 ;
        RECT 12.830 173.515 13.190 173.875 ;
        RECT 13.540 173.515 13.900 173.875 ;
        RECT 14.250 173.515 14.610 173.875 ;
        RECT 14.960 173.515 15.320 173.875 ;
        RECT 15.670 173.515 16.030 173.875 ;
        RECT 16.380 173.515 16.740 173.875 ;
        RECT 17.090 173.515 17.450 173.875 ;
        RECT 17.800 173.515 18.160 173.875 ;
        RECT 18.510 173.515 18.870 173.875 ;
        RECT 19.220 173.515 19.580 173.875 ;
        RECT 19.930 173.515 20.290 173.875 ;
        RECT 20.640 173.515 21.000 173.875 ;
        RECT 21.350 173.515 21.710 173.875 ;
        RECT 22.060 173.515 22.420 173.875 ;
        RECT 22.770 173.515 23.130 173.875 ;
        RECT 23.480 173.515 23.840 173.875 ;
        RECT 24.190 173.515 24.550 173.875 ;
        RECT 24.900 173.515 25.260 173.875 ;
        RECT 25.610 173.515 25.970 173.875 ;
        RECT 26.320 173.515 26.680 173.875 ;
        RECT 27.030 173.515 27.390 173.875 ;
        RECT 27.740 173.515 28.100 173.875 ;
        RECT 28.450 173.515 28.810 173.875 ;
        RECT 29.160 173.515 29.520 173.875 ;
        RECT 29.870 173.515 30.230 173.875 ;
        RECT 30.580 173.515 30.940 173.875 ;
        RECT 31.290 173.515 31.650 173.875 ;
        RECT 32.000 173.515 32.360 173.875 ;
        RECT 32.710 173.515 33.070 173.875 ;
        RECT 33.420 173.515 33.780 173.875 ;
        RECT 34.130 173.515 34.490 173.875 ;
        RECT 34.840 173.515 35.200 173.875 ;
        RECT 35.550 173.515 35.910 173.875 ;
        RECT 36.260 173.515 36.620 173.875 ;
        RECT 36.970 173.515 37.330 173.875 ;
        RECT 37.680 173.515 38.040 173.875 ;
        RECT 38.390 173.515 38.750 173.875 ;
        RECT 39.100 173.515 39.460 173.875 ;
        RECT 39.810 173.515 40.170 173.875 ;
        RECT 40.520 173.515 40.880 173.875 ;
        RECT 41.230 173.515 41.590 173.875 ;
        RECT 41.940 173.515 42.300 173.875 ;
        RECT 42.650 173.515 43.010 173.875 ;
        RECT 43.360 173.515 43.720 173.875 ;
        RECT 44.070 173.515 44.430 173.875 ;
        RECT 44.780 173.515 45.140 173.875 ;
        RECT 45.490 173.515 45.850 173.875 ;
        RECT 46.200 173.515 46.560 173.875 ;
        RECT 46.910 173.515 47.270 173.875 ;
        RECT 47.620 173.515 47.980 173.875 ;
        RECT 48.330 173.515 48.690 173.875 ;
        RECT 49.040 173.515 49.400 173.875 ;
        RECT 49.750 173.515 50.110 173.875 ;
        RECT 50.460 173.515 50.820 173.875 ;
        RECT 51.170 173.515 51.530 173.875 ;
        RECT 51.880 173.515 52.240 173.875 ;
        RECT 52.590 173.515 52.950 173.875 ;
        RECT 53.300 173.515 53.660 173.875 ;
        RECT 54.010 173.515 54.370 173.875 ;
        RECT 54.720 173.515 55.080 173.875 ;
        RECT 55.430 173.515 55.790 173.875 ;
        RECT 56.140 173.515 56.500 173.875 ;
        RECT 56.850 173.515 57.210 173.875 ;
        RECT 57.560 173.515 57.920 173.875 ;
        RECT 58.270 173.515 58.630 173.875 ;
        RECT 58.980 173.515 59.340 173.875 ;
        RECT 59.690 173.515 60.050 173.875 ;
        RECT 60.400 173.515 60.760 173.875 ;
        RECT 61.110 173.515 61.470 173.875 ;
        RECT 61.820 173.515 62.180 173.875 ;
        RECT 62.530 173.515 62.890 173.875 ;
        RECT 63.240 173.515 63.600 173.875 ;
        RECT 63.950 173.515 64.310 173.875 ;
        RECT 64.660 173.515 65.020 173.875 ;
        RECT 65.370 173.515 65.730 173.875 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V3 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.300 66.490 174.000 ;
      LAYER V2 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.300 66.490 174.000 ;
      LAYER V1 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M1 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V5 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V4 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
    END
  END VSSH
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.600 0.700 113.895 ;
        RECT 0.190 92.280 0.700 100.280 ;
        RECT 0.205 81.280 0.700 89.280 ;
        RECT 0.205 70.000 0.700 79.520 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 110.465 69.415 113.895 ;
        RECT 69.420 150.320 69.675 151.785 ;
        RECT 69.300 152.430 69.685 154.220 ;
        RECT 69.300 81.365 69.740 89.280 ;
        RECT 69.300 70.000 69.740 77.985 ;
        RECT 69.300 115.135 69.780 118.565 ;
        RECT 69.300 105.320 69.780 108.750 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 162.720 69.845 170.465 ;
        RECT 69.300 92.360 69.850 100.195 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 118.565 ;
        RECT 69.420 150.320 70.000 151.785 ;
        RECT 69.560 115.135 70.000 154.220 ;
        RECT 69.300 152.430 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.600 0.700 113.895 ;
        RECT 0.190 92.280 0.700 100.280 ;
        RECT 0.205 81.280 0.700 89.280 ;
        RECT 0.205 70.000 0.700 79.520 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 110.465 69.415 113.895 ;
        RECT 69.420 150.320 69.675 151.785 ;
        RECT 69.300 152.430 69.685 154.220 ;
        RECT 69.300 81.365 69.740 89.280 ;
        RECT 69.300 70.000 69.740 77.985 ;
        RECT 69.300 115.135 69.780 118.565 ;
        RECT 69.300 105.320 69.780 108.750 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 162.720 69.845 170.465 ;
        RECT 69.300 92.360 69.850 100.195 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.600 0.700 113.895 ;
        RECT 0.190 92.280 0.700 100.280 ;
        RECT 0.205 81.280 0.700 89.280 ;
        RECT 0.205 70.000 0.700 79.520 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 110.465 69.415 113.895 ;
        RECT 69.420 150.320 69.675 151.785 ;
        RECT 69.300 152.430 69.685 154.220 ;
        RECT 69.300 81.365 69.740 89.280 ;
        RECT 69.300 70.000 69.740 77.985 ;
        RECT 69.300 115.135 69.780 118.565 ;
        RECT 69.300 105.320 69.780 108.750 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 162.720 69.845 170.465 ;
        RECT 69.300 92.360 69.850 100.195 ;
  END 
END PLVSSH

MACRO PLVSSC
  CLASS  PAD ;
  FOREIGN PLVSSC 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    CLASS CORE ;
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V6 ;
        RECT 4.310 173.515 4.670 173.875 ;
        RECT 5.020 173.515 5.380 173.875 ;
        RECT 5.730 173.515 6.090 173.875 ;
        RECT 6.440 173.515 6.800 173.875 ;
        RECT 7.150 173.515 7.510 173.875 ;
        RECT 7.860 173.515 8.220 173.875 ;
        RECT 8.570 173.515 8.930 173.875 ;
        RECT 9.280 173.515 9.640 173.875 ;
        RECT 9.990 173.515 10.350 173.875 ;
        RECT 10.700 173.515 11.060 173.875 ;
        RECT 11.410 173.515 11.770 173.875 ;
        RECT 12.120 173.515 12.480 173.875 ;
        RECT 12.830 173.515 13.190 173.875 ;
        RECT 13.540 173.515 13.900 173.875 ;
        RECT 14.250 173.515 14.610 173.875 ;
        RECT 14.960 173.515 15.320 173.875 ;
        RECT 15.670 173.515 16.030 173.875 ;
        RECT 16.380 173.515 16.740 173.875 ;
        RECT 17.090 173.515 17.450 173.875 ;
        RECT 17.800 173.515 18.160 173.875 ;
        RECT 18.510 173.515 18.870 173.875 ;
        RECT 19.220 173.515 19.580 173.875 ;
        RECT 19.930 173.515 20.290 173.875 ;
        RECT 20.640 173.515 21.000 173.875 ;
        RECT 21.350 173.515 21.710 173.875 ;
        RECT 22.060 173.515 22.420 173.875 ;
        RECT 22.770 173.515 23.130 173.875 ;
        RECT 23.480 173.515 23.840 173.875 ;
        RECT 24.190 173.515 24.550 173.875 ;
        RECT 24.900 173.515 25.260 173.875 ;
        RECT 25.610 173.515 25.970 173.875 ;
        RECT 26.320 173.515 26.680 173.875 ;
        RECT 27.030 173.515 27.390 173.875 ;
        RECT 27.740 173.515 28.100 173.875 ;
        RECT 28.450 173.515 28.810 173.875 ;
        RECT 29.160 173.515 29.520 173.875 ;
        RECT 29.870 173.515 30.230 173.875 ;
        RECT 30.580 173.515 30.940 173.875 ;
        RECT 31.290 173.515 31.650 173.875 ;
        RECT 32.000 173.515 32.360 173.875 ;
        RECT 32.710 173.515 33.070 173.875 ;
        RECT 33.420 173.515 33.780 173.875 ;
        RECT 34.130 173.515 34.490 173.875 ;
        RECT 34.840 173.515 35.200 173.875 ;
        RECT 35.550 173.515 35.910 173.875 ;
        RECT 36.260 173.515 36.620 173.875 ;
        RECT 36.970 173.515 37.330 173.875 ;
        RECT 37.680 173.515 38.040 173.875 ;
        RECT 38.390 173.515 38.750 173.875 ;
        RECT 39.100 173.515 39.460 173.875 ;
        RECT 39.810 173.515 40.170 173.875 ;
        RECT 40.520 173.515 40.880 173.875 ;
        RECT 41.230 173.515 41.590 173.875 ;
        RECT 41.940 173.515 42.300 173.875 ;
        RECT 42.650 173.515 43.010 173.875 ;
        RECT 43.360 173.515 43.720 173.875 ;
        RECT 44.070 173.515 44.430 173.875 ;
        RECT 44.780 173.515 45.140 173.875 ;
        RECT 45.490 173.515 45.850 173.875 ;
        RECT 46.200 173.515 46.560 173.875 ;
        RECT 46.910 173.515 47.270 173.875 ;
        RECT 47.620 173.515 47.980 173.875 ;
        RECT 48.330 173.515 48.690 173.875 ;
        RECT 49.040 173.515 49.400 173.875 ;
        RECT 49.750 173.515 50.110 173.875 ;
        RECT 50.460 173.515 50.820 173.875 ;
        RECT 51.170 173.515 51.530 173.875 ;
        RECT 51.880 173.515 52.240 173.875 ;
        RECT 52.590 173.515 52.950 173.875 ;
        RECT 53.300 173.515 53.660 173.875 ;
        RECT 54.010 173.515 54.370 173.875 ;
        RECT 54.720 173.515 55.080 173.875 ;
        RECT 55.430 173.515 55.790 173.875 ;
        RECT 56.140 173.515 56.500 173.875 ;
        RECT 56.850 173.515 57.210 173.875 ;
        RECT 57.560 173.515 57.920 173.875 ;
        RECT 58.270 173.515 58.630 173.875 ;
        RECT 58.980 173.515 59.340 173.875 ;
        RECT 59.690 173.515 60.050 173.875 ;
        RECT 60.400 173.515 60.760 173.875 ;
        RECT 61.110 173.515 61.470 173.875 ;
        RECT 61.820 173.515 62.180 173.875 ;
        RECT 62.530 173.515 62.890 173.875 ;
        RECT 63.240 173.515 63.600 173.875 ;
        RECT 63.950 173.515 64.310 173.875 ;
        RECT 64.660 173.515 65.020 173.875 ;
        RECT 65.370 173.515 65.730 173.875 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V3 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.300 66.490 174.000 ;
      LAYER V2 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.300 66.490 174.000 ;
      LAYER V1 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M1 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V5 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V4 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
    END
  END GND
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.600 0.700 113.895 ;
        RECT 0.190 92.280 0.700 100.280 ;
        RECT 0.205 81.280 0.700 89.280 ;
        RECT 0.205 70.000 0.700 79.520 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 110.465 69.415 113.895 ;
        RECT 69.420 150.320 69.675 151.785 ;
        RECT 69.300 152.430 69.685 154.220 ;
        RECT 69.300 81.365 69.740 89.280 ;
        RECT 69.300 70.000 69.740 77.985 ;
        RECT 69.300 115.135 69.780 118.565 ;
        RECT 69.300 105.320 69.780 108.750 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 162.720 69.845 170.465 ;
        RECT 69.300 92.360 69.850 100.195 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 118.565 ;
        RECT 69.420 150.320 70.000 151.785 ;
        RECT 69.560 115.135 70.000 154.220 ;
        RECT 69.300 152.430 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.600 0.700 113.895 ;
        RECT 0.190 92.280 0.700 100.280 ;
        RECT 0.205 81.280 0.700 89.280 ;
        RECT 0.205 70.000 0.700 79.520 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 110.465 69.415 113.895 ;
        RECT 69.420 150.320 69.675 151.785 ;
        RECT 69.300 152.430 69.685 154.220 ;
        RECT 69.300 81.365 69.740 89.280 ;
        RECT 69.300 70.000 69.740 77.985 ;
        RECT 69.300 115.135 69.780 118.565 ;
        RECT 69.300 105.320 69.780 108.750 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 162.720 69.845 170.465 ;
        RECT 69.300 92.360 69.850 100.195 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.600 0.700 113.895 ;
        RECT 0.190 92.280 0.700 100.280 ;
        RECT 0.205 81.280 0.700 89.280 ;
        RECT 0.205 70.000 0.700 79.520 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 110.465 69.415 113.895 ;
        RECT 69.420 150.320 69.675 151.785 ;
        RECT 69.300 152.430 69.685 154.220 ;
        RECT 69.300 81.365 69.740 89.280 ;
        RECT 69.300 70.000 69.740 77.985 ;
        RECT 69.300 115.135 69.780 118.565 ;
        RECT 69.300 105.320 69.780 108.750 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 162.720 69.845 170.465 ;
        RECT 69.300 92.360 69.850 100.195 ;
  END 
END PLVSSC

MACRO PLVDDO
  CLASS  PAD ;
  FOREIGN PLVDDO 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN VDDO
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V6 ;
        RECT 4.310 173.515 4.670 173.875 ;
        RECT 5.020 173.515 5.380 173.875 ;
        RECT 5.730 173.515 6.090 173.875 ;
        RECT 6.440 173.515 6.800 173.875 ;
        RECT 7.150 173.515 7.510 173.875 ;
        RECT 7.860 173.515 8.220 173.875 ;
        RECT 8.570 173.515 8.930 173.875 ;
        RECT 9.280 173.515 9.640 173.875 ;
        RECT 9.990 173.515 10.350 173.875 ;
        RECT 10.700 173.515 11.060 173.875 ;
        RECT 11.410 173.515 11.770 173.875 ;
        RECT 12.120 173.515 12.480 173.875 ;
        RECT 12.830 173.515 13.190 173.875 ;
        RECT 13.540 173.515 13.900 173.875 ;
        RECT 14.250 173.515 14.610 173.875 ;
        RECT 14.960 173.515 15.320 173.875 ;
        RECT 15.670 173.515 16.030 173.875 ;
        RECT 16.380 173.515 16.740 173.875 ;
        RECT 17.090 173.515 17.450 173.875 ;
        RECT 17.800 173.515 18.160 173.875 ;
        RECT 18.510 173.515 18.870 173.875 ;
        RECT 19.220 173.515 19.580 173.875 ;
        RECT 19.930 173.515 20.290 173.875 ;
        RECT 20.640 173.515 21.000 173.875 ;
        RECT 21.350 173.515 21.710 173.875 ;
        RECT 22.060 173.515 22.420 173.875 ;
        RECT 22.770 173.515 23.130 173.875 ;
        RECT 23.480 173.515 23.840 173.875 ;
        RECT 24.190 173.515 24.550 173.875 ;
        RECT 24.900 173.515 25.260 173.875 ;
        RECT 25.610 173.515 25.970 173.875 ;
        RECT 26.320 173.515 26.680 173.875 ;
        RECT 27.030 173.515 27.390 173.875 ;
        RECT 27.740 173.515 28.100 173.875 ;
        RECT 28.450 173.515 28.810 173.875 ;
        RECT 29.160 173.515 29.520 173.875 ;
        RECT 29.870 173.515 30.230 173.875 ;
        RECT 30.580 173.515 30.940 173.875 ;
        RECT 31.290 173.515 31.650 173.875 ;
        RECT 32.000 173.515 32.360 173.875 ;
        RECT 32.710 173.515 33.070 173.875 ;
        RECT 33.420 173.515 33.780 173.875 ;
        RECT 34.130 173.515 34.490 173.875 ;
        RECT 34.840 173.515 35.200 173.875 ;
        RECT 35.550 173.515 35.910 173.875 ;
        RECT 36.260 173.515 36.620 173.875 ;
        RECT 36.970 173.515 37.330 173.875 ;
        RECT 37.680 173.515 38.040 173.875 ;
        RECT 38.390 173.515 38.750 173.875 ;
        RECT 39.100 173.515 39.460 173.875 ;
        RECT 39.810 173.515 40.170 173.875 ;
        RECT 40.520 173.515 40.880 173.875 ;
        RECT 41.230 173.515 41.590 173.875 ;
        RECT 41.940 173.515 42.300 173.875 ;
        RECT 42.650 173.515 43.010 173.875 ;
        RECT 43.360 173.515 43.720 173.875 ;
        RECT 44.070 173.515 44.430 173.875 ;
        RECT 44.780 173.515 45.140 173.875 ;
        RECT 45.490 173.515 45.850 173.875 ;
        RECT 46.200 173.515 46.560 173.875 ;
        RECT 46.910 173.515 47.270 173.875 ;
        RECT 47.620 173.515 47.980 173.875 ;
        RECT 48.330 173.515 48.690 173.875 ;
        RECT 49.040 173.515 49.400 173.875 ;
        RECT 49.750 173.515 50.110 173.875 ;
        RECT 50.460 173.515 50.820 173.875 ;
        RECT 51.170 173.515 51.530 173.875 ;
        RECT 51.880 173.515 52.240 173.875 ;
        RECT 52.590 173.515 52.950 173.875 ;
        RECT 53.300 173.515 53.660 173.875 ;
        RECT 54.010 173.515 54.370 173.875 ;
        RECT 54.720 173.515 55.080 173.875 ;
        RECT 55.430 173.515 55.790 173.875 ;
        RECT 56.140 173.515 56.500 173.875 ;
        RECT 56.850 173.515 57.210 173.875 ;
        RECT 57.560 173.515 57.920 173.875 ;
        RECT 58.270 173.515 58.630 173.875 ;
        RECT 58.980 173.515 59.340 173.875 ;
        RECT 59.690 173.515 60.050 173.875 ;
        RECT 60.400 173.515 60.760 173.875 ;
        RECT 61.110 173.515 61.470 173.875 ;
        RECT 61.820 173.515 62.180 173.875 ;
        RECT 62.530 173.515 62.890 173.875 ;
        RECT 63.240 173.515 63.600 173.875 ;
        RECT 63.950 173.515 64.310 173.875 ;
        RECT 64.660 173.515 65.020 173.875 ;
        RECT 65.370 173.515 65.730 173.875 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V3 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.300 66.490 174.000 ;
      LAYER V2 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.300 66.490 174.000 ;
      LAYER V1 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M1 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V5 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V4 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
    END
  END VDDO
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.700 0.700 154.200 ;
        RECT 0.160 115.135 0.700 119.550 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.320 0.700 100.190 ;
        RECT 0.160 81.280 0.700 89.215 ;
        RECT 0.160 70.000 0.700 78.150 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 152.410 69.745 154.200 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
        RECT 69.300 105.190 69.840 108.790 ;
        RECT 69.300 92.280 69.840 100.265 ;
        RECT 69.300 81.365 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.190 ;
        RECT 69.300 162.720 69.845 170.465 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 119.555 ;
        RECT 0.000 115.135 0.440 154.220 ;
        RECT 0.000 150.700 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.905 ;
        RECT 69.560 115.135 70.000 154.220 ;
        RECT 69.300 152.410 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.700 0.700 154.200 ;
        RECT 0.160 115.135 0.700 119.550 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.320 0.700 100.190 ;
        RECT 0.160 81.280 0.700 89.215 ;
        RECT 0.160 70.000 0.700 78.150 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 152.410 69.745 154.200 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
        RECT 69.300 105.190 69.840 108.790 ;
        RECT 69.300 92.280 69.840 100.265 ;
        RECT 69.300 81.365 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.190 ;
        RECT 69.300 162.720 69.845 170.465 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.700 0.700 154.200 ;
        RECT 0.160 115.135 0.700 119.550 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.320 0.700 100.190 ;
        RECT 0.160 81.280 0.700 89.215 ;
        RECT 0.160 70.000 0.700 78.150 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 152.410 69.745 154.200 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
        RECT 69.300 105.190 69.840 108.790 ;
        RECT 69.300 92.280 69.840 100.265 ;
        RECT 69.300 81.365 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.190 ;
        RECT 69.300 162.720 69.845 170.465 ;
  END 
END PLVDDO

MACRO PLVDDH
  CLASS  PAD ;
  FOREIGN PLVDDH 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN VDDH
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V6 ;
        RECT 4.310 173.515 4.670 173.875 ;
        RECT 5.020 173.515 5.380 173.875 ;
        RECT 5.730 173.515 6.090 173.875 ;
        RECT 6.440 173.515 6.800 173.875 ;
        RECT 7.150 173.515 7.510 173.875 ;
        RECT 7.860 173.515 8.220 173.875 ;
        RECT 8.570 173.515 8.930 173.875 ;
        RECT 9.280 173.515 9.640 173.875 ;
        RECT 9.990 173.515 10.350 173.875 ;
        RECT 10.700 173.515 11.060 173.875 ;
        RECT 11.410 173.515 11.770 173.875 ;
        RECT 12.120 173.515 12.480 173.875 ;
        RECT 12.830 173.515 13.190 173.875 ;
        RECT 13.540 173.515 13.900 173.875 ;
        RECT 14.250 173.515 14.610 173.875 ;
        RECT 14.960 173.515 15.320 173.875 ;
        RECT 15.670 173.515 16.030 173.875 ;
        RECT 16.380 173.515 16.740 173.875 ;
        RECT 17.090 173.515 17.450 173.875 ;
        RECT 17.800 173.515 18.160 173.875 ;
        RECT 18.510 173.515 18.870 173.875 ;
        RECT 19.220 173.515 19.580 173.875 ;
        RECT 19.930 173.515 20.290 173.875 ;
        RECT 20.640 173.515 21.000 173.875 ;
        RECT 21.350 173.515 21.710 173.875 ;
        RECT 22.060 173.515 22.420 173.875 ;
        RECT 22.770 173.515 23.130 173.875 ;
        RECT 23.480 173.515 23.840 173.875 ;
        RECT 24.190 173.515 24.550 173.875 ;
        RECT 24.900 173.515 25.260 173.875 ;
        RECT 25.610 173.515 25.970 173.875 ;
        RECT 26.320 173.515 26.680 173.875 ;
        RECT 27.030 173.515 27.390 173.875 ;
        RECT 27.740 173.515 28.100 173.875 ;
        RECT 28.450 173.515 28.810 173.875 ;
        RECT 29.160 173.515 29.520 173.875 ;
        RECT 29.870 173.515 30.230 173.875 ;
        RECT 30.580 173.515 30.940 173.875 ;
        RECT 31.290 173.515 31.650 173.875 ;
        RECT 32.000 173.515 32.360 173.875 ;
        RECT 32.710 173.515 33.070 173.875 ;
        RECT 33.420 173.515 33.780 173.875 ;
        RECT 34.130 173.515 34.490 173.875 ;
        RECT 34.840 173.515 35.200 173.875 ;
        RECT 35.550 173.515 35.910 173.875 ;
        RECT 36.260 173.515 36.620 173.875 ;
        RECT 36.970 173.515 37.330 173.875 ;
        RECT 37.680 173.515 38.040 173.875 ;
        RECT 38.390 173.515 38.750 173.875 ;
        RECT 39.100 173.515 39.460 173.875 ;
        RECT 39.810 173.515 40.170 173.875 ;
        RECT 40.520 173.515 40.880 173.875 ;
        RECT 41.230 173.515 41.590 173.875 ;
        RECT 41.940 173.515 42.300 173.875 ;
        RECT 42.650 173.515 43.010 173.875 ;
        RECT 43.360 173.515 43.720 173.875 ;
        RECT 44.070 173.515 44.430 173.875 ;
        RECT 44.780 173.515 45.140 173.875 ;
        RECT 45.490 173.515 45.850 173.875 ;
        RECT 46.200 173.515 46.560 173.875 ;
        RECT 46.910 173.515 47.270 173.875 ;
        RECT 47.620 173.515 47.980 173.875 ;
        RECT 48.330 173.515 48.690 173.875 ;
        RECT 49.040 173.515 49.400 173.875 ;
        RECT 49.750 173.515 50.110 173.875 ;
        RECT 50.460 173.515 50.820 173.875 ;
        RECT 51.170 173.515 51.530 173.875 ;
        RECT 51.880 173.515 52.240 173.875 ;
        RECT 52.590 173.515 52.950 173.875 ;
        RECT 53.300 173.515 53.660 173.875 ;
        RECT 54.010 173.515 54.370 173.875 ;
        RECT 54.720 173.515 55.080 173.875 ;
        RECT 55.430 173.515 55.790 173.875 ;
        RECT 56.140 173.515 56.500 173.875 ;
        RECT 56.850 173.515 57.210 173.875 ;
        RECT 57.560 173.515 57.920 173.875 ;
        RECT 58.270 173.515 58.630 173.875 ;
        RECT 58.980 173.515 59.340 173.875 ;
        RECT 59.690 173.515 60.050 173.875 ;
        RECT 60.400 173.515 60.760 173.875 ;
        RECT 61.110 173.515 61.470 173.875 ;
        RECT 61.820 173.515 62.180 173.875 ;
        RECT 62.530 173.515 62.890 173.875 ;
        RECT 63.240 173.515 63.600 173.875 ;
        RECT 63.950 173.515 64.310 173.875 ;
        RECT 64.660 173.515 65.020 173.875 ;
        RECT 65.370 173.515 65.730 173.875 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V3 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.300 66.490 174.000 ;
      LAYER V2 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.300 66.490 174.000 ;
      LAYER V1 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M1 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V5 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V4 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
    END
  END VDDH
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.780 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.455 0.700 100.280 ;
        RECT 0.160 81.355 0.700 89.280 ;
        RECT 0.160 70.000 0.700 77.910 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 152.430 69.755 154.220 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
        RECT 69.300 105.215 69.840 108.815 ;
        RECT 69.300 92.280 69.840 100.180 ;
        RECT 69.300 81.335 69.840 89.130 ;
        RECT 69.300 70.000 69.840 77.940 ;
        RECT 69.300 162.720 69.845 170.465 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 119.710 ;
        RECT 0.000 115.135 0.440 154.220 ;
        RECT 0.000 150.780 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.905 ;
        RECT 69.560 115.135 70.000 154.220 ;
        RECT 69.300 152.430 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.780 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.455 0.700 100.280 ;
        RECT 0.160 81.355 0.700 89.280 ;
        RECT 0.160 70.000 0.700 77.910 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 152.430 69.755 154.220 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
        RECT 69.300 105.215 69.840 108.815 ;
        RECT 69.300 92.280 69.840 100.180 ;
        RECT 69.300 81.335 69.840 89.130 ;
        RECT 69.300 70.000 69.840 77.940 ;
        RECT 69.300 162.720 69.845 170.465 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.780 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.710 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.455 0.700 100.280 ;
        RECT 0.160 81.355 0.700 89.280 ;
        RECT 0.160 70.000 0.700 77.910 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 152.430 69.755 154.220 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
        RECT 69.300 105.215 69.840 108.815 ;
        RECT 69.300 92.280 69.840 100.180 ;
        RECT 69.300 81.335 69.840 89.130 ;
        RECT 69.300 70.000 69.840 77.940 ;
        RECT 69.300 162.720 69.845 170.465 ;
  END 
END PLVDDH

MACRO PLVDDC
  CLASS  PAD ;
  FOREIGN PLVDDC 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    CLASS CORE ;
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V6 ;
        RECT 4.310 173.515 4.670 173.875 ;
        RECT 5.020 173.515 5.380 173.875 ;
        RECT 5.730 173.515 6.090 173.875 ;
        RECT 6.440 173.515 6.800 173.875 ;
        RECT 7.150 173.515 7.510 173.875 ;
        RECT 7.860 173.515 8.220 173.875 ;
        RECT 8.570 173.515 8.930 173.875 ;
        RECT 9.280 173.515 9.640 173.875 ;
        RECT 9.990 173.515 10.350 173.875 ;
        RECT 10.700 173.515 11.060 173.875 ;
        RECT 11.410 173.515 11.770 173.875 ;
        RECT 12.120 173.515 12.480 173.875 ;
        RECT 12.830 173.515 13.190 173.875 ;
        RECT 13.540 173.515 13.900 173.875 ;
        RECT 14.250 173.515 14.610 173.875 ;
        RECT 14.960 173.515 15.320 173.875 ;
        RECT 15.670 173.515 16.030 173.875 ;
        RECT 16.380 173.515 16.740 173.875 ;
        RECT 17.090 173.515 17.450 173.875 ;
        RECT 17.800 173.515 18.160 173.875 ;
        RECT 18.510 173.515 18.870 173.875 ;
        RECT 19.220 173.515 19.580 173.875 ;
        RECT 19.930 173.515 20.290 173.875 ;
        RECT 20.640 173.515 21.000 173.875 ;
        RECT 21.350 173.515 21.710 173.875 ;
        RECT 22.060 173.515 22.420 173.875 ;
        RECT 22.770 173.515 23.130 173.875 ;
        RECT 23.480 173.515 23.840 173.875 ;
        RECT 24.190 173.515 24.550 173.875 ;
        RECT 24.900 173.515 25.260 173.875 ;
        RECT 25.610 173.515 25.970 173.875 ;
        RECT 26.320 173.515 26.680 173.875 ;
        RECT 27.030 173.515 27.390 173.875 ;
        RECT 27.740 173.515 28.100 173.875 ;
        RECT 28.450 173.515 28.810 173.875 ;
        RECT 29.160 173.515 29.520 173.875 ;
        RECT 29.870 173.515 30.230 173.875 ;
        RECT 30.580 173.515 30.940 173.875 ;
        RECT 31.290 173.515 31.650 173.875 ;
        RECT 32.000 173.515 32.360 173.875 ;
        RECT 32.710 173.515 33.070 173.875 ;
        RECT 33.420 173.515 33.780 173.875 ;
        RECT 34.130 173.515 34.490 173.875 ;
        RECT 34.840 173.515 35.200 173.875 ;
        RECT 35.550 173.515 35.910 173.875 ;
        RECT 36.260 173.515 36.620 173.875 ;
        RECT 36.970 173.515 37.330 173.875 ;
        RECT 37.680 173.515 38.040 173.875 ;
        RECT 38.390 173.515 38.750 173.875 ;
        RECT 39.100 173.515 39.460 173.875 ;
        RECT 39.810 173.515 40.170 173.875 ;
        RECT 40.520 173.515 40.880 173.875 ;
        RECT 41.230 173.515 41.590 173.875 ;
        RECT 41.940 173.515 42.300 173.875 ;
        RECT 42.650 173.515 43.010 173.875 ;
        RECT 43.360 173.515 43.720 173.875 ;
        RECT 44.070 173.515 44.430 173.875 ;
        RECT 44.780 173.515 45.140 173.875 ;
        RECT 45.490 173.515 45.850 173.875 ;
        RECT 46.200 173.515 46.560 173.875 ;
        RECT 46.910 173.515 47.270 173.875 ;
        RECT 47.620 173.515 47.980 173.875 ;
        RECT 48.330 173.515 48.690 173.875 ;
        RECT 49.040 173.515 49.400 173.875 ;
        RECT 49.750 173.515 50.110 173.875 ;
        RECT 50.460 173.515 50.820 173.875 ;
        RECT 51.170 173.515 51.530 173.875 ;
        RECT 51.880 173.515 52.240 173.875 ;
        RECT 52.590 173.515 52.950 173.875 ;
        RECT 53.300 173.515 53.660 173.875 ;
        RECT 54.010 173.515 54.370 173.875 ;
        RECT 54.720 173.515 55.080 173.875 ;
        RECT 55.430 173.515 55.790 173.875 ;
        RECT 56.140 173.515 56.500 173.875 ;
        RECT 56.850 173.515 57.210 173.875 ;
        RECT 57.560 173.515 57.920 173.875 ;
        RECT 58.270 173.515 58.630 173.875 ;
        RECT 58.980 173.515 59.340 173.875 ;
        RECT 59.690 173.515 60.050 173.875 ;
        RECT 60.400 173.515 60.760 173.875 ;
        RECT 61.110 173.515 61.470 173.875 ;
        RECT 61.820 173.515 62.180 173.875 ;
        RECT 62.530 173.515 62.890 173.875 ;
        RECT 63.240 173.515 63.600 173.875 ;
        RECT 63.950 173.515 64.310 173.875 ;
        RECT 64.660 173.515 65.020 173.875 ;
        RECT 65.370 173.515 65.730 173.875 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V3 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.300 66.490 174.000 ;
      LAYER V2 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.300 66.490 174.000 ;
      LAYER V1 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M1 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V5 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V4 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
    END
  END VDD
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.690 0.700 154.105 ;
        RECT 0.160 115.135 0.700 119.680 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.290 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.200 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
        RECT 69.300 105.215 69.840 108.815 ;
        RECT 69.300 92.300 69.840 100.280 ;
        RECT 69.300 81.345 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 162.720 69.845 170.465 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 119.680 ;
        RECT 0.000 115.135 0.440 154.220 ;
        RECT 0.000 150.690 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.905 ;
        RECT 69.560 115.135 70.000 154.220 ;
        RECT 69.300 152.945 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.690 0.700 154.105 ;
        RECT 0.160 115.135 0.700 119.680 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.290 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.200 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
        RECT 69.300 105.215 69.840 108.815 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 162.720 69.845 170.465 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.690 0.700 154.105 ;
        RECT 0.160 115.135 0.700 119.680 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.355 0.700 100.280 ;
        RECT 0.160 81.305 0.700 89.145 ;
        RECT 0.160 70.000 0.700 78.200 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
        RECT 69.300 105.215 69.840 108.815 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 162.720 69.845 170.465 ;
  END 
END PLVDDC

MACRO PLSPLIT_OSC
  CLASS  PAD ;
  FOREIGN PLSPLIT_OSC 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 1.100 1.100 68.900 172.900 ;
      LAYER M1 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.295 110.315 0.700 113.895 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 110.315 69.705 113.895 ;
        RECT 69.300 155.725 70.000 161.220 ;
      LAYER M3 ;
        RECT 1.100 1.100 68.900 172.900 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 1.100 1.100 68.900 172.900 ;
  END 
END PLSPLIT_OSC

MACRO PLSPLIT70CON
  CLASS  PAD ;
  FOREIGN PLSPLIT70CON 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.455 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.455 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.455 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
  END 
END PLSPLIT70CON

MACRO PLSPLIT70
  CLASS  PAD ;
  FOREIGN PLSPLIT70 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
      LAYER M1 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
      LAYER M3 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
      LAYER M6 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
      LAYER M5 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
      LAYER M7 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
      LAYER M2 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
  END 
END PLSPLIT70

MACRO PLSPLIT35CON
  CLASS  PAD ;
  FOREIGN PLSPLIT35CON 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.715 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 171.175 34.840 172.780 ;
        RECT 34.300 162.720 34.840 170.715 ;
        RECT 34.300 155.725 34.840 161.220 ;
        RECT 34.300 110.315 34.840 113.895 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 171.175 35.000 172.780 ;
        RECT 34.300 162.720 35.000 170.715 ;
        RECT 34.300 155.725 35.000 161.220 ;
        RECT 34.300 110.315 35.000 113.895 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.715 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 171.175 34.840 172.780 ;
        RECT 34.300 162.720 34.840 170.715 ;
        RECT 34.300 155.725 34.840 161.220 ;
        RECT 34.300 110.315 34.840 113.895 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 171.175 35.000 172.780 ;
        RECT 34.300 162.720 35.000 170.715 ;
        RECT 34.300 155.725 35.000 161.220 ;
        RECT 34.300 150.480 35.000 154.220 ;
        RECT 34.300 115.135 35.000 119.705 ;
        RECT 34.300 110.315 35.000 113.895 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 171.175 35.000 172.780 ;
        RECT 34.300 162.720 35.000 170.715 ;
        RECT 34.300 155.725 35.000 161.220 ;
        RECT 34.300 150.480 35.000 154.220 ;
        RECT 34.300 115.135 35.000 119.705 ;
        RECT 34.300 110.315 35.000 113.895 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 171.175 35.000 172.780 ;
        RECT 34.300 162.720 35.000 170.715 ;
        RECT 34.300 155.725 35.000 161.220 ;
        RECT 34.300 150.480 35.000 154.220 ;
        RECT 34.300 115.135 35.000 119.705 ;
        RECT 34.300 110.315 35.000 113.895 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.715 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 171.175 34.840 172.780 ;
        RECT 34.300 162.720 34.840 170.715 ;
        RECT 34.300 155.725 34.840 161.220 ;
        RECT 34.300 110.315 34.840 113.895 ;
  END 
END PLSPLIT35CON

MACRO PLSPLIT35
  CLASS  PAD ;
  FOREIGN PLSPLIT35 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 155.725 34.840 161.220 ;
        RECT 34.300 110.315 34.840 113.895 ;
      LAYER M1 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 155.725 35.000 161.220 ;
        RECT 34.300 110.315 35.000 113.895 ;
      LAYER M3 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 155.725 34.840 161.220 ;
        RECT 34.300 110.315 34.840 113.895 ;
      LAYER M6 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 155.725 35.000 161.220 ;
        RECT 34.300 150.480 35.000 154.220 ;
        RECT 34.300 115.135 35.000 119.705 ;
        RECT 34.300 110.315 35.000 113.895 ;
      LAYER M5 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 155.725 35.000 161.220 ;
        RECT 34.300 150.480 35.000 154.220 ;
        RECT 34.300 115.135 35.000 119.705 ;
        RECT 34.300 110.315 35.000 113.895 ;
      LAYER M7 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 155.725 35.000 161.220 ;
        RECT 34.300 150.480 35.000 154.220 ;
        RECT 34.300 115.135 35.000 119.705 ;
        RECT 34.300 110.315 35.000 113.895 ;
      LAYER M2 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 155.725 34.840 161.220 ;
        RECT 34.300 110.315 34.840 113.895 ;
  END 
END PLSPLIT35

MACRO PLOSCR14M
  CLASS  PAD ;
  FOREIGN PLOSCR14M 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 167.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN XTALIN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
    END
  END XTALIN
  PIN EI
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 87.270 173.380 88.270 174.000 ;
      LAYER V6 ;
        RECT 87.590 173.510 87.950 173.870 ;
      LAYER M4 ;
        RECT 87.270 173.380 88.270 174.000 ;
      LAYER V3 ;
        RECT 87.470 173.800 87.660 173.990 ;
        RECT 87.470 173.390 87.660 173.580 ;
        RECT 87.880 173.800 88.070 173.990 ;
        RECT 87.880 173.390 88.070 173.580 ;
      LAYER M3 ;
        RECT 87.270 173.380 88.270 174.000 ;
      LAYER V2 ;
        RECT 87.470 173.800 87.660 173.990 ;
        RECT 87.470 173.390 87.660 173.580 ;
        RECT 87.880 173.800 88.070 173.990 ;
        RECT 87.880 173.390 88.070 173.580 ;
      LAYER M2 ;
        RECT 87.670 173.300 87.870 174.000 ;
        RECT 87.270 173.380 88.270 174.000 ;
      LAYER V1 ;
        RECT 87.470 173.800 87.660 173.990 ;
        RECT 87.470 173.390 87.660 173.580 ;
        RECT 87.880 173.800 88.070 173.990 ;
        RECT 87.880 173.390 88.070 173.580 ;
      LAYER M1 ;
        RECT 87.270 173.380 88.270 174.000 ;
      LAYER M6 ;
        RECT 87.270 173.380 88.270 174.000 ;
      LAYER V5 ;
        RECT 87.470 173.800 87.660 173.990 ;
        RECT 87.470 173.390 87.660 173.580 ;
        RECT 87.880 173.800 88.070 173.990 ;
        RECT 87.880 173.390 88.070 173.580 ;
      LAYER M5 ;
        RECT 87.270 173.380 88.270 174.000 ;
      LAYER V4 ;
        RECT 87.470 173.800 87.660 173.990 ;
        RECT 87.470 173.390 87.660 173.580 ;
        RECT 87.880 173.800 88.070 173.990 ;
        RECT 87.880 173.390 88.070 173.580 ;
    END
  END EI
  PIN XTALOUT
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 73.000 0.665 137.000 0.700 ;
        RECT 73.010 0.660 136.995 0.700 ;
        RECT 73.010 0.655 136.985 0.700 ;
        RECT 73.020 0.650 136.985 0.700 ;
        RECT 73.020 0.645 136.975 0.700 ;
        RECT 73.030 0.640 136.975 0.700 ;
        RECT 73.030 0.635 136.965 0.700 ;
        RECT 73.040 0.630 136.965 0.700 ;
        RECT 73.040 0.625 136.955 0.700 ;
        RECT 73.050 0.620 136.955 0.700 ;
        RECT 73.050 0.615 136.945 0.700 ;
        RECT 73.060 0.610 136.945 0.700 ;
        RECT 73.060 0.605 136.935 0.700 ;
        RECT 73.070 0.600 136.935 0.700 ;
        RECT 73.070 0.595 136.925 0.700 ;
        RECT 73.080 0.590 136.925 0.700 ;
        RECT 73.080 0.585 136.915 0.700 ;
        RECT 73.090 0.580 136.915 0.700 ;
        RECT 73.090 0.575 136.905 0.700 ;
        RECT 73.100 0.570 136.905 0.700 ;
        RECT 73.100 0.565 136.895 0.700 ;
        RECT 73.110 0.560 136.895 0.700 ;
        RECT 73.110 0.555 136.885 0.700 ;
        RECT 73.120 0.550 136.885 0.700 ;
        RECT 73.120 0.545 136.875 0.700 ;
        RECT 73.130 0.540 136.875 0.700 ;
        RECT 73.130 0.535 136.865 0.700 ;
        RECT 73.140 0.530 136.865 0.700 ;
        RECT 73.140 0.525 136.855 0.700 ;
        RECT 73.150 0.520 136.855 0.700 ;
        RECT 73.150 0.515 136.845 0.700 ;
        RECT 73.160 0.510 136.845 0.700 ;
        RECT 73.160 0.505 136.835 0.700 ;
        RECT 73.170 0.500 136.835 0.700 ;
        RECT 73.170 0.495 136.825 0.700 ;
        RECT 73.180 0.490 136.825 0.700 ;
        RECT 73.180 0.485 136.815 0.700 ;
        RECT 73.190 0.480 136.815 0.700 ;
        RECT 73.190 0.475 136.805 0.700 ;
        RECT 73.200 0.470 136.805 0.700 ;
        RECT 73.200 0.465 136.795 0.700 ;
        RECT 73.210 0.460 136.795 0.700 ;
        RECT 73.210 0.455 136.785 0.700 ;
        RECT 73.220 0.450 136.785 0.700 ;
        RECT 73.220 0.445 136.775 0.700 ;
        RECT 73.230 0.440 136.775 0.700 ;
        RECT 73.230 0.435 136.765 0.700 ;
        RECT 73.240 0.430 136.765 0.700 ;
        RECT 73.240 0.425 136.755 0.700 ;
        RECT 73.250 0.420 136.755 0.700 ;
        RECT 73.250 0.415 136.745 0.700 ;
        RECT 73.260 0.410 136.745 0.700 ;
        RECT 73.260 0.405 136.735 0.700 ;
        RECT 73.270 0.400 136.735 0.700 ;
        RECT 73.270 0.395 136.725 0.700 ;
        RECT 73.280 0.390 136.725 0.700 ;
        RECT 73.280 0.385 136.715 0.700 ;
        RECT 73.290 0.380 136.715 0.700 ;
        RECT 73.290 0.375 136.705 0.700 ;
        RECT 73.300 0.370 136.705 0.700 ;
        RECT 73.300 0.365 136.695 0.700 ;
        RECT 73.310 0.360 136.695 0.700 ;
        RECT 73.310 0.355 136.685 0.700 ;
        RECT 73.320 0.350 136.685 0.700 ;
        RECT 73.320 0.345 136.675 0.700 ;
        RECT 73.330 0.340 136.675 0.700 ;
        RECT 73.330 0.335 136.665 0.700 ;
        RECT 73.340 0.330 136.665 0.700 ;
        RECT 73.340 0.325 136.655 0.700 ;
        RECT 73.350 0.320 136.655 0.700 ;
        RECT 73.350 0.315 136.645 0.700 ;
        RECT 73.360 0.310 136.645 0.700 ;
        RECT 73.360 0.305 136.635 0.700 ;
        RECT 73.370 0.300 136.635 0.700 ;
        RECT 73.370 0.295 136.625 0.700 ;
        RECT 73.380 0.290 136.625 0.700 ;
        RECT 73.380 0.285 136.615 0.700 ;
        RECT 73.390 0.280 136.615 0.700 ;
        RECT 73.390 0.275 136.605 0.700 ;
        RECT 73.400 0.270 136.605 0.700 ;
        RECT 73.400 0.265 136.595 0.700 ;
        RECT 73.410 0.260 136.595 0.700 ;
        RECT 73.410 0.255 136.585 0.700 ;
        RECT 73.420 0.250 136.585 0.700 ;
        RECT 73.420 0.245 136.575 0.700 ;
        RECT 73.430 0.240 136.575 0.700 ;
        RECT 73.430 0.235 136.565 0.700 ;
        RECT 73.440 0.230 136.565 0.700 ;
        RECT 73.440 0.225 136.555 0.700 ;
        RECT 73.450 0.220 136.555 0.700 ;
        RECT 73.450 0.215 136.545 0.700 ;
        RECT 73.460 0.210 136.545 0.700 ;
        RECT 73.460 0.205 136.535 0.700 ;
        RECT 73.470 0.200 136.535 0.700 ;
        RECT 73.470 0.195 136.525 0.700 ;
        RECT 73.480 0.190 136.525 0.700 ;
        RECT 73.480 0.185 136.515 0.700 ;
        RECT 73.490 0.180 136.515 0.700 ;
        RECT 73.490 0.175 136.505 0.700 ;
        RECT 73.500 0.170 136.505 0.700 ;
        RECT 73.500 0.165 136.495 0.700 ;
        RECT 73.510 0.160 136.495 0.700 ;
        RECT 73.510 0.155 136.485 0.700 ;
        RECT 73.520 0.150 136.485 0.700 ;
        RECT 73.520 0.145 136.475 0.700 ;
        RECT 73.530 0.140 136.475 0.700 ;
        RECT 73.530 0.135 136.465 0.700 ;
        RECT 73.540 0.130 136.465 0.700 ;
        RECT 73.540 0.125 136.455 0.700 ;
        RECT 73.550 0.120 136.455 0.700 ;
        RECT 73.550 0.115 136.445 0.700 ;
        RECT 73.560 0.110 136.445 0.700 ;
        RECT 73.560 0.105 136.435 0.700 ;
        RECT 73.570 0.100 136.435 0.700 ;
        RECT 73.570 0.095 136.425 0.700 ;
        RECT 73.580 0.090 136.425 0.700 ;
        RECT 73.580 0.085 136.415 0.700 ;
        RECT 73.590 0.080 136.415 0.700 ;
        RECT 73.590 0.075 136.405 0.700 ;
        RECT 73.600 0.070 136.405 0.700 ;
        RECT 73.600 0.065 136.395 0.700 ;
        RECT 73.610 0.060 136.395 0.700 ;
        RECT 73.610 0.055 136.385 0.700 ;
        RECT 73.620 0.050 136.385 0.700 ;
        RECT 73.620 0.045 136.375 0.700 ;
        RECT 73.630 0.040 136.375 0.700 ;
        RECT 73.630 0.035 136.365 0.700 ;
        RECT 73.640 0.030 136.365 0.700 ;
        RECT 73.640 0.025 136.355 0.700 ;
        RECT 73.650 0.020 136.355 0.700 ;
        RECT 73.650 0.015 136.345 0.700 ;
        RECT 73.660 0.010 136.345 0.700 ;
        RECT 73.660 0.005 136.335 0.700 ;
        RECT 73.665 0.000 136.335 0.700 ;
      LAYER M4 ;
        RECT 73.000 0.665 137.000 0.700 ;
        RECT 73.010 0.660 136.995 0.700 ;
        RECT 73.010 0.655 136.985 0.700 ;
        RECT 73.020 0.650 136.985 0.700 ;
        RECT 73.020 0.645 136.975 0.700 ;
        RECT 73.030 0.640 136.975 0.700 ;
        RECT 73.030 0.635 136.965 0.700 ;
        RECT 73.040 0.630 136.965 0.700 ;
        RECT 73.040 0.625 136.955 0.700 ;
        RECT 73.050 0.620 136.955 0.700 ;
        RECT 73.050 0.615 136.945 0.700 ;
        RECT 73.060 0.610 136.945 0.700 ;
        RECT 73.060 0.605 136.935 0.700 ;
        RECT 73.070 0.600 136.935 0.700 ;
        RECT 73.070 0.595 136.925 0.700 ;
        RECT 73.080 0.590 136.925 0.700 ;
        RECT 73.080 0.585 136.915 0.700 ;
        RECT 73.090 0.580 136.915 0.700 ;
        RECT 73.090 0.575 136.905 0.700 ;
        RECT 73.100 0.570 136.905 0.700 ;
        RECT 73.100 0.565 136.895 0.700 ;
        RECT 73.110 0.560 136.895 0.700 ;
        RECT 73.110 0.555 136.885 0.700 ;
        RECT 73.120 0.550 136.885 0.700 ;
        RECT 73.120 0.545 136.875 0.700 ;
        RECT 73.130 0.540 136.875 0.700 ;
        RECT 73.130 0.535 136.865 0.700 ;
        RECT 73.140 0.530 136.865 0.700 ;
        RECT 73.140 0.525 136.855 0.700 ;
        RECT 73.150 0.520 136.855 0.700 ;
        RECT 73.150 0.515 136.845 0.700 ;
        RECT 73.160 0.510 136.845 0.700 ;
        RECT 73.160 0.505 136.835 0.700 ;
        RECT 73.170 0.500 136.835 0.700 ;
        RECT 73.170 0.495 136.825 0.700 ;
        RECT 73.180 0.490 136.825 0.700 ;
        RECT 73.180 0.485 136.815 0.700 ;
        RECT 73.190 0.480 136.815 0.700 ;
        RECT 73.190 0.475 136.805 0.700 ;
        RECT 73.200 0.470 136.805 0.700 ;
        RECT 73.200 0.465 136.795 0.700 ;
        RECT 73.210 0.460 136.795 0.700 ;
        RECT 73.210 0.455 136.785 0.700 ;
        RECT 73.220 0.450 136.785 0.700 ;
        RECT 73.220 0.445 136.775 0.700 ;
        RECT 73.230 0.440 136.775 0.700 ;
        RECT 73.230 0.435 136.765 0.700 ;
        RECT 73.240 0.430 136.765 0.700 ;
        RECT 73.240 0.425 136.755 0.700 ;
        RECT 73.250 0.420 136.755 0.700 ;
        RECT 73.250 0.415 136.745 0.700 ;
        RECT 73.260 0.410 136.745 0.700 ;
        RECT 73.260 0.405 136.735 0.700 ;
        RECT 73.270 0.400 136.735 0.700 ;
        RECT 73.270 0.395 136.725 0.700 ;
        RECT 73.280 0.390 136.725 0.700 ;
        RECT 73.280 0.385 136.715 0.700 ;
        RECT 73.290 0.380 136.715 0.700 ;
        RECT 73.290 0.375 136.705 0.700 ;
        RECT 73.300 0.370 136.705 0.700 ;
        RECT 73.300 0.365 136.695 0.700 ;
        RECT 73.310 0.360 136.695 0.700 ;
        RECT 73.310 0.355 136.685 0.700 ;
        RECT 73.320 0.350 136.685 0.700 ;
        RECT 73.320 0.345 136.675 0.700 ;
        RECT 73.330 0.340 136.675 0.700 ;
        RECT 73.330 0.335 136.665 0.700 ;
        RECT 73.340 0.330 136.665 0.700 ;
        RECT 73.340 0.325 136.655 0.700 ;
        RECT 73.350 0.320 136.655 0.700 ;
        RECT 73.350 0.315 136.645 0.700 ;
        RECT 73.360 0.310 136.645 0.700 ;
        RECT 73.360 0.305 136.635 0.700 ;
        RECT 73.370 0.300 136.635 0.700 ;
        RECT 73.370 0.295 136.625 0.700 ;
        RECT 73.380 0.290 136.625 0.700 ;
        RECT 73.380 0.285 136.615 0.700 ;
        RECT 73.390 0.280 136.615 0.700 ;
        RECT 73.390 0.275 136.605 0.700 ;
        RECT 73.400 0.270 136.605 0.700 ;
        RECT 73.400 0.265 136.595 0.700 ;
        RECT 73.410 0.260 136.595 0.700 ;
        RECT 73.410 0.255 136.585 0.700 ;
        RECT 73.420 0.250 136.585 0.700 ;
        RECT 73.420 0.245 136.575 0.700 ;
        RECT 73.430 0.240 136.575 0.700 ;
        RECT 73.430 0.235 136.565 0.700 ;
        RECT 73.440 0.230 136.565 0.700 ;
        RECT 73.440 0.225 136.555 0.700 ;
        RECT 73.450 0.220 136.555 0.700 ;
        RECT 73.450 0.215 136.545 0.700 ;
        RECT 73.460 0.210 136.545 0.700 ;
        RECT 73.460 0.205 136.535 0.700 ;
        RECT 73.470 0.200 136.535 0.700 ;
        RECT 73.470 0.195 136.525 0.700 ;
        RECT 73.480 0.190 136.525 0.700 ;
        RECT 73.480 0.185 136.515 0.700 ;
        RECT 73.490 0.180 136.515 0.700 ;
        RECT 73.490 0.175 136.505 0.700 ;
        RECT 73.500 0.170 136.505 0.700 ;
        RECT 73.500 0.165 136.495 0.700 ;
        RECT 73.510 0.160 136.495 0.700 ;
        RECT 73.510 0.155 136.485 0.700 ;
        RECT 73.520 0.150 136.485 0.700 ;
        RECT 73.520 0.145 136.475 0.700 ;
        RECT 73.530 0.140 136.475 0.700 ;
        RECT 73.530 0.135 136.465 0.700 ;
        RECT 73.540 0.130 136.465 0.700 ;
        RECT 73.540 0.125 136.455 0.700 ;
        RECT 73.550 0.120 136.455 0.700 ;
        RECT 73.550 0.115 136.445 0.700 ;
        RECT 73.560 0.110 136.445 0.700 ;
        RECT 73.560 0.105 136.435 0.700 ;
        RECT 73.570 0.100 136.435 0.700 ;
        RECT 73.570 0.095 136.425 0.700 ;
        RECT 73.580 0.090 136.425 0.700 ;
        RECT 73.580 0.085 136.415 0.700 ;
        RECT 73.590 0.080 136.415 0.700 ;
        RECT 73.590 0.075 136.405 0.700 ;
        RECT 73.600 0.070 136.405 0.700 ;
        RECT 73.600 0.065 136.395 0.700 ;
        RECT 73.610 0.060 136.395 0.700 ;
        RECT 73.610 0.055 136.385 0.700 ;
        RECT 73.620 0.050 136.385 0.700 ;
        RECT 73.620 0.045 136.375 0.700 ;
        RECT 73.630 0.040 136.375 0.700 ;
        RECT 73.630 0.035 136.365 0.700 ;
        RECT 73.640 0.030 136.365 0.700 ;
        RECT 73.640 0.025 136.355 0.700 ;
        RECT 73.650 0.020 136.355 0.700 ;
        RECT 73.650 0.015 136.345 0.700 ;
        RECT 73.660 0.010 136.345 0.700 ;
        RECT 73.660 0.005 136.335 0.700 ;
        RECT 73.665 0.000 136.335 0.700 ;
      LAYER M3 ;
        RECT 73.000 0.665 137.000 0.700 ;
        RECT 73.010 0.660 136.995 0.700 ;
        RECT 73.010 0.655 136.985 0.700 ;
        RECT 73.020 0.650 136.985 0.700 ;
        RECT 73.020 0.645 136.975 0.700 ;
        RECT 73.030 0.640 136.975 0.700 ;
        RECT 73.030 0.635 136.965 0.700 ;
        RECT 73.040 0.630 136.965 0.700 ;
        RECT 73.040 0.625 136.955 0.700 ;
        RECT 73.050 0.620 136.955 0.700 ;
        RECT 73.050 0.615 136.945 0.700 ;
        RECT 73.060 0.610 136.945 0.700 ;
        RECT 73.060 0.605 136.935 0.700 ;
        RECT 73.070 0.600 136.935 0.700 ;
        RECT 73.070 0.595 136.925 0.700 ;
        RECT 73.080 0.590 136.925 0.700 ;
        RECT 73.080 0.585 136.915 0.700 ;
        RECT 73.090 0.580 136.915 0.700 ;
        RECT 73.090 0.575 136.905 0.700 ;
        RECT 73.100 0.570 136.905 0.700 ;
        RECT 73.100 0.565 136.895 0.700 ;
        RECT 73.110 0.560 136.895 0.700 ;
        RECT 73.110 0.555 136.885 0.700 ;
        RECT 73.120 0.550 136.885 0.700 ;
        RECT 73.120 0.545 136.875 0.700 ;
        RECT 73.130 0.540 136.875 0.700 ;
        RECT 73.130 0.535 136.865 0.700 ;
        RECT 73.140 0.530 136.865 0.700 ;
        RECT 73.140 0.525 136.855 0.700 ;
        RECT 73.150 0.520 136.855 0.700 ;
        RECT 73.150 0.515 136.845 0.700 ;
        RECT 73.160 0.510 136.845 0.700 ;
        RECT 73.160 0.505 136.835 0.700 ;
        RECT 73.170 0.500 136.835 0.700 ;
        RECT 73.170 0.495 136.825 0.700 ;
        RECT 73.180 0.490 136.825 0.700 ;
        RECT 73.180 0.485 136.815 0.700 ;
        RECT 73.190 0.480 136.815 0.700 ;
        RECT 73.190 0.475 136.805 0.700 ;
        RECT 73.200 0.470 136.805 0.700 ;
        RECT 73.200 0.465 136.795 0.700 ;
        RECT 73.210 0.460 136.795 0.700 ;
        RECT 73.210 0.455 136.785 0.700 ;
        RECT 73.220 0.450 136.785 0.700 ;
        RECT 73.220 0.445 136.775 0.700 ;
        RECT 73.230 0.440 136.775 0.700 ;
        RECT 73.230 0.435 136.765 0.700 ;
        RECT 73.240 0.430 136.765 0.700 ;
        RECT 73.240 0.425 136.755 0.700 ;
        RECT 73.250 0.420 136.755 0.700 ;
        RECT 73.250 0.415 136.745 0.700 ;
        RECT 73.260 0.410 136.745 0.700 ;
        RECT 73.260 0.405 136.735 0.700 ;
        RECT 73.270 0.400 136.735 0.700 ;
        RECT 73.270 0.395 136.725 0.700 ;
        RECT 73.280 0.390 136.725 0.700 ;
        RECT 73.280 0.385 136.715 0.700 ;
        RECT 73.290 0.380 136.715 0.700 ;
        RECT 73.290 0.375 136.705 0.700 ;
        RECT 73.300 0.370 136.705 0.700 ;
        RECT 73.300 0.365 136.695 0.700 ;
        RECT 73.310 0.360 136.695 0.700 ;
        RECT 73.310 0.355 136.685 0.700 ;
        RECT 73.320 0.350 136.685 0.700 ;
        RECT 73.320 0.345 136.675 0.700 ;
        RECT 73.330 0.340 136.675 0.700 ;
        RECT 73.330 0.335 136.665 0.700 ;
        RECT 73.340 0.330 136.665 0.700 ;
        RECT 73.340 0.325 136.655 0.700 ;
        RECT 73.350 0.320 136.655 0.700 ;
        RECT 73.350 0.315 136.645 0.700 ;
        RECT 73.360 0.310 136.645 0.700 ;
        RECT 73.360 0.305 136.635 0.700 ;
        RECT 73.370 0.300 136.635 0.700 ;
        RECT 73.370 0.295 136.625 0.700 ;
        RECT 73.380 0.290 136.625 0.700 ;
        RECT 73.380 0.285 136.615 0.700 ;
        RECT 73.390 0.280 136.615 0.700 ;
        RECT 73.390 0.275 136.605 0.700 ;
        RECT 73.400 0.270 136.605 0.700 ;
        RECT 73.400 0.265 136.595 0.700 ;
        RECT 73.410 0.260 136.595 0.700 ;
        RECT 73.410 0.255 136.585 0.700 ;
        RECT 73.420 0.250 136.585 0.700 ;
        RECT 73.420 0.245 136.575 0.700 ;
        RECT 73.430 0.240 136.575 0.700 ;
        RECT 73.430 0.235 136.565 0.700 ;
        RECT 73.440 0.230 136.565 0.700 ;
        RECT 73.440 0.225 136.555 0.700 ;
        RECT 73.450 0.220 136.555 0.700 ;
        RECT 73.450 0.215 136.545 0.700 ;
        RECT 73.460 0.210 136.545 0.700 ;
        RECT 73.460 0.205 136.535 0.700 ;
        RECT 73.470 0.200 136.535 0.700 ;
        RECT 73.470 0.195 136.525 0.700 ;
        RECT 73.480 0.190 136.525 0.700 ;
        RECT 73.480 0.185 136.515 0.700 ;
        RECT 73.490 0.180 136.515 0.700 ;
        RECT 73.490 0.175 136.505 0.700 ;
        RECT 73.500 0.170 136.505 0.700 ;
        RECT 73.500 0.165 136.495 0.700 ;
        RECT 73.510 0.160 136.495 0.700 ;
        RECT 73.510 0.155 136.485 0.700 ;
        RECT 73.520 0.150 136.485 0.700 ;
        RECT 73.520 0.145 136.475 0.700 ;
        RECT 73.530 0.140 136.475 0.700 ;
        RECT 73.530 0.135 136.465 0.700 ;
        RECT 73.540 0.130 136.465 0.700 ;
        RECT 73.540 0.125 136.455 0.700 ;
        RECT 73.550 0.120 136.455 0.700 ;
        RECT 73.550 0.115 136.445 0.700 ;
        RECT 73.560 0.110 136.445 0.700 ;
        RECT 73.560 0.105 136.435 0.700 ;
        RECT 73.570 0.100 136.435 0.700 ;
        RECT 73.570 0.095 136.425 0.700 ;
        RECT 73.580 0.090 136.425 0.700 ;
        RECT 73.580 0.085 136.415 0.700 ;
        RECT 73.590 0.080 136.415 0.700 ;
        RECT 73.590 0.075 136.405 0.700 ;
        RECT 73.600 0.070 136.405 0.700 ;
        RECT 73.600 0.065 136.395 0.700 ;
        RECT 73.610 0.060 136.395 0.700 ;
        RECT 73.610 0.055 136.385 0.700 ;
        RECT 73.620 0.050 136.385 0.700 ;
        RECT 73.620 0.045 136.375 0.700 ;
        RECT 73.630 0.040 136.375 0.700 ;
        RECT 73.630 0.035 136.365 0.700 ;
        RECT 73.640 0.030 136.365 0.700 ;
        RECT 73.640 0.025 136.355 0.700 ;
        RECT 73.650 0.020 136.355 0.700 ;
        RECT 73.650 0.015 136.345 0.700 ;
        RECT 73.660 0.010 136.345 0.700 ;
        RECT 73.660 0.005 136.335 0.700 ;
        RECT 73.665 0.000 136.335 0.700 ;
      LAYER M2 ;
        RECT 73.000 0.665 137.000 0.700 ;
        RECT 73.010 0.660 136.995 0.700 ;
        RECT 73.010 0.655 136.985 0.700 ;
        RECT 73.020 0.650 136.985 0.700 ;
        RECT 73.020 0.645 136.975 0.700 ;
        RECT 73.030 0.640 136.975 0.700 ;
        RECT 73.030 0.635 136.965 0.700 ;
        RECT 73.040 0.630 136.965 0.700 ;
        RECT 73.040 0.625 136.955 0.700 ;
        RECT 73.050 0.620 136.955 0.700 ;
        RECT 73.050 0.615 136.945 0.700 ;
        RECT 73.060 0.610 136.945 0.700 ;
        RECT 73.060 0.605 136.935 0.700 ;
        RECT 73.070 0.600 136.935 0.700 ;
        RECT 73.070 0.595 136.925 0.700 ;
        RECT 73.080 0.590 136.925 0.700 ;
        RECT 73.080 0.585 136.915 0.700 ;
        RECT 73.090 0.580 136.915 0.700 ;
        RECT 73.090 0.575 136.905 0.700 ;
        RECT 73.100 0.570 136.905 0.700 ;
        RECT 73.100 0.565 136.895 0.700 ;
        RECT 73.110 0.560 136.895 0.700 ;
        RECT 73.110 0.555 136.885 0.700 ;
        RECT 73.120 0.550 136.885 0.700 ;
        RECT 73.120 0.545 136.875 0.700 ;
        RECT 73.130 0.540 136.875 0.700 ;
        RECT 73.130 0.535 136.865 0.700 ;
        RECT 73.140 0.530 136.865 0.700 ;
        RECT 73.140 0.525 136.855 0.700 ;
        RECT 73.150 0.520 136.855 0.700 ;
        RECT 73.150 0.515 136.845 0.700 ;
        RECT 73.160 0.510 136.845 0.700 ;
        RECT 73.160 0.505 136.835 0.700 ;
        RECT 73.170 0.500 136.835 0.700 ;
        RECT 73.170 0.495 136.825 0.700 ;
        RECT 73.180 0.490 136.825 0.700 ;
        RECT 73.180 0.485 136.815 0.700 ;
        RECT 73.190 0.480 136.815 0.700 ;
        RECT 73.190 0.475 136.805 0.700 ;
        RECT 73.200 0.470 136.805 0.700 ;
        RECT 73.200 0.465 136.795 0.700 ;
        RECT 73.210 0.460 136.795 0.700 ;
        RECT 73.210 0.455 136.785 0.700 ;
        RECT 73.220 0.450 136.785 0.700 ;
        RECT 73.220 0.445 136.775 0.700 ;
        RECT 73.230 0.440 136.775 0.700 ;
        RECT 73.230 0.435 136.765 0.700 ;
        RECT 73.240 0.430 136.765 0.700 ;
        RECT 73.240 0.425 136.755 0.700 ;
        RECT 73.250 0.420 136.755 0.700 ;
        RECT 73.250 0.415 136.745 0.700 ;
        RECT 73.260 0.410 136.745 0.700 ;
        RECT 73.260 0.405 136.735 0.700 ;
        RECT 73.270 0.400 136.735 0.700 ;
        RECT 73.270 0.395 136.725 0.700 ;
        RECT 73.280 0.390 136.725 0.700 ;
        RECT 73.280 0.385 136.715 0.700 ;
        RECT 73.290 0.380 136.715 0.700 ;
        RECT 73.290 0.375 136.705 0.700 ;
        RECT 73.300 0.370 136.705 0.700 ;
        RECT 73.300 0.365 136.695 0.700 ;
        RECT 73.310 0.360 136.695 0.700 ;
        RECT 73.310 0.355 136.685 0.700 ;
        RECT 73.320 0.350 136.685 0.700 ;
        RECT 73.320 0.345 136.675 0.700 ;
        RECT 73.330 0.340 136.675 0.700 ;
        RECT 73.330 0.335 136.665 0.700 ;
        RECT 73.340 0.330 136.665 0.700 ;
        RECT 73.340 0.325 136.655 0.700 ;
        RECT 73.350 0.320 136.655 0.700 ;
        RECT 73.350 0.315 136.645 0.700 ;
        RECT 73.360 0.310 136.645 0.700 ;
        RECT 73.360 0.305 136.635 0.700 ;
        RECT 73.370 0.300 136.635 0.700 ;
        RECT 73.370 0.295 136.625 0.700 ;
        RECT 73.380 0.290 136.625 0.700 ;
        RECT 73.380 0.285 136.615 0.700 ;
        RECT 73.390 0.280 136.615 0.700 ;
        RECT 73.390 0.275 136.605 0.700 ;
        RECT 73.400 0.270 136.605 0.700 ;
        RECT 73.400 0.265 136.595 0.700 ;
        RECT 73.410 0.260 136.595 0.700 ;
        RECT 73.410 0.255 136.585 0.700 ;
        RECT 73.420 0.250 136.585 0.700 ;
        RECT 73.420 0.245 136.575 0.700 ;
        RECT 73.430 0.240 136.575 0.700 ;
        RECT 73.430 0.235 136.565 0.700 ;
        RECT 73.440 0.230 136.565 0.700 ;
        RECT 73.440 0.225 136.555 0.700 ;
        RECT 73.450 0.220 136.555 0.700 ;
        RECT 73.450 0.215 136.545 0.700 ;
        RECT 73.460 0.210 136.545 0.700 ;
        RECT 73.460 0.205 136.535 0.700 ;
        RECT 73.470 0.200 136.535 0.700 ;
        RECT 73.470 0.195 136.525 0.700 ;
        RECT 73.480 0.190 136.525 0.700 ;
        RECT 73.480 0.185 136.515 0.700 ;
        RECT 73.490 0.180 136.515 0.700 ;
        RECT 73.490 0.175 136.505 0.700 ;
        RECT 73.500 0.170 136.505 0.700 ;
        RECT 73.500 0.165 136.495 0.700 ;
        RECT 73.510 0.160 136.495 0.700 ;
        RECT 73.510 0.155 136.485 0.700 ;
        RECT 73.520 0.150 136.485 0.700 ;
        RECT 73.520 0.145 136.475 0.700 ;
        RECT 73.530 0.140 136.475 0.700 ;
        RECT 73.530 0.135 136.465 0.700 ;
        RECT 73.540 0.130 136.465 0.700 ;
        RECT 73.540 0.125 136.455 0.700 ;
        RECT 73.550 0.120 136.455 0.700 ;
        RECT 73.550 0.115 136.445 0.700 ;
        RECT 73.560 0.110 136.445 0.700 ;
        RECT 73.560 0.105 136.435 0.700 ;
        RECT 73.570 0.100 136.435 0.700 ;
        RECT 73.570 0.095 136.425 0.700 ;
        RECT 73.580 0.090 136.425 0.700 ;
        RECT 73.580 0.085 136.415 0.700 ;
        RECT 73.590 0.080 136.415 0.700 ;
        RECT 73.590 0.075 136.405 0.700 ;
        RECT 73.600 0.070 136.405 0.700 ;
        RECT 73.600 0.065 136.395 0.700 ;
        RECT 73.610 0.060 136.395 0.700 ;
        RECT 73.610 0.055 136.385 0.700 ;
        RECT 73.620 0.050 136.385 0.700 ;
        RECT 73.620 0.045 136.375 0.700 ;
        RECT 73.630 0.040 136.375 0.700 ;
        RECT 73.630 0.035 136.365 0.700 ;
        RECT 73.640 0.030 136.365 0.700 ;
        RECT 73.640 0.025 136.355 0.700 ;
        RECT 73.650 0.020 136.355 0.700 ;
        RECT 73.650 0.015 136.345 0.700 ;
        RECT 73.660 0.010 136.345 0.700 ;
        RECT 73.660 0.005 136.335 0.700 ;
        RECT 73.665 0.000 136.335 0.700 ;
      LAYER M6 ;
        RECT 73.000 0.665 137.000 0.700 ;
        RECT 73.010 0.660 136.995 0.700 ;
        RECT 73.010 0.655 136.985 0.700 ;
        RECT 73.020 0.650 136.985 0.700 ;
        RECT 73.020 0.645 136.975 0.700 ;
        RECT 73.030 0.640 136.975 0.700 ;
        RECT 73.030 0.635 136.965 0.700 ;
        RECT 73.040 0.630 136.965 0.700 ;
        RECT 73.040 0.625 136.955 0.700 ;
        RECT 73.050 0.620 136.955 0.700 ;
        RECT 73.050 0.615 136.945 0.700 ;
        RECT 73.060 0.610 136.945 0.700 ;
        RECT 73.060 0.605 136.935 0.700 ;
        RECT 73.070 0.600 136.935 0.700 ;
        RECT 73.070 0.595 136.925 0.700 ;
        RECT 73.080 0.590 136.925 0.700 ;
        RECT 73.080 0.585 136.915 0.700 ;
        RECT 73.090 0.580 136.915 0.700 ;
        RECT 73.090 0.575 136.905 0.700 ;
        RECT 73.100 0.570 136.905 0.700 ;
        RECT 73.100 0.565 136.895 0.700 ;
        RECT 73.110 0.560 136.895 0.700 ;
        RECT 73.110 0.555 136.885 0.700 ;
        RECT 73.120 0.550 136.885 0.700 ;
        RECT 73.120 0.545 136.875 0.700 ;
        RECT 73.130 0.540 136.875 0.700 ;
        RECT 73.130 0.535 136.865 0.700 ;
        RECT 73.140 0.530 136.865 0.700 ;
        RECT 73.140 0.525 136.855 0.700 ;
        RECT 73.150 0.520 136.855 0.700 ;
        RECT 73.150 0.515 136.845 0.700 ;
        RECT 73.160 0.510 136.845 0.700 ;
        RECT 73.160 0.505 136.835 0.700 ;
        RECT 73.170 0.500 136.835 0.700 ;
        RECT 73.170 0.495 136.825 0.700 ;
        RECT 73.180 0.490 136.825 0.700 ;
        RECT 73.180 0.485 136.815 0.700 ;
        RECT 73.190 0.480 136.815 0.700 ;
        RECT 73.190 0.475 136.805 0.700 ;
        RECT 73.200 0.470 136.805 0.700 ;
        RECT 73.200 0.465 136.795 0.700 ;
        RECT 73.210 0.460 136.795 0.700 ;
        RECT 73.210 0.455 136.785 0.700 ;
        RECT 73.220 0.450 136.785 0.700 ;
        RECT 73.220 0.445 136.775 0.700 ;
        RECT 73.230 0.440 136.775 0.700 ;
        RECT 73.230 0.435 136.765 0.700 ;
        RECT 73.240 0.430 136.765 0.700 ;
        RECT 73.240 0.425 136.755 0.700 ;
        RECT 73.250 0.420 136.755 0.700 ;
        RECT 73.250 0.415 136.745 0.700 ;
        RECT 73.260 0.410 136.745 0.700 ;
        RECT 73.260 0.405 136.735 0.700 ;
        RECT 73.270 0.400 136.735 0.700 ;
        RECT 73.270 0.395 136.725 0.700 ;
        RECT 73.280 0.390 136.725 0.700 ;
        RECT 73.280 0.385 136.715 0.700 ;
        RECT 73.290 0.380 136.715 0.700 ;
        RECT 73.290 0.375 136.705 0.700 ;
        RECT 73.300 0.370 136.705 0.700 ;
        RECT 73.300 0.365 136.695 0.700 ;
        RECT 73.310 0.360 136.695 0.700 ;
        RECT 73.310 0.355 136.685 0.700 ;
        RECT 73.320 0.350 136.685 0.700 ;
        RECT 73.320 0.345 136.675 0.700 ;
        RECT 73.330 0.340 136.675 0.700 ;
        RECT 73.330 0.335 136.665 0.700 ;
        RECT 73.340 0.330 136.665 0.700 ;
        RECT 73.340 0.325 136.655 0.700 ;
        RECT 73.350 0.320 136.655 0.700 ;
        RECT 73.350 0.315 136.645 0.700 ;
        RECT 73.360 0.310 136.645 0.700 ;
        RECT 73.360 0.305 136.635 0.700 ;
        RECT 73.370 0.300 136.635 0.700 ;
        RECT 73.370 0.295 136.625 0.700 ;
        RECT 73.380 0.290 136.625 0.700 ;
        RECT 73.380 0.285 136.615 0.700 ;
        RECT 73.390 0.280 136.615 0.700 ;
        RECT 73.390 0.275 136.605 0.700 ;
        RECT 73.400 0.270 136.605 0.700 ;
        RECT 73.400 0.265 136.595 0.700 ;
        RECT 73.410 0.260 136.595 0.700 ;
        RECT 73.410 0.255 136.585 0.700 ;
        RECT 73.420 0.250 136.585 0.700 ;
        RECT 73.420 0.245 136.575 0.700 ;
        RECT 73.430 0.240 136.575 0.700 ;
        RECT 73.430 0.235 136.565 0.700 ;
        RECT 73.440 0.230 136.565 0.700 ;
        RECT 73.440 0.225 136.555 0.700 ;
        RECT 73.450 0.220 136.555 0.700 ;
        RECT 73.450 0.215 136.545 0.700 ;
        RECT 73.460 0.210 136.545 0.700 ;
        RECT 73.460 0.205 136.535 0.700 ;
        RECT 73.470 0.200 136.535 0.700 ;
        RECT 73.470 0.195 136.525 0.700 ;
        RECT 73.480 0.190 136.525 0.700 ;
        RECT 73.480 0.185 136.515 0.700 ;
        RECT 73.490 0.180 136.515 0.700 ;
        RECT 73.490 0.175 136.505 0.700 ;
        RECT 73.500 0.170 136.505 0.700 ;
        RECT 73.500 0.165 136.495 0.700 ;
        RECT 73.510 0.160 136.495 0.700 ;
        RECT 73.510 0.155 136.485 0.700 ;
        RECT 73.520 0.150 136.485 0.700 ;
        RECT 73.520 0.145 136.475 0.700 ;
        RECT 73.530 0.140 136.475 0.700 ;
        RECT 73.530 0.135 136.465 0.700 ;
        RECT 73.540 0.130 136.465 0.700 ;
        RECT 73.540 0.125 136.455 0.700 ;
        RECT 73.550 0.120 136.455 0.700 ;
        RECT 73.550 0.115 136.445 0.700 ;
        RECT 73.560 0.110 136.445 0.700 ;
        RECT 73.560 0.105 136.435 0.700 ;
        RECT 73.570 0.100 136.435 0.700 ;
        RECT 73.570 0.095 136.425 0.700 ;
        RECT 73.580 0.090 136.425 0.700 ;
        RECT 73.580 0.085 136.415 0.700 ;
        RECT 73.590 0.080 136.415 0.700 ;
        RECT 73.590 0.075 136.405 0.700 ;
        RECT 73.600 0.070 136.405 0.700 ;
        RECT 73.600 0.065 136.395 0.700 ;
        RECT 73.610 0.060 136.395 0.700 ;
        RECT 73.610 0.055 136.385 0.700 ;
        RECT 73.620 0.050 136.385 0.700 ;
        RECT 73.620 0.045 136.375 0.700 ;
        RECT 73.630 0.040 136.375 0.700 ;
        RECT 73.630 0.035 136.365 0.700 ;
        RECT 73.640 0.030 136.365 0.700 ;
        RECT 73.640 0.025 136.355 0.700 ;
        RECT 73.650 0.020 136.355 0.700 ;
        RECT 73.650 0.015 136.345 0.700 ;
        RECT 73.660 0.010 136.345 0.700 ;
        RECT 73.660 0.005 136.335 0.700 ;
        RECT 73.665 0.000 136.335 0.700 ;
      LAYER M5 ;
        RECT 73.000 0.665 137.000 0.700 ;
        RECT 73.010 0.660 136.995 0.700 ;
        RECT 73.010 0.655 136.985 0.700 ;
        RECT 73.020 0.650 136.985 0.700 ;
        RECT 73.020 0.645 136.975 0.700 ;
        RECT 73.030 0.640 136.975 0.700 ;
        RECT 73.030 0.635 136.965 0.700 ;
        RECT 73.040 0.630 136.965 0.700 ;
        RECT 73.040 0.625 136.955 0.700 ;
        RECT 73.050 0.620 136.955 0.700 ;
        RECT 73.050 0.615 136.945 0.700 ;
        RECT 73.060 0.610 136.945 0.700 ;
        RECT 73.060 0.605 136.935 0.700 ;
        RECT 73.070 0.600 136.935 0.700 ;
        RECT 73.070 0.595 136.925 0.700 ;
        RECT 73.080 0.590 136.925 0.700 ;
        RECT 73.080 0.585 136.915 0.700 ;
        RECT 73.090 0.580 136.915 0.700 ;
        RECT 73.090 0.575 136.905 0.700 ;
        RECT 73.100 0.570 136.905 0.700 ;
        RECT 73.100 0.565 136.895 0.700 ;
        RECT 73.110 0.560 136.895 0.700 ;
        RECT 73.110 0.555 136.885 0.700 ;
        RECT 73.120 0.550 136.885 0.700 ;
        RECT 73.120 0.545 136.875 0.700 ;
        RECT 73.130 0.540 136.875 0.700 ;
        RECT 73.130 0.535 136.865 0.700 ;
        RECT 73.140 0.530 136.865 0.700 ;
        RECT 73.140 0.525 136.855 0.700 ;
        RECT 73.150 0.520 136.855 0.700 ;
        RECT 73.150 0.515 136.845 0.700 ;
        RECT 73.160 0.510 136.845 0.700 ;
        RECT 73.160 0.505 136.835 0.700 ;
        RECT 73.170 0.500 136.835 0.700 ;
        RECT 73.170 0.495 136.825 0.700 ;
        RECT 73.180 0.490 136.825 0.700 ;
        RECT 73.180 0.485 136.815 0.700 ;
        RECT 73.190 0.480 136.815 0.700 ;
        RECT 73.190 0.475 136.805 0.700 ;
        RECT 73.200 0.470 136.805 0.700 ;
        RECT 73.200 0.465 136.795 0.700 ;
        RECT 73.210 0.460 136.795 0.700 ;
        RECT 73.210 0.455 136.785 0.700 ;
        RECT 73.220 0.450 136.785 0.700 ;
        RECT 73.220 0.445 136.775 0.700 ;
        RECT 73.230 0.440 136.775 0.700 ;
        RECT 73.230 0.435 136.765 0.700 ;
        RECT 73.240 0.430 136.765 0.700 ;
        RECT 73.240 0.425 136.755 0.700 ;
        RECT 73.250 0.420 136.755 0.700 ;
        RECT 73.250 0.415 136.745 0.700 ;
        RECT 73.260 0.410 136.745 0.700 ;
        RECT 73.260 0.405 136.735 0.700 ;
        RECT 73.270 0.400 136.735 0.700 ;
        RECT 73.270 0.395 136.725 0.700 ;
        RECT 73.280 0.390 136.725 0.700 ;
        RECT 73.280 0.385 136.715 0.700 ;
        RECT 73.290 0.380 136.715 0.700 ;
        RECT 73.290 0.375 136.705 0.700 ;
        RECT 73.300 0.370 136.705 0.700 ;
        RECT 73.300 0.365 136.695 0.700 ;
        RECT 73.310 0.360 136.695 0.700 ;
        RECT 73.310 0.355 136.685 0.700 ;
        RECT 73.320 0.350 136.685 0.700 ;
        RECT 73.320 0.345 136.675 0.700 ;
        RECT 73.330 0.340 136.675 0.700 ;
        RECT 73.330 0.335 136.665 0.700 ;
        RECT 73.340 0.330 136.665 0.700 ;
        RECT 73.340 0.325 136.655 0.700 ;
        RECT 73.350 0.320 136.655 0.700 ;
        RECT 73.350 0.315 136.645 0.700 ;
        RECT 73.360 0.310 136.645 0.700 ;
        RECT 73.360 0.305 136.635 0.700 ;
        RECT 73.370 0.300 136.635 0.700 ;
        RECT 73.370 0.295 136.625 0.700 ;
        RECT 73.380 0.290 136.625 0.700 ;
        RECT 73.380 0.285 136.615 0.700 ;
        RECT 73.390 0.280 136.615 0.700 ;
        RECT 73.390 0.275 136.605 0.700 ;
        RECT 73.400 0.270 136.605 0.700 ;
        RECT 73.400 0.265 136.595 0.700 ;
        RECT 73.410 0.260 136.595 0.700 ;
        RECT 73.410 0.255 136.585 0.700 ;
        RECT 73.420 0.250 136.585 0.700 ;
        RECT 73.420 0.245 136.575 0.700 ;
        RECT 73.430 0.240 136.575 0.700 ;
        RECT 73.430 0.235 136.565 0.700 ;
        RECT 73.440 0.230 136.565 0.700 ;
        RECT 73.440 0.225 136.555 0.700 ;
        RECT 73.450 0.220 136.555 0.700 ;
        RECT 73.450 0.215 136.545 0.700 ;
        RECT 73.460 0.210 136.545 0.700 ;
        RECT 73.460 0.205 136.535 0.700 ;
        RECT 73.470 0.200 136.535 0.700 ;
        RECT 73.470 0.195 136.525 0.700 ;
        RECT 73.480 0.190 136.525 0.700 ;
        RECT 73.480 0.185 136.515 0.700 ;
        RECT 73.490 0.180 136.515 0.700 ;
        RECT 73.490 0.175 136.505 0.700 ;
        RECT 73.500 0.170 136.505 0.700 ;
        RECT 73.500 0.165 136.495 0.700 ;
        RECT 73.510 0.160 136.495 0.700 ;
        RECT 73.510 0.155 136.485 0.700 ;
        RECT 73.520 0.150 136.485 0.700 ;
        RECT 73.520 0.145 136.475 0.700 ;
        RECT 73.530 0.140 136.475 0.700 ;
        RECT 73.530 0.135 136.465 0.700 ;
        RECT 73.540 0.130 136.465 0.700 ;
        RECT 73.540 0.125 136.455 0.700 ;
        RECT 73.550 0.120 136.455 0.700 ;
        RECT 73.550 0.115 136.445 0.700 ;
        RECT 73.560 0.110 136.445 0.700 ;
        RECT 73.560 0.105 136.435 0.700 ;
        RECT 73.570 0.100 136.435 0.700 ;
        RECT 73.570 0.095 136.425 0.700 ;
        RECT 73.580 0.090 136.425 0.700 ;
        RECT 73.580 0.085 136.415 0.700 ;
        RECT 73.590 0.080 136.415 0.700 ;
        RECT 73.590 0.075 136.405 0.700 ;
        RECT 73.600 0.070 136.405 0.700 ;
        RECT 73.600 0.065 136.395 0.700 ;
        RECT 73.610 0.060 136.395 0.700 ;
        RECT 73.610 0.055 136.385 0.700 ;
        RECT 73.620 0.050 136.385 0.700 ;
        RECT 73.620 0.045 136.375 0.700 ;
        RECT 73.630 0.040 136.375 0.700 ;
        RECT 73.630 0.035 136.365 0.700 ;
        RECT 73.640 0.030 136.365 0.700 ;
        RECT 73.640 0.025 136.355 0.700 ;
        RECT 73.650 0.020 136.355 0.700 ;
        RECT 73.650 0.015 136.345 0.700 ;
        RECT 73.660 0.010 136.345 0.700 ;
        RECT 73.660 0.005 136.335 0.700 ;
        RECT 73.665 0.000 136.335 0.700 ;
    END
  END XTALOUT
  PIN EO
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 115.610 173.380 116.610 174.000 ;
      LAYER V6 ;
        RECT 115.930 173.510 116.290 173.870 ;
      LAYER M4 ;
        RECT 115.610 173.380 116.610 174.000 ;
      LAYER V3 ;
        RECT 115.810 173.800 116.000 173.990 ;
        RECT 115.810 173.390 116.000 173.580 ;
        RECT 116.220 173.800 116.410 173.990 ;
        RECT 116.220 173.390 116.410 173.580 ;
      LAYER M3 ;
        RECT 115.610 173.380 116.610 174.000 ;
      LAYER V2 ;
        RECT 115.810 173.800 116.000 173.990 ;
        RECT 115.810 173.390 116.000 173.580 ;
        RECT 116.220 173.800 116.410 173.990 ;
        RECT 116.220 173.390 116.410 173.580 ;
      LAYER M2 ;
        RECT 116.010 173.300 116.210 174.000 ;
        RECT 115.610 173.380 116.610 174.000 ;
      LAYER V1 ;
        RECT 115.810 173.800 116.000 173.990 ;
        RECT 115.810 173.390 116.000 173.580 ;
        RECT 116.220 173.800 116.410 173.990 ;
        RECT 116.220 173.390 116.410 173.580 ;
      LAYER M1 ;
        RECT 115.610 173.380 116.610 174.000 ;
      LAYER M6 ;
        RECT 115.610 173.380 116.610 174.000 ;
      LAYER V5 ;
        RECT 115.810 173.800 116.000 173.990 ;
        RECT 115.810 173.390 116.000 173.580 ;
        RECT 116.220 173.800 116.410 173.990 ;
        RECT 116.220 173.390 116.410 173.580 ;
      LAYER M5 ;
        RECT 115.610 173.380 116.610 174.000 ;
      LAYER V4 ;
        RECT 115.810 173.800 116.000 173.990 ;
        RECT 115.810 173.390 116.000 173.580 ;
        RECT 116.220 173.800 116.410 173.990 ;
        RECT 116.220 173.390 116.410 173.580 ;
    END
  END EO
  PIN CK
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 103.755 173.380 104.755 174.000 ;
      LAYER V6 ;
        RECT 104.075 173.510 104.435 173.870 ;
      LAYER M4 ;
        RECT 103.755 173.380 104.755 174.000 ;
      LAYER V3 ;
        RECT 103.955 173.800 104.145 173.990 ;
        RECT 103.955 173.390 104.145 173.580 ;
        RECT 104.365 173.800 104.555 173.990 ;
        RECT 104.365 173.390 104.555 173.580 ;
      LAYER M3 ;
        RECT 103.755 173.380 104.755 174.000 ;
      LAYER V2 ;
        RECT 103.955 173.800 104.145 173.990 ;
        RECT 103.955 173.390 104.145 173.580 ;
        RECT 104.365 173.800 104.555 173.990 ;
        RECT 104.365 173.390 104.555 173.580 ;
      LAYER M2 ;
        RECT 103.755 173.300 104.755 174.000 ;
      LAYER V1 ;
        RECT 103.955 173.800 104.145 173.990 ;
        RECT 103.955 173.390 104.145 173.580 ;
        RECT 104.365 173.800 104.555 173.990 ;
        RECT 104.365 173.390 104.555 173.580 ;
      LAYER M1 ;
        RECT 103.755 173.380 104.755 174.000 ;
      LAYER M6 ;
        RECT 103.755 173.380 104.755 174.000 ;
      LAYER V5 ;
        RECT 103.955 173.800 104.145 173.990 ;
        RECT 103.955 173.390 104.145 173.580 ;
        RECT 104.365 173.800 104.555 173.990 ;
        RECT 104.365 173.390 104.555 173.580 ;
      LAYER M5 ;
        RECT 103.755 173.380 104.755 174.000 ;
      LAYER V4 ;
        RECT 103.955 173.800 104.145 173.990 ;
        RECT 103.955 173.390 104.145 173.580 ;
        RECT 104.365 173.800 104.555 173.990 ;
        RECT 104.365 173.390 104.555 173.580 ;
    END
  END CK
  OBS 
      LAYER M4 ;
        RECT 0.160 156.095 0.700 161.085 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.345 0.700 100.135 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 165.900 172.900 ;
        RECT 166.300 151.245 166.735 153.935 ;
        RECT 166.300 83.165 166.750 88.155 ;
        RECT 166.300 155.725 166.815 161.220 ;
      LAYER M1 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.600 155.725 0.700 165.695 ;
        RECT 0.000 115.135 0.700 151.515 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 165.900 172.900 ;
        RECT 166.300 155.725 167.000 161.220 ;
        RECT 166.300 115.135 167.000 154.220 ;
        RECT 166.300 110.315 167.000 113.895 ;
        RECT 166.300 70.000 167.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 156.095 0.700 161.085 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.345 0.700 100.135 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 165.900 172.900 ;
        RECT 166.300 151.245 166.735 153.935 ;
        RECT 166.300 83.165 166.750 88.155 ;
        RECT 166.300 155.725 166.815 161.220 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 165.900 172.900 ;
        RECT 166.300 171.175 167.000 172.780 ;
        RECT 166.300 162.720 167.000 170.715 ;
        RECT 166.300 155.725 167.000 161.220 ;
        RECT 166.300 150.480 167.000 154.220 ;
        RECT 166.300 137.395 167.000 147.565 ;
        RECT 166.300 127.100 167.000 134.395 ;
        RECT 166.300 121.860 167.000 124.100 ;
        RECT 166.300 115.135 167.000 119.705 ;
        RECT 166.300 110.315 167.000 113.895 ;
        RECT 166.300 97.700 167.000 108.815 ;
        RECT 166.300 86.640 167.000 94.700 ;
        RECT 166.300 75.630 167.000 83.640 ;
        RECT 166.300 70.000 167.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 165.900 172.900 ;
        RECT 166.300 171.175 167.000 172.780 ;
        RECT 166.300 162.720 167.000 170.715 ;
        RECT 166.300 155.725 167.000 161.220 ;
        RECT 166.300 150.480 167.000 154.220 ;
        RECT 166.300 143.340 167.000 147.565 ;
        RECT 166.300 131.850 167.000 140.340 ;
        RECT 166.300 121.860 167.000 128.850 ;
        RECT 166.300 115.135 167.000 119.705 ;
        RECT 166.300 110.315 167.000 113.895 ;
        RECT 166.300 103.280 167.000 108.815 ;
        RECT 166.300 92.280 167.000 100.280 ;
        RECT 166.300 81.280 167.000 89.280 ;
        RECT 166.300 70.000 167.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 165.900 172.900 ;
        RECT 166.300 171.175 167.000 172.780 ;
        RECT 166.300 162.720 167.000 170.715 ;
        RECT 166.300 155.725 167.000 161.220 ;
        RECT 166.300 150.480 167.000 154.220 ;
        RECT 166.300 143.340 167.000 147.565 ;
        RECT 166.300 131.850 167.000 140.340 ;
        RECT 166.300 121.860 167.000 128.850 ;
        RECT 166.300 115.135 167.000 119.705 ;
        RECT 166.300 110.315 167.000 113.895 ;
        RECT 166.300 103.280 167.000 108.815 ;
        RECT 166.300 92.280 167.000 100.280 ;
        RECT 166.300 81.280 167.000 89.280 ;
        RECT 166.300 70.000 167.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 156.095 0.700 161.085 ;
        RECT 0.135 115.870 0.700 154.905 ;
        RECT 0.145 115.860 0.700 154.915 ;
        RECT 0.155 115.850 0.700 154.925 ;
        RECT 0.165 115.840 0.700 154.935 ;
        RECT 0.175 115.830 0.700 154.945 ;
        RECT 0.185 115.820 0.700 154.955 ;
        RECT 0.195 115.810 0.700 154.965 ;
        RECT 0.205 115.800 0.700 154.975 ;
        RECT 0.215 115.790 0.700 154.985 ;
        RECT 0.225 115.780 0.700 154.995 ;
        RECT 0.235 115.770 0.700 155.005 ;
        RECT 0.245 115.760 0.700 155.015 ;
        RECT 0.255 115.750 0.700 155.025 ;
        RECT 0.265 115.740 0.700 155.035 ;
        RECT 0.270 115.735 0.700 155.040 ;
        RECT 0.280 115.735 0.700 155.050 ;
        RECT 0.285 115.735 0.700 155.055 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.345 0.700 100.135 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 165.900 172.900 ;
        RECT 166.300 151.245 166.735 153.935 ;
        RECT 166.300 83.165 166.750 88.155 ;
        RECT 166.300 155.725 166.815 161.220 ;
  END 
END PLOSCR14M

MACRO PLOSC14M
  CLASS  PAD ;
  FOREIGN PLOSC14M 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN XTALIN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
    END
  END XTALIN
  PIN EI
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 63.680 173.380 64.680 174.000 ;
      LAYER V6 ;
        RECT 64.000 173.510 64.360 173.870 ;
      LAYER M4 ;
        RECT 63.680 173.380 64.680 174.000 ;
      LAYER V3 ;
        RECT 63.880 173.800 64.070 173.990 ;
        RECT 63.880 173.390 64.070 173.580 ;
        RECT 64.290 173.800 64.480 173.990 ;
        RECT 64.290 173.390 64.480 173.580 ;
      LAYER M3 ;
        RECT 63.680 173.380 64.680 174.000 ;
      LAYER V2 ;
        RECT 63.880 173.800 64.070 173.990 ;
        RECT 63.880 173.390 64.070 173.580 ;
        RECT 64.290 173.800 64.480 173.990 ;
        RECT 64.290 173.390 64.480 173.580 ;
      LAYER M2 ;
        RECT 64.080 173.300 64.280 174.000 ;
        RECT 63.680 173.380 64.680 174.000 ;
      LAYER V1 ;
        RECT 63.880 173.800 64.070 173.990 ;
        RECT 63.880 173.390 64.070 173.580 ;
        RECT 64.290 173.800 64.480 173.990 ;
        RECT 64.290 173.390 64.480 173.580 ;
      LAYER M1 ;
        RECT 63.680 173.380 64.680 174.000 ;
      LAYER M6 ;
        RECT 63.680 173.380 64.680 174.000 ;
      LAYER V5 ;
        RECT 63.880 173.800 64.070 173.990 ;
        RECT 63.880 173.390 64.070 173.580 ;
        RECT 64.290 173.800 64.480 173.990 ;
        RECT 64.290 173.390 64.480 173.580 ;
      LAYER M5 ;
        RECT 63.680 173.380 64.680 174.000 ;
      LAYER V4 ;
        RECT 63.880 173.800 64.070 173.990 ;
        RECT 63.880 173.390 64.070 173.580 ;
        RECT 64.290 173.800 64.480 173.990 ;
        RECT 64.290 173.390 64.480 173.580 ;
    END
  END EI
  PIN XTALOUT
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 73.000 0.665 137.000 0.700 ;
        RECT 73.010 0.660 136.995 0.700 ;
        RECT 73.010 0.655 136.985 0.700 ;
        RECT 73.020 0.650 136.985 0.700 ;
        RECT 73.020 0.645 136.975 0.700 ;
        RECT 73.030 0.640 136.975 0.700 ;
        RECT 73.030 0.635 136.965 0.700 ;
        RECT 73.040 0.630 136.965 0.700 ;
        RECT 73.040 0.625 136.955 0.700 ;
        RECT 73.050 0.620 136.955 0.700 ;
        RECT 73.050 0.615 136.945 0.700 ;
        RECT 73.060 0.610 136.945 0.700 ;
        RECT 73.060 0.605 136.935 0.700 ;
        RECT 73.070 0.600 136.935 0.700 ;
        RECT 73.070 0.595 136.925 0.700 ;
        RECT 73.080 0.590 136.925 0.700 ;
        RECT 73.080 0.585 136.915 0.700 ;
        RECT 73.090 0.580 136.915 0.700 ;
        RECT 73.090 0.575 136.905 0.700 ;
        RECT 73.100 0.570 136.905 0.700 ;
        RECT 73.100 0.565 136.895 0.700 ;
        RECT 73.110 0.560 136.895 0.700 ;
        RECT 73.110 0.555 136.885 0.700 ;
        RECT 73.120 0.550 136.885 0.700 ;
        RECT 73.120 0.545 136.875 0.700 ;
        RECT 73.130 0.540 136.875 0.700 ;
        RECT 73.130 0.535 136.865 0.700 ;
        RECT 73.140 0.530 136.865 0.700 ;
        RECT 73.140 0.525 136.855 0.700 ;
        RECT 73.150 0.520 136.855 0.700 ;
        RECT 73.150 0.515 136.845 0.700 ;
        RECT 73.160 0.510 136.845 0.700 ;
        RECT 73.160 0.505 136.835 0.700 ;
        RECT 73.170 0.500 136.835 0.700 ;
        RECT 73.170 0.495 136.825 0.700 ;
        RECT 73.180 0.490 136.825 0.700 ;
        RECT 73.180 0.485 136.815 0.700 ;
        RECT 73.190 0.480 136.815 0.700 ;
        RECT 73.190 0.475 136.805 0.700 ;
        RECT 73.200 0.470 136.805 0.700 ;
        RECT 73.200 0.465 136.795 0.700 ;
        RECT 73.210 0.460 136.795 0.700 ;
        RECT 73.210 0.455 136.785 0.700 ;
        RECT 73.220 0.450 136.785 0.700 ;
        RECT 73.220 0.445 136.775 0.700 ;
        RECT 73.230 0.440 136.775 0.700 ;
        RECT 73.230 0.435 136.765 0.700 ;
        RECT 73.240 0.430 136.765 0.700 ;
        RECT 73.240 0.425 136.755 0.700 ;
        RECT 73.250 0.420 136.755 0.700 ;
        RECT 73.250 0.415 136.745 0.700 ;
        RECT 73.260 0.410 136.745 0.700 ;
        RECT 73.260 0.405 136.735 0.700 ;
        RECT 73.270 0.400 136.735 0.700 ;
        RECT 73.270 0.395 136.725 0.700 ;
        RECT 73.280 0.390 136.725 0.700 ;
        RECT 73.280 0.385 136.715 0.700 ;
        RECT 73.290 0.380 136.715 0.700 ;
        RECT 73.290 0.375 136.705 0.700 ;
        RECT 73.300 0.370 136.705 0.700 ;
        RECT 73.300 0.365 136.695 0.700 ;
        RECT 73.310 0.360 136.695 0.700 ;
        RECT 73.310 0.355 136.685 0.700 ;
        RECT 73.320 0.350 136.685 0.700 ;
        RECT 73.320 0.345 136.675 0.700 ;
        RECT 73.330 0.340 136.675 0.700 ;
        RECT 73.330 0.335 136.665 0.700 ;
        RECT 73.340 0.330 136.665 0.700 ;
        RECT 73.340 0.325 136.655 0.700 ;
        RECT 73.350 0.320 136.655 0.700 ;
        RECT 73.350 0.315 136.645 0.700 ;
        RECT 73.360 0.310 136.645 0.700 ;
        RECT 73.360 0.305 136.635 0.700 ;
        RECT 73.370 0.300 136.635 0.700 ;
        RECT 73.370 0.295 136.625 0.700 ;
        RECT 73.380 0.290 136.625 0.700 ;
        RECT 73.380 0.285 136.615 0.700 ;
        RECT 73.390 0.280 136.615 0.700 ;
        RECT 73.390 0.275 136.605 0.700 ;
        RECT 73.400 0.270 136.605 0.700 ;
        RECT 73.400 0.265 136.595 0.700 ;
        RECT 73.410 0.260 136.595 0.700 ;
        RECT 73.410 0.255 136.585 0.700 ;
        RECT 73.420 0.250 136.585 0.700 ;
        RECT 73.420 0.245 136.575 0.700 ;
        RECT 73.430 0.240 136.575 0.700 ;
        RECT 73.430 0.235 136.565 0.700 ;
        RECT 73.440 0.230 136.565 0.700 ;
        RECT 73.440 0.225 136.555 0.700 ;
        RECT 73.450 0.220 136.555 0.700 ;
        RECT 73.450 0.215 136.545 0.700 ;
        RECT 73.460 0.210 136.545 0.700 ;
        RECT 73.460 0.205 136.535 0.700 ;
        RECT 73.470 0.200 136.535 0.700 ;
        RECT 73.470 0.195 136.525 0.700 ;
        RECT 73.480 0.190 136.525 0.700 ;
        RECT 73.480 0.185 136.515 0.700 ;
        RECT 73.490 0.180 136.515 0.700 ;
        RECT 73.490 0.175 136.505 0.700 ;
        RECT 73.500 0.170 136.505 0.700 ;
        RECT 73.500 0.165 136.495 0.700 ;
        RECT 73.510 0.160 136.495 0.700 ;
        RECT 73.510 0.155 136.485 0.700 ;
        RECT 73.520 0.150 136.485 0.700 ;
        RECT 73.520 0.145 136.475 0.700 ;
        RECT 73.530 0.140 136.475 0.700 ;
        RECT 73.530 0.135 136.465 0.700 ;
        RECT 73.540 0.130 136.465 0.700 ;
        RECT 73.540 0.125 136.455 0.700 ;
        RECT 73.550 0.120 136.455 0.700 ;
        RECT 73.550 0.115 136.445 0.700 ;
        RECT 73.560 0.110 136.445 0.700 ;
        RECT 73.560 0.105 136.435 0.700 ;
        RECT 73.570 0.100 136.435 0.700 ;
        RECT 73.570 0.095 136.425 0.700 ;
        RECT 73.580 0.090 136.425 0.700 ;
        RECT 73.580 0.085 136.415 0.700 ;
        RECT 73.590 0.080 136.415 0.700 ;
        RECT 73.590 0.075 136.405 0.700 ;
        RECT 73.600 0.070 136.405 0.700 ;
        RECT 73.600 0.065 136.395 0.700 ;
        RECT 73.610 0.060 136.395 0.700 ;
        RECT 73.610 0.055 136.385 0.700 ;
        RECT 73.620 0.050 136.385 0.700 ;
        RECT 73.620 0.045 136.375 0.700 ;
        RECT 73.630 0.040 136.375 0.700 ;
        RECT 73.630 0.035 136.365 0.700 ;
        RECT 73.640 0.030 136.365 0.700 ;
        RECT 73.640 0.025 136.355 0.700 ;
        RECT 73.650 0.020 136.355 0.700 ;
        RECT 73.650 0.015 136.345 0.700 ;
        RECT 73.660 0.010 136.345 0.700 ;
        RECT 73.660 0.005 136.335 0.700 ;
        RECT 73.665 0.000 136.335 0.700 ;
      LAYER M4 ;
        RECT 73.000 0.665 137.000 0.700 ;
        RECT 73.010 0.660 136.995 0.700 ;
        RECT 73.010 0.655 136.985 0.700 ;
        RECT 73.020 0.650 136.985 0.700 ;
        RECT 73.020 0.645 136.975 0.700 ;
        RECT 73.030 0.640 136.975 0.700 ;
        RECT 73.030 0.635 136.965 0.700 ;
        RECT 73.040 0.630 136.965 0.700 ;
        RECT 73.040 0.625 136.955 0.700 ;
        RECT 73.050 0.620 136.955 0.700 ;
        RECT 73.050 0.615 136.945 0.700 ;
        RECT 73.060 0.610 136.945 0.700 ;
        RECT 73.060 0.605 136.935 0.700 ;
        RECT 73.070 0.600 136.935 0.700 ;
        RECT 73.070 0.595 136.925 0.700 ;
        RECT 73.080 0.590 136.925 0.700 ;
        RECT 73.080 0.585 136.915 0.700 ;
        RECT 73.090 0.580 136.915 0.700 ;
        RECT 73.090 0.575 136.905 0.700 ;
        RECT 73.100 0.570 136.905 0.700 ;
        RECT 73.100 0.565 136.895 0.700 ;
        RECT 73.110 0.560 136.895 0.700 ;
        RECT 73.110 0.555 136.885 0.700 ;
        RECT 73.120 0.550 136.885 0.700 ;
        RECT 73.120 0.545 136.875 0.700 ;
        RECT 73.130 0.540 136.875 0.700 ;
        RECT 73.130 0.535 136.865 0.700 ;
        RECT 73.140 0.530 136.865 0.700 ;
        RECT 73.140 0.525 136.855 0.700 ;
        RECT 73.150 0.520 136.855 0.700 ;
        RECT 73.150 0.515 136.845 0.700 ;
        RECT 73.160 0.510 136.845 0.700 ;
        RECT 73.160 0.505 136.835 0.700 ;
        RECT 73.170 0.500 136.835 0.700 ;
        RECT 73.170 0.495 136.825 0.700 ;
        RECT 73.180 0.490 136.825 0.700 ;
        RECT 73.180 0.485 136.815 0.700 ;
        RECT 73.190 0.480 136.815 0.700 ;
        RECT 73.190 0.475 136.805 0.700 ;
        RECT 73.200 0.470 136.805 0.700 ;
        RECT 73.200 0.465 136.795 0.700 ;
        RECT 73.210 0.460 136.795 0.700 ;
        RECT 73.210 0.455 136.785 0.700 ;
        RECT 73.220 0.450 136.785 0.700 ;
        RECT 73.220 0.445 136.775 0.700 ;
        RECT 73.230 0.440 136.775 0.700 ;
        RECT 73.230 0.435 136.765 0.700 ;
        RECT 73.240 0.430 136.765 0.700 ;
        RECT 73.240 0.425 136.755 0.700 ;
        RECT 73.250 0.420 136.755 0.700 ;
        RECT 73.250 0.415 136.745 0.700 ;
        RECT 73.260 0.410 136.745 0.700 ;
        RECT 73.260 0.405 136.735 0.700 ;
        RECT 73.270 0.400 136.735 0.700 ;
        RECT 73.270 0.395 136.725 0.700 ;
        RECT 73.280 0.390 136.725 0.700 ;
        RECT 73.280 0.385 136.715 0.700 ;
        RECT 73.290 0.380 136.715 0.700 ;
        RECT 73.290 0.375 136.705 0.700 ;
        RECT 73.300 0.370 136.705 0.700 ;
        RECT 73.300 0.365 136.695 0.700 ;
        RECT 73.310 0.360 136.695 0.700 ;
        RECT 73.310 0.355 136.685 0.700 ;
        RECT 73.320 0.350 136.685 0.700 ;
        RECT 73.320 0.345 136.675 0.700 ;
        RECT 73.330 0.340 136.675 0.700 ;
        RECT 73.330 0.335 136.665 0.700 ;
        RECT 73.340 0.330 136.665 0.700 ;
        RECT 73.340 0.325 136.655 0.700 ;
        RECT 73.350 0.320 136.655 0.700 ;
        RECT 73.350 0.315 136.645 0.700 ;
        RECT 73.360 0.310 136.645 0.700 ;
        RECT 73.360 0.305 136.635 0.700 ;
        RECT 73.370 0.300 136.635 0.700 ;
        RECT 73.370 0.295 136.625 0.700 ;
        RECT 73.380 0.290 136.625 0.700 ;
        RECT 73.380 0.285 136.615 0.700 ;
        RECT 73.390 0.280 136.615 0.700 ;
        RECT 73.390 0.275 136.605 0.700 ;
        RECT 73.400 0.270 136.605 0.700 ;
        RECT 73.400 0.265 136.595 0.700 ;
        RECT 73.410 0.260 136.595 0.700 ;
        RECT 73.410 0.255 136.585 0.700 ;
        RECT 73.420 0.250 136.585 0.700 ;
        RECT 73.420 0.245 136.575 0.700 ;
        RECT 73.430 0.240 136.575 0.700 ;
        RECT 73.430 0.235 136.565 0.700 ;
        RECT 73.440 0.230 136.565 0.700 ;
        RECT 73.440 0.225 136.555 0.700 ;
        RECT 73.450 0.220 136.555 0.700 ;
        RECT 73.450 0.215 136.545 0.700 ;
        RECT 73.460 0.210 136.545 0.700 ;
        RECT 73.460 0.205 136.535 0.700 ;
        RECT 73.470 0.200 136.535 0.700 ;
        RECT 73.470 0.195 136.525 0.700 ;
        RECT 73.480 0.190 136.525 0.700 ;
        RECT 73.480 0.185 136.515 0.700 ;
        RECT 73.490 0.180 136.515 0.700 ;
        RECT 73.490 0.175 136.505 0.700 ;
        RECT 73.500 0.170 136.505 0.700 ;
        RECT 73.500 0.165 136.495 0.700 ;
        RECT 73.510 0.160 136.495 0.700 ;
        RECT 73.510 0.155 136.485 0.700 ;
        RECT 73.520 0.150 136.485 0.700 ;
        RECT 73.520 0.145 136.475 0.700 ;
        RECT 73.530 0.140 136.475 0.700 ;
        RECT 73.530 0.135 136.465 0.700 ;
        RECT 73.540 0.130 136.465 0.700 ;
        RECT 73.540 0.125 136.455 0.700 ;
        RECT 73.550 0.120 136.455 0.700 ;
        RECT 73.550 0.115 136.445 0.700 ;
        RECT 73.560 0.110 136.445 0.700 ;
        RECT 73.560 0.105 136.435 0.700 ;
        RECT 73.570 0.100 136.435 0.700 ;
        RECT 73.570 0.095 136.425 0.700 ;
        RECT 73.580 0.090 136.425 0.700 ;
        RECT 73.580 0.085 136.415 0.700 ;
        RECT 73.590 0.080 136.415 0.700 ;
        RECT 73.590 0.075 136.405 0.700 ;
        RECT 73.600 0.070 136.405 0.700 ;
        RECT 73.600 0.065 136.395 0.700 ;
        RECT 73.610 0.060 136.395 0.700 ;
        RECT 73.610 0.055 136.385 0.700 ;
        RECT 73.620 0.050 136.385 0.700 ;
        RECT 73.620 0.045 136.375 0.700 ;
        RECT 73.630 0.040 136.375 0.700 ;
        RECT 73.630 0.035 136.365 0.700 ;
        RECT 73.640 0.030 136.365 0.700 ;
        RECT 73.640 0.025 136.355 0.700 ;
        RECT 73.650 0.020 136.355 0.700 ;
        RECT 73.650 0.015 136.345 0.700 ;
        RECT 73.660 0.010 136.345 0.700 ;
        RECT 73.660 0.005 136.335 0.700 ;
        RECT 73.665 0.000 136.335 0.700 ;
      LAYER M3 ;
        RECT 73.000 0.665 137.000 0.700 ;
        RECT 73.010 0.660 136.995 0.700 ;
        RECT 73.010 0.655 136.985 0.700 ;
        RECT 73.020 0.650 136.985 0.700 ;
        RECT 73.020 0.645 136.975 0.700 ;
        RECT 73.030 0.640 136.975 0.700 ;
        RECT 73.030 0.635 136.965 0.700 ;
        RECT 73.040 0.630 136.965 0.700 ;
        RECT 73.040 0.625 136.955 0.700 ;
        RECT 73.050 0.620 136.955 0.700 ;
        RECT 73.050 0.615 136.945 0.700 ;
        RECT 73.060 0.610 136.945 0.700 ;
        RECT 73.060 0.605 136.935 0.700 ;
        RECT 73.070 0.600 136.935 0.700 ;
        RECT 73.070 0.595 136.925 0.700 ;
        RECT 73.080 0.590 136.925 0.700 ;
        RECT 73.080 0.585 136.915 0.700 ;
        RECT 73.090 0.580 136.915 0.700 ;
        RECT 73.090 0.575 136.905 0.700 ;
        RECT 73.100 0.570 136.905 0.700 ;
        RECT 73.100 0.565 136.895 0.700 ;
        RECT 73.110 0.560 136.895 0.700 ;
        RECT 73.110 0.555 136.885 0.700 ;
        RECT 73.120 0.550 136.885 0.700 ;
        RECT 73.120 0.545 136.875 0.700 ;
        RECT 73.130 0.540 136.875 0.700 ;
        RECT 73.130 0.535 136.865 0.700 ;
        RECT 73.140 0.530 136.865 0.700 ;
        RECT 73.140 0.525 136.855 0.700 ;
        RECT 73.150 0.520 136.855 0.700 ;
        RECT 73.150 0.515 136.845 0.700 ;
        RECT 73.160 0.510 136.845 0.700 ;
        RECT 73.160 0.505 136.835 0.700 ;
        RECT 73.170 0.500 136.835 0.700 ;
        RECT 73.170 0.495 136.825 0.700 ;
        RECT 73.180 0.490 136.825 0.700 ;
        RECT 73.180 0.485 136.815 0.700 ;
        RECT 73.190 0.480 136.815 0.700 ;
        RECT 73.190 0.475 136.805 0.700 ;
        RECT 73.200 0.470 136.805 0.700 ;
        RECT 73.200 0.465 136.795 0.700 ;
        RECT 73.210 0.460 136.795 0.700 ;
        RECT 73.210 0.455 136.785 0.700 ;
        RECT 73.220 0.450 136.785 0.700 ;
        RECT 73.220 0.445 136.775 0.700 ;
        RECT 73.230 0.440 136.775 0.700 ;
        RECT 73.230 0.435 136.765 0.700 ;
        RECT 73.240 0.430 136.765 0.700 ;
        RECT 73.240 0.425 136.755 0.700 ;
        RECT 73.250 0.420 136.755 0.700 ;
        RECT 73.250 0.415 136.745 0.700 ;
        RECT 73.260 0.410 136.745 0.700 ;
        RECT 73.260 0.405 136.735 0.700 ;
        RECT 73.270 0.400 136.735 0.700 ;
        RECT 73.270 0.395 136.725 0.700 ;
        RECT 73.280 0.390 136.725 0.700 ;
        RECT 73.280 0.385 136.715 0.700 ;
        RECT 73.290 0.380 136.715 0.700 ;
        RECT 73.290 0.375 136.705 0.700 ;
        RECT 73.300 0.370 136.705 0.700 ;
        RECT 73.300 0.365 136.695 0.700 ;
        RECT 73.310 0.360 136.695 0.700 ;
        RECT 73.310 0.355 136.685 0.700 ;
        RECT 73.320 0.350 136.685 0.700 ;
        RECT 73.320 0.345 136.675 0.700 ;
        RECT 73.330 0.340 136.675 0.700 ;
        RECT 73.330 0.335 136.665 0.700 ;
        RECT 73.340 0.330 136.665 0.700 ;
        RECT 73.340 0.325 136.655 0.700 ;
        RECT 73.350 0.320 136.655 0.700 ;
        RECT 73.350 0.315 136.645 0.700 ;
        RECT 73.360 0.310 136.645 0.700 ;
        RECT 73.360 0.305 136.635 0.700 ;
        RECT 73.370 0.300 136.635 0.700 ;
        RECT 73.370 0.295 136.625 0.700 ;
        RECT 73.380 0.290 136.625 0.700 ;
        RECT 73.380 0.285 136.615 0.700 ;
        RECT 73.390 0.280 136.615 0.700 ;
        RECT 73.390 0.275 136.605 0.700 ;
        RECT 73.400 0.270 136.605 0.700 ;
        RECT 73.400 0.265 136.595 0.700 ;
        RECT 73.410 0.260 136.595 0.700 ;
        RECT 73.410 0.255 136.585 0.700 ;
        RECT 73.420 0.250 136.585 0.700 ;
        RECT 73.420 0.245 136.575 0.700 ;
        RECT 73.430 0.240 136.575 0.700 ;
        RECT 73.430 0.235 136.565 0.700 ;
        RECT 73.440 0.230 136.565 0.700 ;
        RECT 73.440 0.225 136.555 0.700 ;
        RECT 73.450 0.220 136.555 0.700 ;
        RECT 73.450 0.215 136.545 0.700 ;
        RECT 73.460 0.210 136.545 0.700 ;
        RECT 73.460 0.205 136.535 0.700 ;
        RECT 73.470 0.200 136.535 0.700 ;
        RECT 73.470 0.195 136.525 0.700 ;
        RECT 73.480 0.190 136.525 0.700 ;
        RECT 73.480 0.185 136.515 0.700 ;
        RECT 73.490 0.180 136.515 0.700 ;
        RECT 73.490 0.175 136.505 0.700 ;
        RECT 73.500 0.170 136.505 0.700 ;
        RECT 73.500 0.165 136.495 0.700 ;
        RECT 73.510 0.160 136.495 0.700 ;
        RECT 73.510 0.155 136.485 0.700 ;
        RECT 73.520 0.150 136.485 0.700 ;
        RECT 73.520 0.145 136.475 0.700 ;
        RECT 73.530 0.140 136.475 0.700 ;
        RECT 73.530 0.135 136.465 0.700 ;
        RECT 73.540 0.130 136.465 0.700 ;
        RECT 73.540 0.125 136.455 0.700 ;
        RECT 73.550 0.120 136.455 0.700 ;
        RECT 73.550 0.115 136.445 0.700 ;
        RECT 73.560 0.110 136.445 0.700 ;
        RECT 73.560 0.105 136.435 0.700 ;
        RECT 73.570 0.100 136.435 0.700 ;
        RECT 73.570 0.095 136.425 0.700 ;
        RECT 73.580 0.090 136.425 0.700 ;
        RECT 73.580 0.085 136.415 0.700 ;
        RECT 73.590 0.080 136.415 0.700 ;
        RECT 73.590 0.075 136.405 0.700 ;
        RECT 73.600 0.070 136.405 0.700 ;
        RECT 73.600 0.065 136.395 0.700 ;
        RECT 73.610 0.060 136.395 0.700 ;
        RECT 73.610 0.055 136.385 0.700 ;
        RECT 73.620 0.050 136.385 0.700 ;
        RECT 73.620 0.045 136.375 0.700 ;
        RECT 73.630 0.040 136.375 0.700 ;
        RECT 73.630 0.035 136.365 0.700 ;
        RECT 73.640 0.030 136.365 0.700 ;
        RECT 73.640 0.025 136.355 0.700 ;
        RECT 73.650 0.020 136.355 0.700 ;
        RECT 73.650 0.015 136.345 0.700 ;
        RECT 73.660 0.010 136.345 0.700 ;
        RECT 73.660 0.005 136.335 0.700 ;
        RECT 73.665 0.000 136.335 0.700 ;
      LAYER M2 ;
        RECT 73.000 0.665 137.000 0.700 ;
        RECT 73.010 0.660 136.995 0.700 ;
        RECT 73.010 0.655 136.985 0.700 ;
        RECT 73.020 0.650 136.985 0.700 ;
        RECT 73.020 0.645 136.975 0.700 ;
        RECT 73.030 0.640 136.975 0.700 ;
        RECT 73.030 0.635 136.965 0.700 ;
        RECT 73.040 0.630 136.965 0.700 ;
        RECT 73.040 0.625 136.955 0.700 ;
        RECT 73.050 0.620 136.955 0.700 ;
        RECT 73.050 0.615 136.945 0.700 ;
        RECT 73.060 0.610 136.945 0.700 ;
        RECT 73.060 0.605 136.935 0.700 ;
        RECT 73.070 0.600 136.935 0.700 ;
        RECT 73.070 0.595 136.925 0.700 ;
        RECT 73.080 0.590 136.925 0.700 ;
        RECT 73.080 0.585 136.915 0.700 ;
        RECT 73.090 0.580 136.915 0.700 ;
        RECT 73.090 0.575 136.905 0.700 ;
        RECT 73.100 0.570 136.905 0.700 ;
        RECT 73.100 0.565 136.895 0.700 ;
        RECT 73.110 0.560 136.895 0.700 ;
        RECT 73.110 0.555 136.885 0.700 ;
        RECT 73.120 0.550 136.885 0.700 ;
        RECT 73.120 0.545 136.875 0.700 ;
        RECT 73.130 0.540 136.875 0.700 ;
        RECT 73.130 0.535 136.865 0.700 ;
        RECT 73.140 0.530 136.865 0.700 ;
        RECT 73.140 0.525 136.855 0.700 ;
        RECT 73.150 0.520 136.855 0.700 ;
        RECT 73.150 0.515 136.845 0.700 ;
        RECT 73.160 0.510 136.845 0.700 ;
        RECT 73.160 0.505 136.835 0.700 ;
        RECT 73.170 0.500 136.835 0.700 ;
        RECT 73.170 0.495 136.825 0.700 ;
        RECT 73.180 0.490 136.825 0.700 ;
        RECT 73.180 0.485 136.815 0.700 ;
        RECT 73.190 0.480 136.815 0.700 ;
        RECT 73.190 0.475 136.805 0.700 ;
        RECT 73.200 0.470 136.805 0.700 ;
        RECT 73.200 0.465 136.795 0.700 ;
        RECT 73.210 0.460 136.795 0.700 ;
        RECT 73.210 0.455 136.785 0.700 ;
        RECT 73.220 0.450 136.785 0.700 ;
        RECT 73.220 0.445 136.775 0.700 ;
        RECT 73.230 0.440 136.775 0.700 ;
        RECT 73.230 0.435 136.765 0.700 ;
        RECT 73.240 0.430 136.765 0.700 ;
        RECT 73.240 0.425 136.755 0.700 ;
        RECT 73.250 0.420 136.755 0.700 ;
        RECT 73.250 0.415 136.745 0.700 ;
        RECT 73.260 0.410 136.745 0.700 ;
        RECT 73.260 0.405 136.735 0.700 ;
        RECT 73.270 0.400 136.735 0.700 ;
        RECT 73.270 0.395 136.725 0.700 ;
        RECT 73.280 0.390 136.725 0.700 ;
        RECT 73.280 0.385 136.715 0.700 ;
        RECT 73.290 0.380 136.715 0.700 ;
        RECT 73.290 0.375 136.705 0.700 ;
        RECT 73.300 0.370 136.705 0.700 ;
        RECT 73.300 0.365 136.695 0.700 ;
        RECT 73.310 0.360 136.695 0.700 ;
        RECT 73.310 0.355 136.685 0.700 ;
        RECT 73.320 0.350 136.685 0.700 ;
        RECT 73.320 0.345 136.675 0.700 ;
        RECT 73.330 0.340 136.675 0.700 ;
        RECT 73.330 0.335 136.665 0.700 ;
        RECT 73.340 0.330 136.665 0.700 ;
        RECT 73.340 0.325 136.655 0.700 ;
        RECT 73.350 0.320 136.655 0.700 ;
        RECT 73.350 0.315 136.645 0.700 ;
        RECT 73.360 0.310 136.645 0.700 ;
        RECT 73.360 0.305 136.635 0.700 ;
        RECT 73.370 0.300 136.635 0.700 ;
        RECT 73.370 0.295 136.625 0.700 ;
        RECT 73.380 0.290 136.625 0.700 ;
        RECT 73.380 0.285 136.615 0.700 ;
        RECT 73.390 0.280 136.615 0.700 ;
        RECT 73.390 0.275 136.605 0.700 ;
        RECT 73.400 0.270 136.605 0.700 ;
        RECT 73.400 0.265 136.595 0.700 ;
        RECT 73.410 0.260 136.595 0.700 ;
        RECT 73.410 0.255 136.585 0.700 ;
        RECT 73.420 0.250 136.585 0.700 ;
        RECT 73.420 0.245 136.575 0.700 ;
        RECT 73.430 0.240 136.575 0.700 ;
        RECT 73.430 0.235 136.565 0.700 ;
        RECT 73.440 0.230 136.565 0.700 ;
        RECT 73.440 0.225 136.555 0.700 ;
        RECT 73.450 0.220 136.555 0.700 ;
        RECT 73.450 0.215 136.545 0.700 ;
        RECT 73.460 0.210 136.545 0.700 ;
        RECT 73.460 0.205 136.535 0.700 ;
        RECT 73.470 0.200 136.535 0.700 ;
        RECT 73.470 0.195 136.525 0.700 ;
        RECT 73.480 0.190 136.525 0.700 ;
        RECT 73.480 0.185 136.515 0.700 ;
        RECT 73.490 0.180 136.515 0.700 ;
        RECT 73.490 0.175 136.505 0.700 ;
        RECT 73.500 0.170 136.505 0.700 ;
        RECT 73.500 0.165 136.495 0.700 ;
        RECT 73.510 0.160 136.495 0.700 ;
        RECT 73.510 0.155 136.485 0.700 ;
        RECT 73.520 0.150 136.485 0.700 ;
        RECT 73.520 0.145 136.475 0.700 ;
        RECT 73.530 0.140 136.475 0.700 ;
        RECT 73.530 0.135 136.465 0.700 ;
        RECT 73.540 0.130 136.465 0.700 ;
        RECT 73.540 0.125 136.455 0.700 ;
        RECT 73.550 0.120 136.455 0.700 ;
        RECT 73.550 0.115 136.445 0.700 ;
        RECT 73.560 0.110 136.445 0.700 ;
        RECT 73.560 0.105 136.435 0.700 ;
        RECT 73.570 0.100 136.435 0.700 ;
        RECT 73.570 0.095 136.425 0.700 ;
        RECT 73.580 0.090 136.425 0.700 ;
        RECT 73.580 0.085 136.415 0.700 ;
        RECT 73.590 0.080 136.415 0.700 ;
        RECT 73.590 0.075 136.405 0.700 ;
        RECT 73.600 0.070 136.405 0.700 ;
        RECT 73.600 0.065 136.395 0.700 ;
        RECT 73.610 0.060 136.395 0.700 ;
        RECT 73.610 0.055 136.385 0.700 ;
        RECT 73.620 0.050 136.385 0.700 ;
        RECT 73.620 0.045 136.375 0.700 ;
        RECT 73.630 0.040 136.375 0.700 ;
        RECT 73.630 0.035 136.365 0.700 ;
        RECT 73.640 0.030 136.365 0.700 ;
        RECT 73.640 0.025 136.355 0.700 ;
        RECT 73.650 0.020 136.355 0.700 ;
        RECT 73.650 0.015 136.345 0.700 ;
        RECT 73.660 0.010 136.345 0.700 ;
        RECT 73.660 0.005 136.335 0.700 ;
        RECT 73.665 0.000 136.335 0.700 ;
      LAYER M6 ;
        RECT 73.000 0.665 137.000 0.700 ;
        RECT 73.010 0.660 136.995 0.700 ;
        RECT 73.010 0.655 136.985 0.700 ;
        RECT 73.020 0.650 136.985 0.700 ;
        RECT 73.020 0.645 136.975 0.700 ;
        RECT 73.030 0.640 136.975 0.700 ;
        RECT 73.030 0.635 136.965 0.700 ;
        RECT 73.040 0.630 136.965 0.700 ;
        RECT 73.040 0.625 136.955 0.700 ;
        RECT 73.050 0.620 136.955 0.700 ;
        RECT 73.050 0.615 136.945 0.700 ;
        RECT 73.060 0.610 136.945 0.700 ;
        RECT 73.060 0.605 136.935 0.700 ;
        RECT 73.070 0.600 136.935 0.700 ;
        RECT 73.070 0.595 136.925 0.700 ;
        RECT 73.080 0.590 136.925 0.700 ;
        RECT 73.080 0.585 136.915 0.700 ;
        RECT 73.090 0.580 136.915 0.700 ;
        RECT 73.090 0.575 136.905 0.700 ;
        RECT 73.100 0.570 136.905 0.700 ;
        RECT 73.100 0.565 136.895 0.700 ;
        RECT 73.110 0.560 136.895 0.700 ;
        RECT 73.110 0.555 136.885 0.700 ;
        RECT 73.120 0.550 136.885 0.700 ;
        RECT 73.120 0.545 136.875 0.700 ;
        RECT 73.130 0.540 136.875 0.700 ;
        RECT 73.130 0.535 136.865 0.700 ;
        RECT 73.140 0.530 136.865 0.700 ;
        RECT 73.140 0.525 136.855 0.700 ;
        RECT 73.150 0.520 136.855 0.700 ;
        RECT 73.150 0.515 136.845 0.700 ;
        RECT 73.160 0.510 136.845 0.700 ;
        RECT 73.160 0.505 136.835 0.700 ;
        RECT 73.170 0.500 136.835 0.700 ;
        RECT 73.170 0.495 136.825 0.700 ;
        RECT 73.180 0.490 136.825 0.700 ;
        RECT 73.180 0.485 136.815 0.700 ;
        RECT 73.190 0.480 136.815 0.700 ;
        RECT 73.190 0.475 136.805 0.700 ;
        RECT 73.200 0.470 136.805 0.700 ;
        RECT 73.200 0.465 136.795 0.700 ;
        RECT 73.210 0.460 136.795 0.700 ;
        RECT 73.210 0.455 136.785 0.700 ;
        RECT 73.220 0.450 136.785 0.700 ;
        RECT 73.220 0.445 136.775 0.700 ;
        RECT 73.230 0.440 136.775 0.700 ;
        RECT 73.230 0.435 136.765 0.700 ;
        RECT 73.240 0.430 136.765 0.700 ;
        RECT 73.240 0.425 136.755 0.700 ;
        RECT 73.250 0.420 136.755 0.700 ;
        RECT 73.250 0.415 136.745 0.700 ;
        RECT 73.260 0.410 136.745 0.700 ;
        RECT 73.260 0.405 136.735 0.700 ;
        RECT 73.270 0.400 136.735 0.700 ;
        RECT 73.270 0.395 136.725 0.700 ;
        RECT 73.280 0.390 136.725 0.700 ;
        RECT 73.280 0.385 136.715 0.700 ;
        RECT 73.290 0.380 136.715 0.700 ;
        RECT 73.290 0.375 136.705 0.700 ;
        RECT 73.300 0.370 136.705 0.700 ;
        RECT 73.300 0.365 136.695 0.700 ;
        RECT 73.310 0.360 136.695 0.700 ;
        RECT 73.310 0.355 136.685 0.700 ;
        RECT 73.320 0.350 136.685 0.700 ;
        RECT 73.320 0.345 136.675 0.700 ;
        RECT 73.330 0.340 136.675 0.700 ;
        RECT 73.330 0.335 136.665 0.700 ;
        RECT 73.340 0.330 136.665 0.700 ;
        RECT 73.340 0.325 136.655 0.700 ;
        RECT 73.350 0.320 136.655 0.700 ;
        RECT 73.350 0.315 136.645 0.700 ;
        RECT 73.360 0.310 136.645 0.700 ;
        RECT 73.360 0.305 136.635 0.700 ;
        RECT 73.370 0.300 136.635 0.700 ;
        RECT 73.370 0.295 136.625 0.700 ;
        RECT 73.380 0.290 136.625 0.700 ;
        RECT 73.380 0.285 136.615 0.700 ;
        RECT 73.390 0.280 136.615 0.700 ;
        RECT 73.390 0.275 136.605 0.700 ;
        RECT 73.400 0.270 136.605 0.700 ;
        RECT 73.400 0.265 136.595 0.700 ;
        RECT 73.410 0.260 136.595 0.700 ;
        RECT 73.410 0.255 136.585 0.700 ;
        RECT 73.420 0.250 136.585 0.700 ;
        RECT 73.420 0.245 136.575 0.700 ;
        RECT 73.430 0.240 136.575 0.700 ;
        RECT 73.430 0.235 136.565 0.700 ;
        RECT 73.440 0.230 136.565 0.700 ;
        RECT 73.440 0.225 136.555 0.700 ;
        RECT 73.450 0.220 136.555 0.700 ;
        RECT 73.450 0.215 136.545 0.700 ;
        RECT 73.460 0.210 136.545 0.700 ;
        RECT 73.460 0.205 136.535 0.700 ;
        RECT 73.470 0.200 136.535 0.700 ;
        RECT 73.470 0.195 136.525 0.700 ;
        RECT 73.480 0.190 136.525 0.700 ;
        RECT 73.480 0.185 136.515 0.700 ;
        RECT 73.490 0.180 136.515 0.700 ;
        RECT 73.490 0.175 136.505 0.700 ;
        RECT 73.500 0.170 136.505 0.700 ;
        RECT 73.500 0.165 136.495 0.700 ;
        RECT 73.510 0.160 136.495 0.700 ;
        RECT 73.510 0.155 136.485 0.700 ;
        RECT 73.520 0.150 136.485 0.700 ;
        RECT 73.520 0.145 136.475 0.700 ;
        RECT 73.530 0.140 136.475 0.700 ;
        RECT 73.530 0.135 136.465 0.700 ;
        RECT 73.540 0.130 136.465 0.700 ;
        RECT 73.540 0.125 136.455 0.700 ;
        RECT 73.550 0.120 136.455 0.700 ;
        RECT 73.550 0.115 136.445 0.700 ;
        RECT 73.560 0.110 136.445 0.700 ;
        RECT 73.560 0.105 136.435 0.700 ;
        RECT 73.570 0.100 136.435 0.700 ;
        RECT 73.570 0.095 136.425 0.700 ;
        RECT 73.580 0.090 136.425 0.700 ;
        RECT 73.580 0.085 136.415 0.700 ;
        RECT 73.590 0.080 136.415 0.700 ;
        RECT 73.590 0.075 136.405 0.700 ;
        RECT 73.600 0.070 136.405 0.700 ;
        RECT 73.600 0.065 136.395 0.700 ;
        RECT 73.610 0.060 136.395 0.700 ;
        RECT 73.610 0.055 136.385 0.700 ;
        RECT 73.620 0.050 136.385 0.700 ;
        RECT 73.620 0.045 136.375 0.700 ;
        RECT 73.630 0.040 136.375 0.700 ;
        RECT 73.630 0.035 136.365 0.700 ;
        RECT 73.640 0.030 136.365 0.700 ;
        RECT 73.640 0.025 136.355 0.700 ;
        RECT 73.650 0.020 136.355 0.700 ;
        RECT 73.650 0.015 136.345 0.700 ;
        RECT 73.660 0.010 136.345 0.700 ;
        RECT 73.660 0.005 136.335 0.700 ;
        RECT 73.665 0.000 136.335 0.700 ;
      LAYER M5 ;
        RECT 73.000 0.665 137.000 0.700 ;
        RECT 73.010 0.660 136.995 0.700 ;
        RECT 73.010 0.655 136.985 0.700 ;
        RECT 73.020 0.650 136.985 0.700 ;
        RECT 73.020 0.645 136.975 0.700 ;
        RECT 73.030 0.640 136.975 0.700 ;
        RECT 73.030 0.635 136.965 0.700 ;
        RECT 73.040 0.630 136.965 0.700 ;
        RECT 73.040 0.625 136.955 0.700 ;
        RECT 73.050 0.620 136.955 0.700 ;
        RECT 73.050 0.615 136.945 0.700 ;
        RECT 73.060 0.610 136.945 0.700 ;
        RECT 73.060 0.605 136.935 0.700 ;
        RECT 73.070 0.600 136.935 0.700 ;
        RECT 73.070 0.595 136.925 0.700 ;
        RECT 73.080 0.590 136.925 0.700 ;
        RECT 73.080 0.585 136.915 0.700 ;
        RECT 73.090 0.580 136.915 0.700 ;
        RECT 73.090 0.575 136.905 0.700 ;
        RECT 73.100 0.570 136.905 0.700 ;
        RECT 73.100 0.565 136.895 0.700 ;
        RECT 73.110 0.560 136.895 0.700 ;
        RECT 73.110 0.555 136.885 0.700 ;
        RECT 73.120 0.550 136.885 0.700 ;
        RECT 73.120 0.545 136.875 0.700 ;
        RECT 73.130 0.540 136.875 0.700 ;
        RECT 73.130 0.535 136.865 0.700 ;
        RECT 73.140 0.530 136.865 0.700 ;
        RECT 73.140 0.525 136.855 0.700 ;
        RECT 73.150 0.520 136.855 0.700 ;
        RECT 73.150 0.515 136.845 0.700 ;
        RECT 73.160 0.510 136.845 0.700 ;
        RECT 73.160 0.505 136.835 0.700 ;
        RECT 73.170 0.500 136.835 0.700 ;
        RECT 73.170 0.495 136.825 0.700 ;
        RECT 73.180 0.490 136.825 0.700 ;
        RECT 73.180 0.485 136.815 0.700 ;
        RECT 73.190 0.480 136.815 0.700 ;
        RECT 73.190 0.475 136.805 0.700 ;
        RECT 73.200 0.470 136.805 0.700 ;
        RECT 73.200 0.465 136.795 0.700 ;
        RECT 73.210 0.460 136.795 0.700 ;
        RECT 73.210 0.455 136.785 0.700 ;
        RECT 73.220 0.450 136.785 0.700 ;
        RECT 73.220 0.445 136.775 0.700 ;
        RECT 73.230 0.440 136.775 0.700 ;
        RECT 73.230 0.435 136.765 0.700 ;
        RECT 73.240 0.430 136.765 0.700 ;
        RECT 73.240 0.425 136.755 0.700 ;
        RECT 73.250 0.420 136.755 0.700 ;
        RECT 73.250 0.415 136.745 0.700 ;
        RECT 73.260 0.410 136.745 0.700 ;
        RECT 73.260 0.405 136.735 0.700 ;
        RECT 73.270 0.400 136.735 0.700 ;
        RECT 73.270 0.395 136.725 0.700 ;
        RECT 73.280 0.390 136.725 0.700 ;
        RECT 73.280 0.385 136.715 0.700 ;
        RECT 73.290 0.380 136.715 0.700 ;
        RECT 73.290 0.375 136.705 0.700 ;
        RECT 73.300 0.370 136.705 0.700 ;
        RECT 73.300 0.365 136.695 0.700 ;
        RECT 73.310 0.360 136.695 0.700 ;
        RECT 73.310 0.355 136.685 0.700 ;
        RECT 73.320 0.350 136.685 0.700 ;
        RECT 73.320 0.345 136.675 0.700 ;
        RECT 73.330 0.340 136.675 0.700 ;
        RECT 73.330 0.335 136.665 0.700 ;
        RECT 73.340 0.330 136.665 0.700 ;
        RECT 73.340 0.325 136.655 0.700 ;
        RECT 73.350 0.320 136.655 0.700 ;
        RECT 73.350 0.315 136.645 0.700 ;
        RECT 73.360 0.310 136.645 0.700 ;
        RECT 73.360 0.305 136.635 0.700 ;
        RECT 73.370 0.300 136.635 0.700 ;
        RECT 73.370 0.295 136.625 0.700 ;
        RECT 73.380 0.290 136.625 0.700 ;
        RECT 73.380 0.285 136.615 0.700 ;
        RECT 73.390 0.280 136.615 0.700 ;
        RECT 73.390 0.275 136.605 0.700 ;
        RECT 73.400 0.270 136.605 0.700 ;
        RECT 73.400 0.265 136.595 0.700 ;
        RECT 73.410 0.260 136.595 0.700 ;
        RECT 73.410 0.255 136.585 0.700 ;
        RECT 73.420 0.250 136.585 0.700 ;
        RECT 73.420 0.245 136.575 0.700 ;
        RECT 73.430 0.240 136.575 0.700 ;
        RECT 73.430 0.235 136.565 0.700 ;
        RECT 73.440 0.230 136.565 0.700 ;
        RECT 73.440 0.225 136.555 0.700 ;
        RECT 73.450 0.220 136.555 0.700 ;
        RECT 73.450 0.215 136.545 0.700 ;
        RECT 73.460 0.210 136.545 0.700 ;
        RECT 73.460 0.205 136.535 0.700 ;
        RECT 73.470 0.200 136.535 0.700 ;
        RECT 73.470 0.195 136.525 0.700 ;
        RECT 73.480 0.190 136.525 0.700 ;
        RECT 73.480 0.185 136.515 0.700 ;
        RECT 73.490 0.180 136.515 0.700 ;
        RECT 73.490 0.175 136.505 0.700 ;
        RECT 73.500 0.170 136.505 0.700 ;
        RECT 73.500 0.165 136.495 0.700 ;
        RECT 73.510 0.160 136.495 0.700 ;
        RECT 73.510 0.155 136.485 0.700 ;
        RECT 73.520 0.150 136.485 0.700 ;
        RECT 73.520 0.145 136.475 0.700 ;
        RECT 73.530 0.140 136.475 0.700 ;
        RECT 73.530 0.135 136.465 0.700 ;
        RECT 73.540 0.130 136.465 0.700 ;
        RECT 73.540 0.125 136.455 0.700 ;
        RECT 73.550 0.120 136.455 0.700 ;
        RECT 73.550 0.115 136.445 0.700 ;
        RECT 73.560 0.110 136.445 0.700 ;
        RECT 73.560 0.105 136.435 0.700 ;
        RECT 73.570 0.100 136.435 0.700 ;
        RECT 73.570 0.095 136.425 0.700 ;
        RECT 73.580 0.090 136.425 0.700 ;
        RECT 73.580 0.085 136.415 0.700 ;
        RECT 73.590 0.080 136.415 0.700 ;
        RECT 73.590 0.075 136.405 0.700 ;
        RECT 73.600 0.070 136.405 0.700 ;
        RECT 73.600 0.065 136.395 0.700 ;
        RECT 73.610 0.060 136.395 0.700 ;
        RECT 73.610 0.055 136.385 0.700 ;
        RECT 73.620 0.050 136.385 0.700 ;
        RECT 73.620 0.045 136.375 0.700 ;
        RECT 73.630 0.040 136.375 0.700 ;
        RECT 73.630 0.035 136.365 0.700 ;
        RECT 73.640 0.030 136.365 0.700 ;
        RECT 73.640 0.025 136.355 0.700 ;
        RECT 73.650 0.020 136.355 0.700 ;
        RECT 73.650 0.015 136.345 0.700 ;
        RECT 73.660 0.010 136.345 0.700 ;
        RECT 73.660 0.005 136.335 0.700 ;
        RECT 73.665 0.000 136.335 0.700 ;
    END
  END XTALOUT
  PIN EO
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 92.020 173.380 93.020 174.000 ;
      LAYER V6 ;
        RECT 92.340 173.510 92.700 173.870 ;
      LAYER M4 ;
        RECT 92.020 173.380 93.020 174.000 ;
      LAYER V3 ;
        RECT 92.220 173.800 92.410 173.990 ;
        RECT 92.220 173.390 92.410 173.580 ;
        RECT 92.630 173.800 92.820 173.990 ;
        RECT 92.630 173.390 92.820 173.580 ;
      LAYER M3 ;
        RECT 92.020 173.380 93.020 174.000 ;
      LAYER V2 ;
        RECT 92.220 173.800 92.410 173.990 ;
        RECT 92.220 173.390 92.410 173.580 ;
        RECT 92.630 173.800 92.820 173.990 ;
        RECT 92.630 173.390 92.820 173.580 ;
      LAYER M2 ;
        RECT 92.420 173.300 92.620 174.000 ;
        RECT 92.020 173.380 93.020 174.000 ;
      LAYER V1 ;
        RECT 92.220 173.800 92.410 173.990 ;
        RECT 92.220 173.390 92.410 173.580 ;
        RECT 92.630 173.800 92.820 173.990 ;
        RECT 92.630 173.390 92.820 173.580 ;
      LAYER M1 ;
        RECT 92.020 173.380 93.020 174.000 ;
      LAYER M6 ;
        RECT 92.020 173.380 93.020 174.000 ;
      LAYER V5 ;
        RECT 92.220 173.800 92.410 173.990 ;
        RECT 92.220 173.390 92.410 173.580 ;
        RECT 92.630 173.800 92.820 173.990 ;
        RECT 92.630 173.390 92.820 173.580 ;
      LAYER M5 ;
        RECT 92.020 173.380 93.020 174.000 ;
      LAYER V4 ;
        RECT 92.220 173.800 92.410 173.990 ;
        RECT 92.220 173.390 92.410 173.580 ;
        RECT 92.630 173.800 92.820 173.990 ;
        RECT 92.630 173.390 92.820 173.580 ;
    END
  END EO
  PIN CK
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 80.165 173.380 81.165 174.000 ;
      LAYER V6 ;
        RECT 80.485 173.510 80.845 173.870 ;
      LAYER M4 ;
        RECT 80.165 173.380 81.165 174.000 ;
      LAYER V3 ;
        RECT 80.365 173.800 80.555 173.990 ;
        RECT 80.365 173.390 80.555 173.580 ;
        RECT 80.775 173.800 80.965 173.990 ;
        RECT 80.775 173.390 80.965 173.580 ;
      LAYER M3 ;
        RECT 80.165 173.380 81.165 174.000 ;
      LAYER V2 ;
        RECT 80.365 173.800 80.555 173.990 ;
        RECT 80.365 173.390 80.555 173.580 ;
        RECT 80.775 173.800 80.965 173.990 ;
        RECT 80.775 173.390 80.965 173.580 ;
      LAYER M2 ;
        RECT 80.165 173.300 81.165 174.000 ;
      LAYER V1 ;
        RECT 80.365 173.800 80.555 173.990 ;
        RECT 80.365 173.390 80.555 173.580 ;
        RECT 80.775 173.800 80.965 173.990 ;
        RECT 80.775 173.390 80.965 173.580 ;
      LAYER M1 ;
        RECT 80.165 173.380 81.165 174.000 ;
      LAYER M6 ;
        RECT 80.165 173.380 81.165 174.000 ;
      LAYER V5 ;
        RECT 80.365 173.800 80.555 173.990 ;
        RECT 80.365 173.390 80.555 173.580 ;
        RECT 80.775 173.800 80.965 173.990 ;
        RECT 80.775 173.390 80.965 173.580 ;
      LAYER M5 ;
        RECT 80.165 173.380 81.165 174.000 ;
      LAYER V4 ;
        RECT 80.365 173.800 80.555 173.990 ;
        RECT 80.365 173.390 80.555 173.580 ;
        RECT 80.775 173.800 80.965 173.990 ;
        RECT 80.775 173.390 80.965 173.580 ;
    END
  END CK
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.540 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.345 0.700 100.135 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 138.900 172.900 ;
        RECT 139.300 162.720 139.840 170.465 ;
        RECT 139.300 110.315 139.840 113.895 ;
        RECT 139.300 105.215 139.840 108.815 ;
        RECT 139.300 92.280 139.840 100.280 ;
        RECT 139.300 81.280 139.840 89.280 ;
        RECT 139.300 70.000 139.840 78.280 ;
        RECT 139.300 171.175 139.845 172.780 ;
        RECT 139.300 155.725 139.845 161.220 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 138.900 172.900 ;
        RECT 139.300 171.175 140.000 172.780 ;
        RECT 139.300 162.720 140.000 170.715 ;
        RECT 139.300 155.725 140.000 161.220 ;
        RECT 139.300 115.135 140.000 154.220 ;
        RECT 139.300 110.315 140.000 113.895 ;
        RECT 139.300 70.000 140.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.540 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.345 0.700 100.135 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 138.900 172.900 ;
        RECT 139.300 162.720 139.840 170.465 ;
        RECT 139.300 110.315 139.840 113.895 ;
        RECT 139.300 105.215 139.840 108.815 ;
        RECT 139.300 92.280 139.840 100.280 ;
        RECT 139.300 81.280 139.840 89.280 ;
        RECT 139.300 70.000 139.840 78.280 ;
        RECT 139.300 171.175 139.845 172.780 ;
        RECT 139.300 155.725 139.845 161.220 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 138.900 172.900 ;
        RECT 139.300 171.175 140.000 172.780 ;
        RECT 139.300 162.720 140.000 170.715 ;
        RECT 139.300 155.725 140.000 161.220 ;
        RECT 139.300 150.480 140.000 154.220 ;
        RECT 139.300 137.395 140.000 147.565 ;
        RECT 139.300 127.100 140.000 134.395 ;
        RECT 139.300 121.860 140.000 124.100 ;
        RECT 139.300 115.135 140.000 119.705 ;
        RECT 139.300 110.315 140.000 113.895 ;
        RECT 139.300 97.700 140.000 108.815 ;
        RECT 139.300 86.640 140.000 94.700 ;
        RECT 139.300 75.630 140.000 83.640 ;
        RECT 139.300 70.000 140.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 138.900 172.900 ;
        RECT 139.300 171.175 140.000 172.780 ;
        RECT 139.300 162.720 140.000 170.715 ;
        RECT 139.300 155.725 140.000 161.220 ;
        RECT 139.300 150.480 140.000 154.220 ;
        RECT 139.300 143.340 140.000 147.565 ;
        RECT 139.300 131.850 140.000 140.340 ;
        RECT 139.300 121.860 140.000 128.850 ;
        RECT 139.300 115.135 140.000 119.705 ;
        RECT 139.300 110.315 140.000 113.895 ;
        RECT 139.300 103.280 140.000 108.815 ;
        RECT 139.300 92.280 140.000 100.280 ;
        RECT 139.300 81.280 140.000 89.280 ;
        RECT 139.300 70.000 140.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 138.900 172.900 ;
        RECT 139.300 171.175 140.000 172.780 ;
        RECT 139.300 162.720 140.000 170.715 ;
        RECT 139.300 155.725 140.000 161.220 ;
        RECT 139.300 150.480 140.000 154.220 ;
        RECT 139.300 143.340 140.000 147.565 ;
        RECT 139.300 131.850 140.000 140.340 ;
        RECT 139.300 121.860 140.000 128.850 ;
        RECT 139.300 115.135 140.000 119.705 ;
        RECT 139.300 110.315 140.000 113.895 ;
        RECT 139.300 103.280 140.000 108.815 ;
        RECT 139.300 92.280 140.000 100.280 ;
        RECT 139.300 81.280 140.000 89.280 ;
        RECT 139.300 70.000 140.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.540 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.135 115.870 0.700 154.930 ;
        RECT 0.145 115.860 0.700 154.940 ;
        RECT 0.155 115.850 0.700 154.950 ;
        RECT 0.165 115.840 0.700 154.960 ;
        RECT 0.175 115.830 0.700 154.970 ;
        RECT 0.185 115.820 0.700 154.980 ;
        RECT 0.195 115.810 0.700 154.990 ;
        RECT 0.205 115.800 0.700 155.000 ;
        RECT 0.215 115.790 0.700 155.010 ;
        RECT 0.225 115.780 0.700 155.020 ;
        RECT 0.235 115.770 0.700 155.030 ;
        RECT 0.245 115.760 0.700 155.040 ;
        RECT 0.255 115.750 0.700 155.050 ;
        RECT 0.270 115.735 0.700 155.055 ;
        RECT 0.260 115.745 0.700 155.055 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.345 0.700 100.135 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 138.900 172.900 ;
        RECT 139.300 162.720 139.840 170.465 ;
        RECT 139.300 110.315 139.840 113.895 ;
        RECT 139.300 105.215 139.840 108.815 ;
        RECT 139.300 92.280 139.840 100.280 ;
        RECT 139.300 81.280 139.840 89.280 ;
        RECT 139.300 70.000 139.840 78.280 ;
        RECT 139.300 171.175 139.845 172.780 ;
        RECT 139.300 155.725 139.845 161.220 ;
        RECT 139.300 115.735 139.730 155.055 ;
        RECT 139.300 115.870 139.865 154.930 ;
        RECT 139.300 115.865 139.860 154.935 ;
        RECT 139.300 115.855 139.850 154.945 ;
        RECT 139.300 115.845 139.840 154.955 ;
        RECT 139.300 115.835 139.830 154.965 ;
        RECT 139.300 115.825 139.820 154.975 ;
        RECT 139.300 115.815 139.810 154.985 ;
        RECT 139.300 115.805 139.800 154.995 ;
        RECT 139.300 115.795 139.790 155.005 ;
        RECT 139.300 115.785 139.780 155.015 ;
        RECT 139.300 115.775 139.770 155.025 ;
        RECT 139.300 115.765 139.760 155.035 ;
        RECT 139.300 115.755 139.750 155.045 ;
        RECT 139.300 115.745 139.740 155.055 ;
  END 
END PLOSC14M

MACRO PLFILLER70
  CLASS  PAD ;
  FOREIGN PLFILLER70 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.395 150.750 0.700 154.220 ;
        RECT 0.395 143.565 0.700 147.565 ;
        RECT 0.395 131.850 0.700 140.340 ;
        RECT 0.395 121.860 0.700 128.665 ;
        RECT 0.395 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.395 103.850 0.700 108.420 ;
        RECT 0.395 92.280 0.700 100.280 ;
        RECT 0.395 81.280 0.700 89.280 ;
        RECT 0.395 70.280 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 150.750 69.605 154.220 ;
        RECT 69.300 143.565 69.605 147.565 ;
        RECT 69.300 131.850 69.605 140.340 ;
        RECT 69.300 121.860 69.605 128.665 ;
        RECT 69.300 115.135 69.605 119.705 ;
        RECT 69.300 81.280 69.685 89.280 ;
        RECT 69.300 103.850 69.750 108.420 ;
        RECT 69.300 92.280 69.770 100.280 ;
        RECT 69.300 70.280 69.810 78.280 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.395 150.720 0.700 154.220 ;
        RECT 0.395 143.565 0.700 147.565 ;
        RECT 0.395 131.850 0.700 140.340 ;
        RECT 0.395 121.860 0.700 128.665 ;
        RECT 0.395 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.395 103.850 0.700 108.420 ;
        RECT 0.395 92.280 0.700 100.280 ;
        RECT 0.395 81.280 0.700 89.280 ;
        RECT 0.395 70.280 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 150.720 69.605 154.220 ;
        RECT 69.300 143.565 69.605 147.565 ;
        RECT 69.300 131.850 69.605 140.340 ;
        RECT 69.300 121.860 69.605 128.665 ;
        RECT 69.300 115.135 69.605 119.705 ;
        RECT 69.300 81.280 69.685 89.280 ;
        RECT 69.300 103.850 69.750 108.420 ;
        RECT 69.300 92.280 69.770 100.280 ;
        RECT 69.300 70.280 69.810 78.280 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.395 150.720 0.700 154.220 ;
        RECT 0.395 143.565 0.700 147.565 ;
        RECT 0.395 131.850 0.700 140.340 ;
        RECT 0.395 121.860 0.700 128.665 ;
        RECT 0.395 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.395 103.850 0.700 108.420 ;
        RECT 0.395 92.280 0.700 100.280 ;
        RECT 0.395 81.280 0.700 89.280 ;
        RECT 0.395 70.280 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 150.720 69.605 154.220 ;
        RECT 69.300 143.565 69.605 147.565 ;
        RECT 69.300 131.850 69.605 140.340 ;
        RECT 69.300 121.860 69.605 128.665 ;
        RECT 69.300 115.135 69.605 119.705 ;
        RECT 69.300 81.280 69.685 89.280 ;
        RECT 69.300 103.850 69.750 108.420 ;
        RECT 69.300 92.280 69.770 100.280 ;
        RECT 69.300 70.280 69.810 78.280 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
  END 
END PLFILLER70

MACRO PLFILLER35
  CLASS  PAD ;
  FOREIGN PLFILLER35 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.395 150.750 0.700 154.220 ;
        RECT 0.395 143.565 0.700 147.565 ;
        RECT 0.395 131.850 0.700 140.340 ;
        RECT 0.395 121.860 0.700 128.665 ;
        RECT 0.395 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.395 103.850 0.700 108.420 ;
        RECT 0.395 92.280 0.700 100.280 ;
        RECT 0.395 81.280 0.700 89.280 ;
        RECT 0.395 70.280 0.700 78.280 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 150.750 34.605 154.220 ;
        RECT 34.300 143.565 34.605 147.565 ;
        RECT 34.300 131.850 34.605 140.340 ;
        RECT 34.300 121.860 34.605 128.665 ;
        RECT 34.300 115.135 34.605 119.705 ;
        RECT 34.300 81.280 34.685 89.280 ;
        RECT 34.300 103.850 34.750 108.420 ;
        RECT 34.300 92.280 34.770 100.280 ;
        RECT 34.300 70.280 34.810 78.280 ;
        RECT 34.300 171.175 34.840 172.780 ;
        RECT 34.300 162.720 34.840 170.465 ;
        RECT 34.300 155.725 34.840 161.220 ;
        RECT 34.300 110.315 34.840 113.895 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 171.175 35.000 172.780 ;
        RECT 34.300 162.720 35.000 170.715 ;
        RECT 34.300 155.725 35.000 161.220 ;
        RECT 34.300 115.135 35.000 154.220 ;
        RECT 34.300 110.315 35.000 113.895 ;
        RECT 34.300 70.000 35.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.395 150.720 0.700 154.220 ;
        RECT 0.395 143.565 0.700 147.565 ;
        RECT 0.395 131.850 0.700 140.340 ;
        RECT 0.395 121.860 0.700 128.665 ;
        RECT 0.395 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.395 103.850 0.700 108.420 ;
        RECT 0.395 92.280 0.700 100.280 ;
        RECT 0.395 81.280 0.700 89.280 ;
        RECT 0.395 70.280 0.700 78.280 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 150.720 34.605 154.220 ;
        RECT 34.300 143.565 34.605 147.565 ;
        RECT 34.300 131.850 34.605 140.340 ;
        RECT 34.300 121.860 34.605 128.665 ;
        RECT 34.300 115.135 34.605 119.705 ;
        RECT 34.300 81.280 34.685 89.280 ;
        RECT 34.300 103.850 34.750 108.420 ;
        RECT 34.300 92.280 34.770 100.280 ;
        RECT 34.300 70.280 34.810 78.280 ;
        RECT 34.300 171.175 34.840 172.780 ;
        RECT 34.300 162.720 34.840 170.465 ;
        RECT 34.300 155.725 34.840 161.220 ;
        RECT 34.300 110.315 34.840 113.895 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 171.175 35.000 172.780 ;
        RECT 34.300 162.720 35.000 170.715 ;
        RECT 34.300 155.725 35.000 161.220 ;
        RECT 34.300 150.480 35.000 154.220 ;
        RECT 34.300 137.395 35.000 147.565 ;
        RECT 34.300 127.100 35.000 134.395 ;
        RECT 34.300 121.860 35.000 124.100 ;
        RECT 34.300 115.135 35.000 119.705 ;
        RECT 34.300 110.315 35.000 113.895 ;
        RECT 34.300 97.700 35.000 108.815 ;
        RECT 34.300 86.640 35.000 94.700 ;
        RECT 34.300 75.630 35.000 83.640 ;
        RECT 34.300 70.000 35.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 171.175 35.000 172.780 ;
        RECT 34.300 162.720 35.000 170.715 ;
        RECT 34.300 155.725 35.000 161.220 ;
        RECT 34.300 150.480 35.000 154.220 ;
        RECT 34.300 143.340 35.000 147.565 ;
        RECT 34.300 131.850 35.000 140.340 ;
        RECT 34.300 121.860 35.000 128.850 ;
        RECT 34.300 115.135 35.000 119.705 ;
        RECT 34.300 110.315 35.000 113.895 ;
        RECT 34.300 103.280 35.000 108.815 ;
        RECT 34.300 92.280 35.000 100.280 ;
        RECT 34.300 81.280 35.000 89.280 ;
        RECT 34.300 70.000 35.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 171.175 35.000 172.780 ;
        RECT 34.300 162.720 35.000 170.715 ;
        RECT 34.300 155.725 35.000 161.220 ;
        RECT 34.300 150.480 35.000 154.220 ;
        RECT 34.300 143.340 35.000 147.565 ;
        RECT 34.300 131.850 35.000 140.340 ;
        RECT 34.300 121.860 35.000 128.850 ;
        RECT 34.300 115.135 35.000 119.705 ;
        RECT 34.300 110.315 35.000 113.895 ;
        RECT 34.300 103.280 35.000 108.815 ;
        RECT 34.300 92.280 35.000 100.280 ;
        RECT 34.300 81.280 35.000 89.280 ;
        RECT 34.300 70.000 35.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.395 150.720 0.700 154.220 ;
        RECT 0.395 143.565 0.700 147.565 ;
        RECT 0.395 131.850 0.700 140.340 ;
        RECT 0.395 121.860 0.700 128.665 ;
        RECT 0.395 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.395 103.850 0.700 108.420 ;
        RECT 0.395 92.280 0.700 100.280 ;
        RECT 0.395 81.280 0.700 89.280 ;
        RECT 0.395 70.280 0.700 78.280 ;
        RECT 1.100 1.100 33.900 172.900 ;
        RECT 34.300 150.720 34.605 154.220 ;
        RECT 34.300 143.565 34.605 147.565 ;
        RECT 34.300 131.850 34.605 140.340 ;
        RECT 34.300 121.860 34.605 128.665 ;
        RECT 34.300 115.135 34.605 119.705 ;
        RECT 34.300 81.280 34.685 89.280 ;
        RECT 34.300 103.850 34.750 108.420 ;
        RECT 34.300 92.280 34.770 100.280 ;
        RECT 34.300 70.280 34.810 78.280 ;
        RECT 34.300 171.175 34.840 172.780 ;
        RECT 34.300 162.720 34.840 170.465 ;
        RECT 34.300 155.725 34.840 161.220 ;
        RECT 34.300 110.315 34.840 113.895 ;
  END 
END PLFILLER35

MACRO PLFILLER20
  CLASS  PAD ;
  FOREIGN PLFILLER20 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.395 150.750 0.700 154.220 ;
        RECT 0.395 143.565 0.700 147.565 ;
        RECT 0.395 131.850 0.700 140.340 ;
        RECT 0.395 121.860 0.700 128.665 ;
        RECT 0.395 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.395 103.850 0.700 108.420 ;
        RECT 0.395 92.280 0.700 100.280 ;
        RECT 0.395 81.280 0.700 89.280 ;
        RECT 0.395 70.280 0.700 78.280 ;
        RECT 1.100 1.100 18.900 172.900 ;
        RECT 19.300 150.750 19.605 154.220 ;
        RECT 19.300 143.565 19.605 147.565 ;
        RECT 19.300 131.850 19.605 140.340 ;
        RECT 19.300 121.860 19.605 128.665 ;
        RECT 19.300 115.135 19.605 119.705 ;
        RECT 19.300 81.280 19.685 89.280 ;
        RECT 19.300 103.850 19.750 108.420 ;
        RECT 19.300 92.280 19.770 100.280 ;
        RECT 19.300 70.280 19.810 78.280 ;
        RECT 19.300 171.175 19.840 172.780 ;
        RECT 19.300 162.720 19.840 170.465 ;
        RECT 19.300 155.725 19.840 161.220 ;
        RECT 19.300 110.315 19.840 113.895 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 18.900 172.900 ;
        RECT 19.300 171.175 20.000 172.780 ;
        RECT 19.300 162.720 20.000 170.715 ;
        RECT 19.300 155.725 20.000 161.220 ;
        RECT 19.300 115.135 20.000 154.220 ;
        RECT 19.300 110.315 20.000 113.895 ;
        RECT 19.300 70.000 20.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.395 150.720 0.700 154.220 ;
        RECT 0.395 143.565 0.700 147.565 ;
        RECT 0.395 131.850 0.700 140.340 ;
        RECT 0.395 121.860 0.700 128.665 ;
        RECT 0.395 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.395 103.850 0.700 108.420 ;
        RECT 0.395 92.280 0.700 100.280 ;
        RECT 0.395 81.280 0.700 89.280 ;
        RECT 0.395 70.280 0.700 78.280 ;
        RECT 1.100 1.100 18.900 172.900 ;
        RECT 19.300 150.720 19.605 154.220 ;
        RECT 19.300 143.565 19.605 147.565 ;
        RECT 19.300 131.850 19.605 140.340 ;
        RECT 19.300 121.860 19.605 128.665 ;
        RECT 19.300 115.135 19.605 119.705 ;
        RECT 19.300 81.280 19.685 89.280 ;
        RECT 19.300 103.850 19.750 108.420 ;
        RECT 19.300 92.280 19.770 100.280 ;
        RECT 19.300 70.280 19.810 78.280 ;
        RECT 19.300 171.175 19.840 172.780 ;
        RECT 19.300 162.720 19.840 170.465 ;
        RECT 19.300 155.725 19.840 161.220 ;
        RECT 19.300 110.315 19.840 113.895 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 18.900 172.900 ;
        RECT 19.300 171.175 20.000 172.780 ;
        RECT 19.300 162.720 20.000 170.715 ;
        RECT 19.300 155.725 20.000 161.220 ;
        RECT 19.300 150.480 20.000 154.220 ;
        RECT 19.300 137.395 20.000 147.565 ;
        RECT 19.300 127.100 20.000 134.395 ;
        RECT 19.300 121.860 20.000 124.100 ;
        RECT 19.300 115.135 20.000 119.705 ;
        RECT 19.300 110.315 20.000 113.895 ;
        RECT 19.300 97.700 20.000 108.815 ;
        RECT 19.300 86.640 20.000 94.700 ;
        RECT 19.300 75.630 20.000 83.640 ;
        RECT 19.300 70.000 20.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 18.900 172.900 ;
        RECT 19.300 171.175 20.000 172.780 ;
        RECT 19.300 162.720 20.000 170.715 ;
        RECT 19.300 155.725 20.000 161.220 ;
        RECT 19.300 150.480 20.000 154.220 ;
        RECT 19.300 143.340 20.000 147.565 ;
        RECT 19.300 131.850 20.000 140.340 ;
        RECT 19.300 121.860 20.000 128.850 ;
        RECT 19.300 115.135 20.000 119.705 ;
        RECT 19.300 110.315 20.000 113.895 ;
        RECT 19.300 103.280 20.000 108.815 ;
        RECT 19.300 92.280 20.000 100.280 ;
        RECT 19.300 81.280 20.000 89.280 ;
        RECT 19.300 70.000 20.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 18.900 172.900 ;
        RECT 19.300 171.175 20.000 172.780 ;
        RECT 19.300 162.720 20.000 170.715 ;
        RECT 19.300 155.725 20.000 161.220 ;
        RECT 19.300 150.480 20.000 154.220 ;
        RECT 19.300 143.340 20.000 147.565 ;
        RECT 19.300 131.850 20.000 140.340 ;
        RECT 19.300 121.860 20.000 128.850 ;
        RECT 19.300 115.135 20.000 119.705 ;
        RECT 19.300 110.315 20.000 113.895 ;
        RECT 19.300 103.280 20.000 108.815 ;
        RECT 19.300 92.280 20.000 100.280 ;
        RECT 19.300 81.280 20.000 89.280 ;
        RECT 19.300 70.000 20.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.395 150.720 0.700 154.220 ;
        RECT 0.395 143.565 0.700 147.565 ;
        RECT 0.395 131.850 0.700 140.340 ;
        RECT 0.395 121.860 0.700 128.665 ;
        RECT 0.395 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.395 103.850 0.700 108.420 ;
        RECT 0.395 92.280 0.700 100.280 ;
        RECT 0.395 81.280 0.700 89.280 ;
        RECT 0.395 70.280 0.700 78.280 ;
        RECT 1.100 1.100 18.900 172.900 ;
        RECT 19.300 150.720 19.605 154.220 ;
        RECT 19.300 143.565 19.605 147.565 ;
        RECT 19.300 131.850 19.605 140.340 ;
        RECT 19.300 121.860 19.605 128.665 ;
        RECT 19.300 115.135 19.605 119.705 ;
        RECT 19.300 81.280 19.685 89.280 ;
        RECT 19.300 103.850 19.750 108.420 ;
        RECT 19.300 92.280 19.770 100.280 ;
        RECT 19.300 70.280 19.810 78.280 ;
        RECT 19.300 171.175 19.840 172.780 ;
        RECT 19.300 162.720 19.840 170.465 ;
        RECT 19.300 155.725 19.840 161.220 ;
        RECT 19.300 110.315 19.840 113.895 ;
  END 
END PLFILLER20

MACRO PLFILLER10
  CLASS  PAD ;
  FOREIGN PLFILLER10 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.395 150.750 0.700 154.220 ;
        RECT 0.395 143.565 0.700 147.565 ;
        RECT 0.395 131.850 0.700 140.340 ;
        RECT 0.395 121.860 0.700 128.665 ;
        RECT 0.395 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.395 103.850 0.700 108.420 ;
        RECT 0.395 92.280 0.700 100.280 ;
        RECT 0.395 81.280 0.700 89.280 ;
        RECT 0.395 70.280 0.700 78.280 ;
        RECT 1.100 1.100 8.900 172.900 ;
        RECT 9.300 150.750 9.605 154.220 ;
        RECT 9.300 143.565 9.605 147.565 ;
        RECT 9.300 131.850 9.605 140.340 ;
        RECT 9.300 121.860 9.605 128.665 ;
        RECT 9.300 115.135 9.605 119.705 ;
        RECT 9.300 81.280 9.685 89.280 ;
        RECT 9.300 103.850 9.750 108.420 ;
        RECT 9.300 92.280 9.770 100.280 ;
        RECT 9.300 70.280 9.810 78.280 ;
        RECT 9.300 171.175 9.840 172.780 ;
        RECT 9.300 162.720 9.840 170.465 ;
        RECT 9.300 155.725 9.840 161.220 ;
        RECT 9.300 110.315 9.840 113.895 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 8.900 172.900 ;
        RECT 9.300 171.175 10.000 172.780 ;
        RECT 9.300 162.720 10.000 170.715 ;
        RECT 9.300 155.725 10.000 161.220 ;
        RECT 9.300 115.135 10.000 154.220 ;
        RECT 9.300 110.315 10.000 113.895 ;
        RECT 9.300 70.000 10.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.395 150.720 0.700 154.220 ;
        RECT 0.395 143.565 0.700 147.565 ;
        RECT 0.395 131.850 0.700 140.340 ;
        RECT 0.395 121.860 0.700 128.665 ;
        RECT 0.395 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.395 103.850 0.700 108.420 ;
        RECT 0.395 92.280 0.700 100.280 ;
        RECT 0.395 81.280 0.700 89.280 ;
        RECT 0.395 70.280 0.700 78.280 ;
        RECT 1.100 1.100 8.900 172.900 ;
        RECT 9.300 150.720 9.605 154.220 ;
        RECT 9.300 143.565 9.605 147.565 ;
        RECT 9.300 131.850 9.605 140.340 ;
        RECT 9.300 121.860 9.605 128.665 ;
        RECT 9.300 115.135 9.605 119.705 ;
        RECT 9.300 81.280 9.685 89.280 ;
        RECT 9.300 103.850 9.750 108.420 ;
        RECT 9.300 92.280 9.770 100.280 ;
        RECT 9.300 70.280 9.810 78.280 ;
        RECT 9.300 171.175 9.840 172.780 ;
        RECT 9.300 162.720 9.840 170.465 ;
        RECT 9.300 155.725 9.840 161.220 ;
        RECT 9.300 110.315 9.840 113.895 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 8.900 172.900 ;
        RECT 9.300 171.175 10.000 172.780 ;
        RECT 9.300 162.720 10.000 170.715 ;
        RECT 9.300 155.725 10.000 161.220 ;
        RECT 9.300 150.480 10.000 154.220 ;
        RECT 9.300 137.395 10.000 147.565 ;
        RECT 9.300 127.100 10.000 134.395 ;
        RECT 9.300 121.860 10.000 124.100 ;
        RECT 9.300 115.135 10.000 119.705 ;
        RECT 9.300 110.315 10.000 113.895 ;
        RECT 9.300 97.700 10.000 108.815 ;
        RECT 9.300 86.640 10.000 94.700 ;
        RECT 9.300 75.630 10.000 83.640 ;
        RECT 9.300 70.000 10.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 8.900 172.900 ;
        RECT 9.300 171.175 10.000 172.780 ;
        RECT 9.300 162.720 10.000 170.715 ;
        RECT 9.300 155.725 10.000 161.220 ;
        RECT 9.300 150.480 10.000 154.220 ;
        RECT 9.300 143.340 10.000 147.565 ;
        RECT 9.300 131.850 10.000 140.340 ;
        RECT 9.300 121.860 10.000 128.850 ;
        RECT 9.300 115.135 10.000 119.705 ;
        RECT 9.300 110.315 10.000 113.895 ;
        RECT 9.300 103.280 10.000 108.815 ;
        RECT 9.300 92.280 10.000 100.280 ;
        RECT 9.300 81.280 10.000 89.280 ;
        RECT 9.300 70.000 10.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 8.900 172.900 ;
        RECT 9.300 171.175 10.000 172.780 ;
        RECT 9.300 162.720 10.000 170.715 ;
        RECT 9.300 155.725 10.000 161.220 ;
        RECT 9.300 150.480 10.000 154.220 ;
        RECT 9.300 143.340 10.000 147.565 ;
        RECT 9.300 131.850 10.000 140.340 ;
        RECT 9.300 121.860 10.000 128.850 ;
        RECT 9.300 115.135 10.000 119.705 ;
        RECT 9.300 110.315 10.000 113.895 ;
        RECT 9.300 103.280 10.000 108.815 ;
        RECT 9.300 92.280 10.000 100.280 ;
        RECT 9.300 81.280 10.000 89.280 ;
        RECT 9.300 70.000 10.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.395 150.720 0.700 154.220 ;
        RECT 0.395 143.565 0.700 147.565 ;
        RECT 0.395 131.850 0.700 140.340 ;
        RECT 0.395 121.860 0.700 128.665 ;
        RECT 0.395 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.395 103.850 0.700 108.420 ;
        RECT 0.395 92.280 0.700 100.280 ;
        RECT 0.395 81.280 0.700 89.280 ;
        RECT 0.395 70.280 0.700 78.280 ;
        RECT 1.100 1.100 8.900 172.900 ;
        RECT 9.300 150.720 9.605 154.220 ;
        RECT 9.300 143.565 9.605 147.565 ;
        RECT 9.300 131.850 9.605 140.340 ;
        RECT 9.300 121.860 9.605 128.665 ;
        RECT 9.300 115.135 9.605 119.705 ;
        RECT 9.300 81.280 9.685 89.280 ;
        RECT 9.300 103.850 9.750 108.420 ;
        RECT 9.300 92.280 9.770 100.280 ;
        RECT 9.300 70.280 9.810 78.280 ;
        RECT 9.300 171.175 9.840 172.780 ;
        RECT 9.300 162.720 9.840 170.465 ;
        RECT 9.300 155.725 9.840 161.220 ;
        RECT 9.300 110.315 9.840 113.895 ;
  END 
END PLFILLER10

MACRO PLFILLER5
  CLASS  PAD ;
  FOREIGN PLFILLER5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.395 150.750 0.700 154.220 ;
        RECT 0.395 143.565 0.700 147.565 ;
        RECT 0.395 131.850 0.700 140.340 ;
        RECT 0.395 121.860 0.700 128.665 ;
        RECT 0.395 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.395 103.850 0.700 108.420 ;
        RECT 0.395 92.280 0.700 100.280 ;
        RECT 0.395 81.280 0.700 89.280 ;
        RECT 0.395 70.280 0.700 78.280 ;
        RECT 1.100 1.100 3.900 172.900 ;
        RECT 4.300 150.750 4.605 154.220 ;
        RECT 4.300 143.565 4.605 147.565 ;
        RECT 4.300 131.850 4.605 140.340 ;
        RECT 4.300 121.860 4.605 128.665 ;
        RECT 4.300 115.135 4.605 119.705 ;
        RECT 4.300 81.280 4.685 89.280 ;
        RECT 4.300 103.850 4.750 108.420 ;
        RECT 4.300 92.280 4.770 100.280 ;
        RECT 4.300 70.280 4.810 78.280 ;
        RECT 4.300 171.175 4.840 172.780 ;
        RECT 4.300 162.720 4.840 170.465 ;
        RECT 4.300 155.725 4.840 161.220 ;
        RECT 4.300 110.315 4.840 113.895 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 3.900 172.900 ;
        RECT 4.300 171.175 5.000 172.780 ;
        RECT 4.300 162.720 5.000 170.715 ;
        RECT 4.300 155.725 5.000 161.220 ;
        RECT 4.300 115.135 5.000 154.220 ;
        RECT 4.300 110.315 5.000 113.895 ;
        RECT 4.300 70.000 5.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.395 150.720 0.700 154.220 ;
        RECT 0.395 143.565 0.700 147.565 ;
        RECT 0.395 131.850 0.700 140.340 ;
        RECT 0.395 121.860 0.700 128.665 ;
        RECT 0.395 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.395 103.850 0.700 108.420 ;
        RECT 0.395 92.280 0.700 100.280 ;
        RECT 0.395 81.280 0.700 89.280 ;
        RECT 0.395 70.280 0.700 78.280 ;
        RECT 1.100 1.100 3.900 172.900 ;
        RECT 4.300 150.720 4.605 154.220 ;
        RECT 4.300 143.565 4.605 147.565 ;
        RECT 4.300 131.850 4.605 140.340 ;
        RECT 4.300 121.860 4.605 128.665 ;
        RECT 4.300 115.135 4.605 119.705 ;
        RECT 4.300 81.280 4.685 89.280 ;
        RECT 4.300 103.850 4.750 108.420 ;
        RECT 4.300 92.280 4.770 100.280 ;
        RECT 4.300 70.280 4.810 78.280 ;
        RECT 4.300 171.175 4.840 172.780 ;
        RECT 4.300 162.720 4.840 170.465 ;
        RECT 4.300 155.725 4.840 161.220 ;
        RECT 4.300 110.315 4.840 113.895 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 3.900 172.900 ;
        RECT 4.300 171.175 5.000 172.780 ;
        RECT 4.300 162.720 5.000 170.715 ;
        RECT 4.300 155.725 5.000 161.220 ;
        RECT 4.300 150.480 5.000 154.220 ;
        RECT 4.300 137.395 5.000 147.565 ;
        RECT 4.300 127.100 5.000 134.395 ;
        RECT 4.300 121.860 5.000 124.100 ;
        RECT 4.300 115.135 5.000 119.705 ;
        RECT 4.300 110.315 5.000 113.895 ;
        RECT 4.300 97.700 5.000 108.815 ;
        RECT 4.300 86.640 5.000 94.700 ;
        RECT 4.300 75.630 5.000 83.640 ;
        RECT 4.300 70.000 5.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 3.900 172.900 ;
        RECT 4.300 171.175 5.000 172.780 ;
        RECT 4.300 162.720 5.000 170.715 ;
        RECT 4.300 155.725 5.000 161.220 ;
        RECT 4.300 150.480 5.000 154.220 ;
        RECT 4.300 143.340 5.000 147.565 ;
        RECT 4.300 131.850 5.000 140.340 ;
        RECT 4.300 121.860 5.000 128.850 ;
        RECT 4.300 115.135 5.000 119.705 ;
        RECT 4.300 110.315 5.000 113.895 ;
        RECT 4.300 103.280 5.000 108.815 ;
        RECT 4.300 92.280 5.000 100.280 ;
        RECT 4.300 81.280 5.000 89.280 ;
        RECT 4.300 70.000 5.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 3.900 172.900 ;
        RECT 4.300 171.175 5.000 172.780 ;
        RECT 4.300 162.720 5.000 170.715 ;
        RECT 4.300 155.725 5.000 161.220 ;
        RECT 4.300 150.480 5.000 154.220 ;
        RECT 4.300 143.340 5.000 147.565 ;
        RECT 4.300 131.850 5.000 140.340 ;
        RECT 4.300 121.860 5.000 128.850 ;
        RECT 4.300 115.135 5.000 119.705 ;
        RECT 4.300 110.315 5.000 113.895 ;
        RECT 4.300 103.280 5.000 108.815 ;
        RECT 4.300 92.280 5.000 100.280 ;
        RECT 4.300 81.280 5.000 89.280 ;
        RECT 4.300 70.000 5.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.395 150.720 0.700 154.220 ;
        RECT 0.395 143.565 0.700 147.565 ;
        RECT 0.395 131.850 0.700 140.340 ;
        RECT 0.395 121.860 0.700 128.665 ;
        RECT 0.395 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.395 103.850 0.700 108.420 ;
        RECT 0.395 92.280 0.700 100.280 ;
        RECT 0.395 81.280 0.700 89.280 ;
        RECT 0.395 70.280 0.700 78.280 ;
        RECT 1.100 1.100 3.900 172.900 ;
        RECT 4.300 150.720 4.605 154.220 ;
        RECT 4.300 143.565 4.605 147.565 ;
        RECT 4.300 131.850 4.605 140.340 ;
        RECT 4.300 121.860 4.605 128.665 ;
        RECT 4.300 115.135 4.605 119.705 ;
        RECT 4.300 81.280 4.685 89.280 ;
        RECT 4.300 103.850 4.750 108.420 ;
        RECT 4.300 92.280 4.770 100.280 ;
        RECT 4.300 70.280 4.810 78.280 ;
        RECT 4.300 171.175 4.840 172.780 ;
        RECT 4.300 162.720 4.840 170.465 ;
        RECT 4.300 155.725 4.840 161.220 ;
        RECT 4.300 110.315 4.840 113.895 ;
  END 
END PLFILLER5

MACRO PLFILLER0005
  CLASS  PAD ;
  FOREIGN PLFILLER0005 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.005 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M1 ;
        RECT 0.000 171.175 0.005 172.780 ;
        RECT 0.000 162.720 0.005 170.715 ;
        RECT 0.000 155.725 0.005 161.220 ;
        RECT 0.000 115.135 0.005 154.220 ;
        RECT 0.000 110.315 0.005 113.895 ;
        RECT 0.000 70.000 0.005 108.815 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.005 172.780 ;
        RECT 0.000 162.720 0.005 170.715 ;
        RECT 0.000 155.725 0.005 161.220 ;
        RECT 0.000 150.480 0.005 154.220 ;
        RECT 0.000 137.395 0.005 147.565 ;
        RECT 0.000 127.100 0.005 134.395 ;
        RECT 0.000 121.860 0.005 124.100 ;
        RECT 0.000 115.135 0.005 119.705 ;
        RECT 0.000 110.315 0.005 113.895 ;
        RECT 0.000 97.700 0.005 108.815 ;
        RECT 0.000 86.640 0.005 94.700 ;
        RECT 0.000 75.630 0.005 83.640 ;
        RECT 0.000 70.000 0.005 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.005 172.780 ;
        RECT 0.000 162.720 0.005 170.715 ;
        RECT 0.000 155.725 0.005 161.220 ;
        RECT 0.000 150.480 0.005 154.220 ;
        RECT 0.000 143.340 0.005 147.565 ;
        RECT 0.000 131.850 0.005 140.340 ;
        RECT 0.000 121.860 0.005 128.850 ;
        RECT 0.000 115.135 0.005 119.705 ;
        RECT 0.000 110.315 0.005 113.895 ;
        RECT 0.000 103.280 0.005 108.815 ;
        RECT 0.000 92.280 0.005 100.280 ;
        RECT 0.000 81.280 0.005 89.280 ;
        RECT 0.000 70.000 0.005 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.005 172.780 ;
        RECT 0.000 162.720 0.005 170.715 ;
        RECT 0.000 155.725 0.005 161.220 ;
        RECT 0.000 150.480 0.005 154.220 ;
        RECT 0.000 143.340 0.005 147.565 ;
        RECT 0.000 131.850 0.005 140.340 ;
        RECT 0.000 121.860 0.005 128.850 ;
        RECT 0.000 115.135 0.005 119.705 ;
        RECT 0.000 110.315 0.005 113.895 ;
        RECT 0.000 103.280 0.005 108.815 ;
        RECT 0.000 92.280 0.005 100.280 ;
        RECT 0.000 81.280 0.005 89.280 ;
        RECT 0.000 70.000 0.005 78.280 ;
  END 
END PLFILLER0005

MACRO PLFILLER1
  CLASS  PAD ;
  FOREIGN PLFILLER1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 0.155 171.175 0.845 172.780 ;
        RECT 0.155 162.720 0.845 170.465 ;
        RECT 0.155 155.725 0.845 161.220 ;
        RECT 0.155 150.745 0.845 154.220 ;
        RECT 0.155 115.135 0.845 119.690 ;
        RECT 0.155 110.315 0.845 113.895 ;
        RECT 0.155 104.990 0.845 108.815 ;
        RECT 0.155 92.280 0.845 100.280 ;
        RECT 0.155 81.280 0.845 89.280 ;
        RECT 0.155 70.280 0.845 78.280 ;
      LAYER M1 ;
        RECT 0.000 171.175 1.000 172.780 ;
        RECT 0.000 162.720 1.000 170.715 ;
        RECT 0.000 155.725 1.000 161.220 ;
        RECT 0.000 115.135 1.000 154.220 ;
        RECT 0.000 110.315 1.000 113.895 ;
        RECT 0.000 70.000 1.000 108.815 ;
      LAYER M3 ;
        RECT 0.155 171.175 0.845 172.780 ;
        RECT 0.155 162.720 0.845 170.465 ;
        RECT 0.155 155.725 0.845 161.220 ;
        RECT 0.155 150.745 0.845 154.220 ;
        RECT 0.155 115.135 0.845 119.690 ;
        RECT 0.155 110.315 0.845 113.895 ;
        RECT 0.155 104.990 0.845 108.815 ;
        RECT 0.155 92.280 0.845 100.280 ;
        RECT 0.155 81.280 0.845 89.280 ;
        RECT 0.155 70.280 0.845 78.280 ;
      LAYER M6 ;
        RECT 0.000 171.175 1.000 172.780 ;
        RECT 0.000 162.720 1.000 170.715 ;
        RECT 0.000 155.725 1.000 161.220 ;
        RECT 0.000 150.480 1.000 154.220 ;
        RECT 0.000 137.395 1.000 147.565 ;
        RECT 0.000 127.100 1.000 134.395 ;
        RECT 0.000 121.860 1.000 124.100 ;
        RECT 0.000 115.135 1.000 119.705 ;
        RECT 0.000 110.315 1.000 113.895 ;
        RECT 0.000 97.700 1.000 108.815 ;
        RECT 0.000 86.640 1.000 94.700 ;
        RECT 0.000 75.630 1.000 83.640 ;
        RECT 0.000 70.000 1.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 1.000 172.780 ;
        RECT 0.000 162.720 1.000 170.715 ;
        RECT 0.000 155.725 1.000 161.220 ;
        RECT 0.000 150.480 1.000 154.220 ;
        RECT 0.000 143.565 1.000 147.565 ;
        RECT 0.000 131.850 1.000 140.340 ;
        RECT 0.000 121.860 1.000 128.850 ;
        RECT 0.000 115.135 1.000 119.705 ;
        RECT 0.000 110.315 1.000 113.895 ;
        RECT 0.000 103.280 1.000 108.815 ;
        RECT 0.000 92.280 1.000 100.280 ;
        RECT 0.000 81.280 1.000 89.280 ;
        RECT 0.000 70.000 1.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 1.000 172.780 ;
        RECT 0.000 162.720 1.000 170.715 ;
        RECT 0.000 155.725 1.000 161.220 ;
        RECT 0.000 150.480 1.000 154.220 ;
        RECT 0.000 143.565 1.000 147.565 ;
        RECT 0.000 131.850 1.000 140.340 ;
        RECT 0.000 121.860 1.000 128.850 ;
        RECT 0.000 115.135 1.000 119.705 ;
        RECT 0.000 110.315 1.000 113.895 ;
        RECT 0.000 103.280 1.000 108.815 ;
        RECT 0.000 92.280 1.000 100.280 ;
        RECT 0.000 81.280 1.000 89.280 ;
        RECT 0.000 70.520 1.000 78.280 ;
      LAYER M2 ;
        RECT 0.155 171.175 0.845 172.780 ;
        RECT 0.155 162.720 0.845 170.465 ;
        RECT 0.155 155.725 0.845 161.220 ;
        RECT 0.155 150.745 0.845 154.220 ;
        RECT 0.155 115.135 0.845 119.690 ;
        RECT 0.155 110.315 0.845 113.895 ;
        RECT 0.155 104.990 0.845 108.815 ;
        RECT 0.155 92.280 0.845 100.280 ;
        RECT 0.155 81.280 0.845 89.280 ;
        RECT 0.155 70.280 0.845 78.280 ;
  END 
END PLFILLER1

MACRO PLFILLER01
  CLASS  PAD ;
  FOREIGN PLFILLER01 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.100 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M1 ;
        RECT 0.000 171.175 0.100 172.780 ;
        RECT 0.000 162.720 0.100 170.715 ;
        RECT 0.000 155.725 0.100 161.220 ;
        RECT 0.000 115.135 0.100 154.220 ;
        RECT 0.000 110.315 0.100 113.895 ;
        RECT 0.000 70.000 0.100 108.815 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.100 172.780 ;
        RECT 0.000 162.720 0.100 170.715 ;
        RECT 0.000 155.725 0.100 161.220 ;
        RECT 0.000 150.480 0.100 154.220 ;
        RECT 0.000 137.395 0.100 147.565 ;
        RECT 0.000 127.100 0.100 134.395 ;
        RECT 0.000 121.860 0.100 124.100 ;
        RECT 0.000 115.135 0.100 119.705 ;
        RECT 0.000 110.315 0.100 113.895 ;
        RECT 0.000 97.700 0.100 108.815 ;
        RECT 0.000 86.640 0.100 94.700 ;
        RECT 0.000 75.630 0.100 83.640 ;
        RECT 0.000 70.000 0.100 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.100 172.780 ;
        RECT 0.000 162.720 0.100 170.715 ;
        RECT 0.000 155.725 0.100 161.220 ;
        RECT 0.000 150.480 0.100 154.220 ;
        RECT 0.000 143.340 0.100 147.565 ;
        RECT 0.000 131.850 0.100 140.340 ;
        RECT 0.000 121.860 0.100 128.850 ;
        RECT 0.000 115.135 0.100 119.705 ;
        RECT 0.000 110.315 0.100 113.895 ;
        RECT 0.000 103.280 0.100 108.815 ;
        RECT 0.000 92.280 0.100 100.280 ;
        RECT 0.000 81.280 0.100 89.280 ;
        RECT 0.000 70.000 0.100 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.100 172.780 ;
        RECT 0.000 162.720 0.100 170.715 ;
        RECT 0.000 155.725 0.100 161.220 ;
        RECT 0.000 150.480 0.100 154.220 ;
        RECT 0.000 143.340 0.100 147.565 ;
        RECT 0.000 131.850 0.100 140.340 ;
        RECT 0.000 121.860 0.100 128.850 ;
        RECT 0.000 115.135 0.100 119.705 ;
        RECT 0.000 110.315 0.100 113.895 ;
        RECT 0.000 103.280 0.100 108.815 ;
        RECT 0.000 92.280 0.100 100.280 ;
        RECT 0.000 81.280 0.100 89.280 ;
        RECT 0.000 70.000 0.100 78.280 ;
  END 
END PLFILLER01

MACRO PLFILLER001
  CLASS  PAD ;
  FOREIGN PLFILLER001 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.010 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M1 ;
        RECT 0.000 171.175 0.010 172.780 ;
        RECT 0.000 162.720 0.010 170.715 ;
        RECT 0.000 155.725 0.010 161.220 ;
        RECT 0.000 115.135 0.010 154.220 ;
        RECT 0.000 110.315 0.010 113.895 ;
        RECT 0.000 70.000 0.010 108.815 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.010 172.780 ;
        RECT 0.000 162.720 0.010 170.715 ;
        RECT 0.000 155.725 0.010 161.220 ;
        RECT 0.000 150.480 0.010 154.220 ;
        RECT 0.000 137.395 0.010 147.565 ;
        RECT 0.000 127.100 0.010 134.395 ;
        RECT 0.000 121.860 0.010 124.100 ;
        RECT 0.000 115.135 0.010 119.705 ;
        RECT 0.000 110.315 0.010 113.895 ;
        RECT 0.000 97.700 0.010 108.815 ;
        RECT 0.000 86.640 0.010 94.700 ;
        RECT 0.000 75.630 0.010 83.640 ;
        RECT 0.000 70.000 0.010 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.010 172.780 ;
        RECT 0.000 162.720 0.010 170.715 ;
        RECT 0.000 155.725 0.010 161.220 ;
        RECT 0.000 150.480 0.010 154.220 ;
        RECT 0.000 143.340 0.010 147.565 ;
        RECT 0.000 131.850 0.010 140.340 ;
        RECT 0.000 121.860 0.010 128.850 ;
        RECT 0.000 115.135 0.010 119.705 ;
        RECT 0.000 110.315 0.010 113.895 ;
        RECT 0.000 103.280 0.010 108.815 ;
        RECT 0.000 92.280 0.010 100.280 ;
        RECT 0.000 81.280 0.010 89.280 ;
        RECT 0.000 70.000 0.010 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.010 172.780 ;
        RECT 0.000 162.720 0.010 170.715 ;
        RECT 0.000 155.725 0.010 161.220 ;
        RECT 0.000 150.480 0.010 154.220 ;
        RECT 0.000 143.340 0.010 147.565 ;
        RECT 0.000 131.850 0.010 140.340 ;
        RECT 0.000 121.860 0.010 128.850 ;
        RECT 0.000 115.135 0.010 119.705 ;
        RECT 0.000 110.315 0.010 113.895 ;
        RECT 0.000 103.280 0.010 108.815 ;
        RECT 0.000 92.280 0.010 100.280 ;
        RECT 0.000 81.280 0.010 89.280 ;
        RECT 0.000 70.000 0.010 78.280 ;
  END 
END PLFILLER001

MACRO PLESDCLAMP
  CLASS  PAD ;
  FOREIGN PLESDCLAMP 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 1.100 1.100 68.900 172.900 ;
      LAYER M1 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 0.000 0.400 70.000 0.700 ;
        RECT 0.000 0.400 0.700 2.300 ;
        RECT 69.300 0.400 70.000 2.300 ;
        RECT 0.000 12.300 0.700 13.100 ;
        RECT 69.300 12.300 70.000 13.100 ;
        RECT 0.000 23.100 0.700 23.900 ;
        RECT 69.300 23.100 70.000 23.900 ;
        RECT 0.000 33.900 0.700 37.100 ;
        RECT 69.300 33.900 70.000 37.100 ;
        RECT 0.000 47.100 0.700 47.900 ;
        RECT 69.300 47.100 70.000 47.900 ;
        RECT 0.000 57.900 0.700 58.700 ;
        RECT 69.300 57.900 70.000 58.700 ;
        RECT 0.000 68.700 0.700 70.700 ;
        RECT 69.300 68.700 70.000 70.700 ;
        RECT 0.000 0.400 0.330 108.815 ;
        RECT 69.670 0.400 70.000 108.815 ;
        RECT 69.300 108.450 70.000 108.815 ;
      LAYER M3 ;
        RECT 1.100 1.100 68.900 172.900 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 1.100 1.100 68.900 172.900 ;
  END 
END PLESDCLAMP

MACRO PLCORNER
  CLASS  ENDCAP BOTTOMLEFT ;
  FOREIGN PLCORNER 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 174.000 BY 174.000 ;
  SYMMETRY Y R90  ;
  SITE CornerSite ;
  OBS 
      LAYER M4 ;
        RECT 107.665 0.000 170.335 173.895 ;
        RECT 0.000 107.665 173.895 170.335 ;
        RECT 0.105 0.105 173.895 173.895 ;
      LAYER M1 ;
        RECT 0.090 70.000 174.000 108.815 ;
        RECT 0.090 110.315 174.000 113.895 ;
        RECT 0.090 115.135 174.000 154.220 ;
        RECT 0.090 155.725 174.000 161.220 ;
        RECT 0.090 162.720 174.000 170.715 ;
        RECT 0.090 171.175 174.000 172.780 ;
        RECT 0.090 0.090 173.910 173.910 ;
        RECT 70.000 0.090 108.815 174.000 ;
        RECT 110.315 0.090 113.895 174.000 ;
        RECT 115.135 0.090 154.220 174.000 ;
        RECT 155.725 0.090 161.220 174.000 ;
        RECT 162.720 0.090 170.715 174.000 ;
        RECT 171.175 0.090 172.780 174.000 ;
      LAYER M3 ;
        RECT 107.665 0.000 170.335 173.895 ;
        RECT 0.000 107.665 173.895 170.335 ;
        RECT 0.105 0.105 173.895 173.895 ;
      LAYER M6 ;
        RECT 162.720 0.000 170.335 174.000 ;
        RECT 107.665 0.000 170.335 173.895 ;
        RECT 0.105 70.000 174.000 72.630 ;
        RECT 0.105 75.630 174.000 83.640 ;
        RECT 0.105 86.640 174.000 94.700 ;
        RECT 0.105 97.700 174.000 108.815 ;
        RECT 0.000 107.665 174.000 108.815 ;
        RECT 0.000 110.315 174.000 113.895 ;
        RECT 0.000 115.135 174.000 119.705 ;
        RECT 0.000 121.860 174.000 124.100 ;
        RECT 0.000 127.100 174.000 134.395 ;
        RECT 0.000 137.395 174.000 147.565 ;
        RECT 0.000 150.480 174.000 154.220 ;
        RECT 0.000 155.725 174.000 161.220 ;
        RECT 0.000 107.665 173.895 170.335 ;
        RECT 0.000 162.720 174.000 170.335 ;
        RECT 0.105 162.720 174.000 170.715 ;
        RECT 0.105 171.175 174.000 172.780 ;
        RECT 0.105 0.105 173.895 173.895 ;
        RECT 70.000 0.105 72.630 174.000 ;
        RECT 75.630 0.105 83.640 174.000 ;
        RECT 86.640 0.105 94.700 174.000 ;
        RECT 107.665 0.000 108.035 174.000 ;
        RECT 96.920 0.105 108.035 174.000 ;
        RECT 110.315 0.000 113.895 174.000 ;
        RECT 115.135 0.000 119.705 174.000 ;
        RECT 121.860 0.000 124.100 174.000 ;
        RECT 127.100 0.000 134.395 174.000 ;
        RECT 137.395 0.000 147.565 174.000 ;
        RECT 150.480 0.000 154.220 174.000 ;
        RECT 155.725 0.000 161.220 174.000 ;
        RECT 162.720 0.105 170.715 174.000 ;
        RECT 171.175 0.105 172.780 174.000 ;
      LAYER M5 ;
        RECT 162.720 0.000 170.335 174.000 ;
        RECT 107.665 0.000 170.335 173.895 ;
        RECT 0.105 70.000 174.000 78.280 ;
        RECT 0.105 81.280 174.000 89.280 ;
        RECT 0.105 92.280 174.000 100.280 ;
        RECT 0.105 103.280 174.000 108.815 ;
        RECT 0.000 107.665 174.000 108.815 ;
        RECT 0.000 110.315 174.000 113.895 ;
        RECT 0.000 115.135 174.000 119.705 ;
        RECT 0.000 121.860 174.000 128.850 ;
        RECT 0.000 131.850 174.000 140.340 ;
        RECT 0.000 143.340 174.000 147.565 ;
        RECT 0.000 150.480 174.000 154.220 ;
        RECT 0.000 155.725 174.000 161.220 ;
        RECT 0.000 107.665 173.895 170.335 ;
        RECT 0.000 162.720 174.000 170.335 ;
        RECT 0.105 162.720 174.000 170.715 ;
        RECT 0.105 171.175 174.000 172.780 ;
        RECT 0.105 0.105 173.895 173.895 ;
        RECT 70.000 0.105 78.280 174.000 ;
        RECT 81.280 0.105 89.280 174.000 ;
        RECT 92.280 0.105 100.280 174.000 ;
        RECT 107.665 0.000 108.815 174.000 ;
        RECT 103.280 0.105 108.815 174.000 ;
        RECT 110.315 0.000 113.895 174.000 ;
        RECT 115.135 0.000 119.705 174.000 ;
        RECT 121.860 0.000 128.850 174.000 ;
        RECT 131.850 0.000 140.340 174.000 ;
        RECT 143.340 0.000 147.565 174.000 ;
        RECT 150.480 0.000 154.220 174.000 ;
        RECT 155.725 0.000 161.220 174.000 ;
        RECT 162.720 0.105 170.715 174.000 ;
        RECT 171.175 0.105 172.780 174.000 ;
      LAYER M7 ;
        RECT 162.720 0.000 170.335 174.000 ;
        RECT 107.665 0.000 170.335 173.770 ;
        RECT 0.230 70.000 174.000 78.280 ;
        RECT 0.230 81.280 174.000 89.280 ;
        RECT 0.230 92.280 174.000 100.280 ;
        RECT 0.230 103.280 174.000 108.815 ;
        RECT 0.000 107.665 174.000 108.815 ;
        RECT 0.000 110.315 174.000 113.895 ;
        RECT 0.000 115.135 174.000 119.705 ;
        RECT 0.000 121.860 174.000 128.850 ;
        RECT 0.000 131.850 174.000 140.340 ;
        RECT 0.000 143.340 174.000 147.565 ;
        RECT 0.000 150.480 174.000 154.220 ;
        RECT 0.000 155.725 174.000 161.220 ;
        RECT 0.000 107.665 173.770 170.335 ;
        RECT 0.000 162.720 174.000 170.335 ;
        RECT 0.230 162.720 174.000 170.715 ;
        RECT 0.230 171.175 174.000 172.780 ;
        RECT 0.230 0.230 173.770 173.770 ;
        RECT 70.000 0.230 78.280 174.000 ;
        RECT 81.280 0.230 89.280 174.000 ;
        RECT 92.280 0.230 100.280 174.000 ;
        RECT 107.665 0.000 108.815 174.000 ;
        RECT 103.280 0.230 108.815 174.000 ;
        RECT 110.315 0.000 113.895 174.000 ;
        RECT 115.135 0.000 119.705 174.000 ;
        RECT 121.860 0.000 128.850 174.000 ;
        RECT 131.850 0.000 140.340 174.000 ;
        RECT 143.340 0.000 147.565 174.000 ;
        RECT 150.480 0.000 154.220 174.000 ;
        RECT 155.725 0.000 161.220 174.000 ;
        RECT 162.720 0.230 170.715 174.000 ;
        RECT 171.175 0.230 172.780 174.000 ;
      LAYER M2 ;
        RECT 107.665 0.000 170.335 173.895 ;
        RECT 0.000 107.665 173.895 170.335 ;
        RECT 0.105 0.105 173.895 173.895 ;
        RECT 110.315 0.000 113.895 173.900 ;
  END 
END PLCORNER

MACRO PLBIAR
  CLASS  PAD ;
  FOREIGN PLBIAR 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
    END
  END P
  PIN AI
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V6 ;
        RECT 4.310 173.515 4.670 173.875 ;
        RECT 5.020 173.515 5.380 173.875 ;
        RECT 5.730 173.515 6.090 173.875 ;
        RECT 6.440 173.515 6.800 173.875 ;
        RECT 7.150 173.515 7.510 173.875 ;
        RECT 7.860 173.515 8.220 173.875 ;
        RECT 8.570 173.515 8.930 173.875 ;
        RECT 9.280 173.515 9.640 173.875 ;
        RECT 9.990 173.515 10.350 173.875 ;
        RECT 10.700 173.515 11.060 173.875 ;
        RECT 11.410 173.515 11.770 173.875 ;
        RECT 12.120 173.515 12.480 173.875 ;
        RECT 12.830 173.515 13.190 173.875 ;
        RECT 13.540 173.515 13.900 173.875 ;
        RECT 14.250 173.515 14.610 173.875 ;
        RECT 14.960 173.515 15.320 173.875 ;
        RECT 15.670 173.515 16.030 173.875 ;
        RECT 16.380 173.515 16.740 173.875 ;
        RECT 17.090 173.515 17.450 173.875 ;
        RECT 17.800 173.515 18.160 173.875 ;
        RECT 18.510 173.515 18.870 173.875 ;
        RECT 19.220 173.515 19.580 173.875 ;
        RECT 19.930 173.515 20.290 173.875 ;
        RECT 20.640 173.515 21.000 173.875 ;
        RECT 21.350 173.515 21.710 173.875 ;
        RECT 22.060 173.515 22.420 173.875 ;
        RECT 22.770 173.515 23.130 173.875 ;
        RECT 23.480 173.515 23.840 173.875 ;
        RECT 24.190 173.515 24.550 173.875 ;
        RECT 24.900 173.515 25.260 173.875 ;
        RECT 25.610 173.515 25.970 173.875 ;
        RECT 26.320 173.515 26.680 173.875 ;
        RECT 27.030 173.515 27.390 173.875 ;
        RECT 27.740 173.515 28.100 173.875 ;
        RECT 28.450 173.515 28.810 173.875 ;
        RECT 29.160 173.515 29.520 173.875 ;
        RECT 29.870 173.515 30.230 173.875 ;
        RECT 30.580 173.515 30.940 173.875 ;
        RECT 31.290 173.515 31.650 173.875 ;
        RECT 32.000 173.515 32.360 173.875 ;
        RECT 32.710 173.515 33.070 173.875 ;
        RECT 33.420 173.515 33.780 173.875 ;
        RECT 34.130 173.515 34.490 173.875 ;
        RECT 34.840 173.515 35.200 173.875 ;
        RECT 35.550 173.515 35.910 173.875 ;
        RECT 36.260 173.515 36.620 173.875 ;
        RECT 36.970 173.515 37.330 173.875 ;
        RECT 37.680 173.515 38.040 173.875 ;
        RECT 38.390 173.515 38.750 173.875 ;
        RECT 39.100 173.515 39.460 173.875 ;
        RECT 39.810 173.515 40.170 173.875 ;
        RECT 40.520 173.515 40.880 173.875 ;
        RECT 41.230 173.515 41.590 173.875 ;
        RECT 41.940 173.515 42.300 173.875 ;
        RECT 42.650 173.515 43.010 173.875 ;
        RECT 43.360 173.515 43.720 173.875 ;
        RECT 44.070 173.515 44.430 173.875 ;
        RECT 44.780 173.515 45.140 173.875 ;
        RECT 45.490 173.515 45.850 173.875 ;
        RECT 46.200 173.515 46.560 173.875 ;
        RECT 46.910 173.515 47.270 173.875 ;
        RECT 47.620 173.515 47.980 173.875 ;
        RECT 48.330 173.515 48.690 173.875 ;
        RECT 49.040 173.515 49.400 173.875 ;
        RECT 49.750 173.515 50.110 173.875 ;
        RECT 50.460 173.515 50.820 173.875 ;
        RECT 51.170 173.515 51.530 173.875 ;
        RECT 51.880 173.515 52.240 173.875 ;
        RECT 52.590 173.515 52.950 173.875 ;
        RECT 53.300 173.515 53.660 173.875 ;
        RECT 54.010 173.515 54.370 173.875 ;
        RECT 54.720 173.515 55.080 173.875 ;
        RECT 55.430 173.515 55.790 173.875 ;
        RECT 56.140 173.515 56.500 173.875 ;
        RECT 56.850 173.515 57.210 173.875 ;
        RECT 57.560 173.515 57.920 173.875 ;
        RECT 58.270 173.515 58.630 173.875 ;
        RECT 58.980 173.515 59.340 173.875 ;
        RECT 59.690 173.515 60.050 173.875 ;
        RECT 60.400 173.515 60.760 173.875 ;
        RECT 61.110 173.515 61.470 173.875 ;
        RECT 61.820 173.515 62.180 173.875 ;
        RECT 62.530 173.515 62.890 173.875 ;
        RECT 63.240 173.515 63.600 173.875 ;
        RECT 63.950 173.515 64.310 173.875 ;
        RECT 64.660 173.515 65.020 173.875 ;
        RECT 65.370 173.515 65.730 173.875 ;
      LAYER M4 ;
        RECT 3.510 173.300 66.490 174.000 ;
      LAYER V3 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M3 ;
        RECT 3.510 173.300 66.490 174.000 ;
      LAYER V2 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M2 ;
        RECT 3.510 173.300 66.490 174.000 ;
      LAYER V1 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M1 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER M6 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V5 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M5 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V4 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
    END
  END AI
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 168.090 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 152.430 69.840 154.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
        RECT 69.300 105.215 69.840 108.815 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 162.720 69.845 168.090 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 168.090 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 152.430 69.840 154.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
        RECT 69.300 105.215 69.840 108.815 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 162.720 69.845 168.090 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 168.090 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.300 152.430 69.840 154.220 ;
        RECT 69.300 110.315 69.840 113.895 ;
        RECT 69.300 105.215 69.840 108.815 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 162.720 69.845 168.090 ;
  END 
END PLBIAR

MACRO PLBIA
  CLASS  PAD ;
  FOREIGN PLBIA 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V6 ;
        RECT 4.310 173.515 4.670 173.875 ;
        RECT 5.020 173.515 5.380 173.875 ;
        RECT 5.730 173.515 6.090 173.875 ;
        RECT 6.440 173.515 6.800 173.875 ;
        RECT 7.150 173.515 7.510 173.875 ;
        RECT 7.860 173.515 8.220 173.875 ;
        RECT 8.570 173.515 8.930 173.875 ;
        RECT 9.280 173.515 9.640 173.875 ;
        RECT 9.990 173.515 10.350 173.875 ;
        RECT 10.700 173.515 11.060 173.875 ;
        RECT 11.410 173.515 11.770 173.875 ;
        RECT 12.120 173.515 12.480 173.875 ;
        RECT 12.830 173.515 13.190 173.875 ;
        RECT 13.540 173.515 13.900 173.875 ;
        RECT 14.250 173.515 14.610 173.875 ;
        RECT 14.960 173.515 15.320 173.875 ;
        RECT 15.670 173.515 16.030 173.875 ;
        RECT 16.380 173.515 16.740 173.875 ;
        RECT 17.090 173.515 17.450 173.875 ;
        RECT 17.800 173.515 18.160 173.875 ;
        RECT 18.510 173.515 18.870 173.875 ;
        RECT 19.220 173.515 19.580 173.875 ;
        RECT 19.930 173.515 20.290 173.875 ;
        RECT 20.640 173.515 21.000 173.875 ;
        RECT 21.350 173.515 21.710 173.875 ;
        RECT 22.060 173.515 22.420 173.875 ;
        RECT 22.770 173.515 23.130 173.875 ;
        RECT 23.480 173.515 23.840 173.875 ;
        RECT 24.190 173.515 24.550 173.875 ;
        RECT 24.900 173.515 25.260 173.875 ;
        RECT 25.610 173.515 25.970 173.875 ;
        RECT 26.320 173.515 26.680 173.875 ;
        RECT 27.030 173.515 27.390 173.875 ;
        RECT 27.740 173.515 28.100 173.875 ;
        RECT 28.450 173.515 28.810 173.875 ;
        RECT 29.160 173.515 29.520 173.875 ;
        RECT 29.870 173.515 30.230 173.875 ;
        RECT 30.580 173.515 30.940 173.875 ;
        RECT 31.290 173.515 31.650 173.875 ;
        RECT 32.000 173.515 32.360 173.875 ;
        RECT 32.710 173.515 33.070 173.875 ;
        RECT 33.420 173.515 33.780 173.875 ;
        RECT 34.130 173.515 34.490 173.875 ;
        RECT 34.840 173.515 35.200 173.875 ;
        RECT 35.550 173.515 35.910 173.875 ;
        RECT 36.260 173.515 36.620 173.875 ;
        RECT 36.970 173.515 37.330 173.875 ;
        RECT 37.680 173.515 38.040 173.875 ;
        RECT 38.390 173.515 38.750 173.875 ;
        RECT 39.100 173.515 39.460 173.875 ;
        RECT 39.810 173.515 40.170 173.875 ;
        RECT 40.520 173.515 40.880 173.875 ;
        RECT 41.230 173.515 41.590 173.875 ;
        RECT 41.940 173.515 42.300 173.875 ;
        RECT 42.650 173.515 43.010 173.875 ;
        RECT 43.360 173.515 43.720 173.875 ;
        RECT 44.070 173.515 44.430 173.875 ;
        RECT 44.780 173.515 45.140 173.875 ;
        RECT 45.490 173.515 45.850 173.875 ;
        RECT 46.200 173.515 46.560 173.875 ;
        RECT 46.910 173.515 47.270 173.875 ;
        RECT 47.620 173.515 47.980 173.875 ;
        RECT 48.330 173.515 48.690 173.875 ;
        RECT 49.040 173.515 49.400 173.875 ;
        RECT 49.750 173.515 50.110 173.875 ;
        RECT 50.460 173.515 50.820 173.875 ;
        RECT 51.170 173.515 51.530 173.875 ;
        RECT 51.880 173.515 52.240 173.875 ;
        RECT 52.590 173.515 52.950 173.875 ;
        RECT 53.300 173.515 53.660 173.875 ;
        RECT 54.010 173.515 54.370 173.875 ;
        RECT 54.720 173.515 55.080 173.875 ;
        RECT 55.430 173.515 55.790 173.875 ;
        RECT 56.140 173.515 56.500 173.875 ;
        RECT 56.850 173.515 57.210 173.875 ;
        RECT 57.560 173.515 57.920 173.875 ;
        RECT 58.270 173.515 58.630 173.875 ;
        RECT 58.980 173.515 59.340 173.875 ;
        RECT 59.690 173.515 60.050 173.875 ;
        RECT 60.400 173.515 60.760 173.875 ;
        RECT 61.110 173.515 61.470 173.875 ;
        RECT 61.820 173.515 62.180 173.875 ;
        RECT 62.530 173.515 62.890 173.875 ;
        RECT 63.240 173.515 63.600 173.875 ;
        RECT 63.950 173.515 64.310 173.875 ;
        RECT 64.660 173.515 65.020 173.875 ;
        RECT 65.370 173.515 65.730 173.875 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V3 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.300 66.490 174.000 ;
      LAYER V2 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.300 66.490 174.000 ;
      LAYER V1 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M1 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V5 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
        RECT 3.510 173.380 66.490 174.000 ;
      LAYER V4 ;
        RECT 4.360 173.800 4.550 173.990 ;
        RECT 4.360 173.390 4.550 173.580 ;
        RECT 4.770 173.800 4.960 173.990 ;
        RECT 4.770 173.390 4.960 173.580 ;
        RECT 5.180 173.800 5.370 173.990 ;
        RECT 5.180 173.390 5.370 173.580 ;
        RECT 5.590 173.800 5.780 173.990 ;
        RECT 5.590 173.390 5.780 173.580 ;
        RECT 6.000 173.800 6.190 173.990 ;
        RECT 6.000 173.390 6.190 173.580 ;
        RECT 6.410 173.800 6.600 173.990 ;
        RECT 6.410 173.390 6.600 173.580 ;
        RECT 6.820 173.800 7.010 173.990 ;
        RECT 6.820 173.390 7.010 173.580 ;
        RECT 7.230 173.800 7.420 173.990 ;
        RECT 7.230 173.390 7.420 173.580 ;
        RECT 7.640 173.800 7.830 173.990 ;
        RECT 7.640 173.390 7.830 173.580 ;
        RECT 8.050 173.800 8.240 173.990 ;
        RECT 8.050 173.390 8.240 173.580 ;
        RECT 8.460 173.800 8.650 173.990 ;
        RECT 8.460 173.390 8.650 173.580 ;
        RECT 8.870 173.800 9.060 173.990 ;
        RECT 8.870 173.390 9.060 173.580 ;
        RECT 9.280 173.800 9.470 173.990 ;
        RECT 9.280 173.390 9.470 173.580 ;
        RECT 9.690 173.800 9.880 173.990 ;
        RECT 9.690 173.390 9.880 173.580 ;
        RECT 10.100 173.800 10.290 173.990 ;
        RECT 10.100 173.390 10.290 173.580 ;
        RECT 10.510 173.800 10.700 173.990 ;
        RECT 10.510 173.390 10.700 173.580 ;
        RECT 10.920 173.800 11.110 173.990 ;
        RECT 10.920 173.390 11.110 173.580 ;
        RECT 11.330 173.800 11.520 173.990 ;
        RECT 11.330 173.390 11.520 173.580 ;
        RECT 11.740 173.800 11.930 173.990 ;
        RECT 11.740 173.390 11.930 173.580 ;
        RECT 12.150 173.800 12.340 173.990 ;
        RECT 12.150 173.390 12.340 173.580 ;
        RECT 12.560 173.800 12.750 173.990 ;
        RECT 12.560 173.390 12.750 173.580 ;
        RECT 12.970 173.800 13.160 173.990 ;
        RECT 12.970 173.390 13.160 173.580 ;
        RECT 13.380 173.800 13.570 173.990 ;
        RECT 13.380 173.390 13.570 173.580 ;
        RECT 13.790 173.800 13.980 173.990 ;
        RECT 13.790 173.390 13.980 173.580 ;
        RECT 14.200 173.800 14.390 173.990 ;
        RECT 14.200 173.390 14.390 173.580 ;
        RECT 14.610 173.800 14.800 173.990 ;
        RECT 14.610 173.390 14.800 173.580 ;
        RECT 15.020 173.800 15.210 173.990 ;
        RECT 15.020 173.390 15.210 173.580 ;
        RECT 15.430 173.800 15.620 173.990 ;
        RECT 15.430 173.390 15.620 173.580 ;
        RECT 15.840 173.800 16.030 173.990 ;
        RECT 15.840 173.390 16.030 173.580 ;
        RECT 16.250 173.800 16.440 173.990 ;
        RECT 16.250 173.390 16.440 173.580 ;
        RECT 16.660 173.800 16.850 173.990 ;
        RECT 16.660 173.390 16.850 173.580 ;
        RECT 17.070 173.800 17.260 173.990 ;
        RECT 17.070 173.390 17.260 173.580 ;
        RECT 17.480 173.800 17.670 173.990 ;
        RECT 17.480 173.390 17.670 173.580 ;
        RECT 17.890 173.800 18.080 173.990 ;
        RECT 17.890 173.390 18.080 173.580 ;
        RECT 18.300 173.800 18.490 173.990 ;
        RECT 18.300 173.390 18.490 173.580 ;
        RECT 18.710 173.800 18.900 173.990 ;
        RECT 18.710 173.390 18.900 173.580 ;
        RECT 19.120 173.800 19.310 173.990 ;
        RECT 19.120 173.390 19.310 173.580 ;
        RECT 19.530 173.800 19.720 173.990 ;
        RECT 19.530 173.390 19.720 173.580 ;
        RECT 19.940 173.800 20.130 173.990 ;
        RECT 19.940 173.390 20.130 173.580 ;
        RECT 20.350 173.800 20.540 173.990 ;
        RECT 20.350 173.390 20.540 173.580 ;
        RECT 20.760 173.800 20.950 173.990 ;
        RECT 20.760 173.390 20.950 173.580 ;
        RECT 21.170 173.800 21.360 173.990 ;
        RECT 21.170 173.390 21.360 173.580 ;
        RECT 21.580 173.800 21.770 173.990 ;
        RECT 21.580 173.390 21.770 173.580 ;
        RECT 21.990 173.800 22.180 173.990 ;
        RECT 21.990 173.390 22.180 173.580 ;
        RECT 22.400 173.800 22.590 173.990 ;
        RECT 22.400 173.390 22.590 173.580 ;
        RECT 22.810 173.800 23.000 173.990 ;
        RECT 22.810 173.390 23.000 173.580 ;
        RECT 23.220 173.800 23.410 173.990 ;
        RECT 23.220 173.390 23.410 173.580 ;
        RECT 23.630 173.800 23.820 173.990 ;
        RECT 23.630 173.390 23.820 173.580 ;
        RECT 24.040 173.800 24.230 173.990 ;
        RECT 24.040 173.390 24.230 173.580 ;
        RECT 24.450 173.800 24.640 173.990 ;
        RECT 24.450 173.390 24.640 173.580 ;
        RECT 24.860 173.800 25.050 173.990 ;
        RECT 24.860 173.390 25.050 173.580 ;
        RECT 25.270 173.800 25.460 173.990 ;
        RECT 25.270 173.390 25.460 173.580 ;
        RECT 25.680 173.800 25.870 173.990 ;
        RECT 25.680 173.390 25.870 173.580 ;
        RECT 26.090 173.800 26.280 173.990 ;
        RECT 26.090 173.390 26.280 173.580 ;
        RECT 26.500 173.800 26.690 173.990 ;
        RECT 26.500 173.390 26.690 173.580 ;
        RECT 26.910 173.800 27.100 173.990 ;
        RECT 26.910 173.390 27.100 173.580 ;
        RECT 27.320 173.800 27.510 173.990 ;
        RECT 27.320 173.390 27.510 173.580 ;
        RECT 27.730 173.800 27.920 173.990 ;
        RECT 27.730 173.390 27.920 173.580 ;
        RECT 28.140 173.800 28.330 173.990 ;
        RECT 28.140 173.390 28.330 173.580 ;
        RECT 28.550 173.800 28.740 173.990 ;
        RECT 28.550 173.390 28.740 173.580 ;
        RECT 28.960 173.800 29.150 173.990 ;
        RECT 28.960 173.390 29.150 173.580 ;
        RECT 29.370 173.800 29.560 173.990 ;
        RECT 29.370 173.390 29.560 173.580 ;
        RECT 29.780 173.800 29.970 173.990 ;
        RECT 29.780 173.390 29.970 173.580 ;
        RECT 30.190 173.800 30.380 173.990 ;
        RECT 30.190 173.390 30.380 173.580 ;
        RECT 30.600 173.800 30.790 173.990 ;
        RECT 30.600 173.390 30.790 173.580 ;
        RECT 31.010 173.800 31.200 173.990 ;
        RECT 31.010 173.390 31.200 173.580 ;
        RECT 31.420 173.800 31.610 173.990 ;
        RECT 31.420 173.390 31.610 173.580 ;
        RECT 31.830 173.800 32.020 173.990 ;
        RECT 31.830 173.390 32.020 173.580 ;
        RECT 32.240 173.800 32.430 173.990 ;
        RECT 32.240 173.390 32.430 173.580 ;
        RECT 32.650 173.800 32.840 173.990 ;
        RECT 32.650 173.390 32.840 173.580 ;
        RECT 33.060 173.800 33.250 173.990 ;
        RECT 33.060 173.390 33.250 173.580 ;
        RECT 33.470 173.800 33.660 173.990 ;
        RECT 33.470 173.390 33.660 173.580 ;
        RECT 33.880 173.800 34.070 173.990 ;
        RECT 33.880 173.390 34.070 173.580 ;
        RECT 34.290 173.800 34.480 173.990 ;
        RECT 34.290 173.390 34.480 173.580 ;
        RECT 34.700 173.800 34.890 173.990 ;
        RECT 34.700 173.390 34.890 173.580 ;
        RECT 35.110 173.800 35.300 173.990 ;
        RECT 35.110 173.390 35.300 173.580 ;
        RECT 35.520 173.800 35.710 173.990 ;
        RECT 35.520 173.390 35.710 173.580 ;
        RECT 35.930 173.800 36.120 173.990 ;
        RECT 35.930 173.390 36.120 173.580 ;
        RECT 36.340 173.800 36.530 173.990 ;
        RECT 36.340 173.390 36.530 173.580 ;
        RECT 36.750 173.800 36.940 173.990 ;
        RECT 36.750 173.390 36.940 173.580 ;
        RECT 37.160 173.800 37.350 173.990 ;
        RECT 37.160 173.390 37.350 173.580 ;
        RECT 37.570 173.800 37.760 173.990 ;
        RECT 37.570 173.390 37.760 173.580 ;
        RECT 37.980 173.800 38.170 173.990 ;
        RECT 37.980 173.390 38.170 173.580 ;
        RECT 38.390 173.800 38.580 173.990 ;
        RECT 38.390 173.390 38.580 173.580 ;
        RECT 38.800 173.800 38.990 173.990 ;
        RECT 38.800 173.390 38.990 173.580 ;
        RECT 39.210 173.800 39.400 173.990 ;
        RECT 39.210 173.390 39.400 173.580 ;
        RECT 39.620 173.800 39.810 173.990 ;
        RECT 39.620 173.390 39.810 173.580 ;
        RECT 40.030 173.800 40.220 173.990 ;
        RECT 40.030 173.390 40.220 173.580 ;
        RECT 40.440 173.800 40.630 173.990 ;
        RECT 40.440 173.390 40.630 173.580 ;
        RECT 40.850 173.800 41.040 173.990 ;
        RECT 40.850 173.390 41.040 173.580 ;
        RECT 41.260 173.800 41.450 173.990 ;
        RECT 41.260 173.390 41.450 173.580 ;
        RECT 41.670 173.800 41.860 173.990 ;
        RECT 41.670 173.390 41.860 173.580 ;
        RECT 42.080 173.800 42.270 173.990 ;
        RECT 42.080 173.390 42.270 173.580 ;
        RECT 42.490 173.800 42.680 173.990 ;
        RECT 42.490 173.390 42.680 173.580 ;
        RECT 42.900 173.800 43.090 173.990 ;
        RECT 42.900 173.390 43.090 173.580 ;
        RECT 43.310 173.800 43.500 173.990 ;
        RECT 43.310 173.390 43.500 173.580 ;
        RECT 43.720 173.800 43.910 173.990 ;
        RECT 43.720 173.390 43.910 173.580 ;
        RECT 44.130 173.800 44.320 173.990 ;
        RECT 44.130 173.390 44.320 173.580 ;
        RECT 44.540 173.800 44.730 173.990 ;
        RECT 44.540 173.390 44.730 173.580 ;
        RECT 44.950 173.800 45.140 173.990 ;
        RECT 44.950 173.390 45.140 173.580 ;
        RECT 45.360 173.800 45.550 173.990 ;
        RECT 45.360 173.390 45.550 173.580 ;
        RECT 45.770 173.800 45.960 173.990 ;
        RECT 45.770 173.390 45.960 173.580 ;
        RECT 46.180 173.800 46.370 173.990 ;
        RECT 46.180 173.390 46.370 173.580 ;
        RECT 46.590 173.800 46.780 173.990 ;
        RECT 46.590 173.390 46.780 173.580 ;
        RECT 47.000 173.800 47.190 173.990 ;
        RECT 47.000 173.390 47.190 173.580 ;
        RECT 47.410 173.800 47.600 173.990 ;
        RECT 47.410 173.390 47.600 173.580 ;
        RECT 47.820 173.800 48.010 173.990 ;
        RECT 47.820 173.390 48.010 173.580 ;
        RECT 48.230 173.800 48.420 173.990 ;
        RECT 48.230 173.390 48.420 173.580 ;
        RECT 48.640 173.800 48.830 173.990 ;
        RECT 48.640 173.390 48.830 173.580 ;
        RECT 49.050 173.800 49.240 173.990 ;
        RECT 49.050 173.390 49.240 173.580 ;
        RECT 49.460 173.800 49.650 173.990 ;
        RECT 49.460 173.390 49.650 173.580 ;
        RECT 49.870 173.800 50.060 173.990 ;
        RECT 49.870 173.390 50.060 173.580 ;
        RECT 50.280 173.800 50.470 173.990 ;
        RECT 50.280 173.390 50.470 173.580 ;
        RECT 50.690 173.800 50.880 173.990 ;
        RECT 50.690 173.390 50.880 173.580 ;
        RECT 51.100 173.800 51.290 173.990 ;
        RECT 51.100 173.390 51.290 173.580 ;
        RECT 51.510 173.800 51.700 173.990 ;
        RECT 51.510 173.390 51.700 173.580 ;
        RECT 51.920 173.800 52.110 173.990 ;
        RECT 51.920 173.390 52.110 173.580 ;
        RECT 52.330 173.800 52.520 173.990 ;
        RECT 52.330 173.390 52.520 173.580 ;
        RECT 52.740 173.800 52.930 173.990 ;
        RECT 52.740 173.390 52.930 173.580 ;
        RECT 53.150 173.800 53.340 173.990 ;
        RECT 53.150 173.390 53.340 173.580 ;
        RECT 53.560 173.800 53.750 173.990 ;
        RECT 53.560 173.390 53.750 173.580 ;
        RECT 53.970 173.800 54.160 173.990 ;
        RECT 53.970 173.390 54.160 173.580 ;
        RECT 54.380 173.800 54.570 173.990 ;
        RECT 54.380 173.390 54.570 173.580 ;
        RECT 54.790 173.800 54.980 173.990 ;
        RECT 54.790 173.390 54.980 173.580 ;
        RECT 55.200 173.800 55.390 173.990 ;
        RECT 55.200 173.390 55.390 173.580 ;
        RECT 55.610 173.800 55.800 173.990 ;
        RECT 55.610 173.390 55.800 173.580 ;
        RECT 56.020 173.800 56.210 173.990 ;
        RECT 56.020 173.390 56.210 173.580 ;
        RECT 56.430 173.800 56.620 173.990 ;
        RECT 56.430 173.390 56.620 173.580 ;
        RECT 56.840 173.800 57.030 173.990 ;
        RECT 56.840 173.390 57.030 173.580 ;
        RECT 57.250 173.800 57.440 173.990 ;
        RECT 57.250 173.390 57.440 173.580 ;
        RECT 57.660 173.800 57.850 173.990 ;
        RECT 57.660 173.390 57.850 173.580 ;
        RECT 58.070 173.800 58.260 173.990 ;
        RECT 58.070 173.390 58.260 173.580 ;
        RECT 58.480 173.800 58.670 173.990 ;
        RECT 58.480 173.390 58.670 173.580 ;
        RECT 58.890 173.800 59.080 173.990 ;
        RECT 58.890 173.390 59.080 173.580 ;
        RECT 59.300 173.800 59.490 173.990 ;
        RECT 59.300 173.390 59.490 173.580 ;
        RECT 59.710 173.800 59.900 173.990 ;
        RECT 59.710 173.390 59.900 173.580 ;
        RECT 60.120 173.800 60.310 173.990 ;
        RECT 60.120 173.390 60.310 173.580 ;
        RECT 60.530 173.800 60.720 173.990 ;
        RECT 60.530 173.390 60.720 173.580 ;
        RECT 60.940 173.800 61.130 173.990 ;
        RECT 60.940 173.390 61.130 173.580 ;
        RECT 61.350 173.800 61.540 173.990 ;
        RECT 61.350 173.390 61.540 173.580 ;
        RECT 61.760 173.800 61.950 173.990 ;
        RECT 61.760 173.390 61.950 173.580 ;
        RECT 62.170 173.800 62.360 173.990 ;
        RECT 62.170 173.390 62.360 173.580 ;
        RECT 62.580 173.800 62.770 173.990 ;
        RECT 62.580 173.390 62.770 173.580 ;
        RECT 62.990 173.800 63.180 173.990 ;
        RECT 62.990 173.390 63.180 173.580 ;
        RECT 63.400 173.800 63.590 173.990 ;
        RECT 63.400 173.390 63.590 173.580 ;
        RECT 63.810 173.800 64.000 173.990 ;
        RECT 63.810 173.390 64.000 173.580 ;
        RECT 64.220 173.800 64.410 173.990 ;
        RECT 64.220 173.390 64.410 173.580 ;
        RECT 64.630 173.800 64.820 173.990 ;
        RECT 64.630 173.390 64.820 173.580 ;
        RECT 65.040 173.800 65.230 173.990 ;
        RECT 65.040 173.390 65.230 173.580 ;
        RECT 65.450 173.800 65.640 173.990 ;
        RECT 65.450 173.390 65.640 173.580 ;
    END
  END P
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.715 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.790 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.895 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.285 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.520 150.720 69.840 154.220 ;
        RECT 69.520 115.135 69.840 119.725 ;
        RECT 69.300 110.315 69.840 113.895 ;
        RECT 69.300 105.215 69.840 108.815 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 162.720 69.845 170.715 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.855 ;
        RECT 69.300 152.430 70.000 152.730 ;
        RECT 69.520 115.135 70.000 154.220 ;
        RECT 69.300 153.920 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.715 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.790 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.895 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.285 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.520 150.720 69.840 154.220 ;
        RECT 69.520 115.135 69.840 119.725 ;
        RECT 69.300 110.315 69.840 113.895 ;
        RECT 69.300 105.215 69.840 108.815 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 162.720 69.845 170.715 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.715 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.790 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.895 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.285 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 155.725 69.840 161.220 ;
        RECT 69.520 150.720 69.840 154.220 ;
        RECT 69.520 115.135 69.840 119.725 ;
        RECT 69.300 110.315 69.840 113.895 ;
        RECT 69.300 105.215 69.840 108.815 ;
        RECT 69.300 92.280 69.840 100.415 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 162.720 69.845 170.715 ;
  END 
END PLBIA

MACRO PLBI24S
  CLASS  PAD ;
  FOREIGN PLBI24S 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V6 ;
        RECT 9.520 173.510 9.880 173.870 ;
      LAYER M4 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V3 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M3 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V2 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M2 ;
        RECT 9.600 173.300 9.800 174.000 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V1 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M1 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER M6 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V5 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M5 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V4 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V6 ;
        RECT 66.240 173.510 66.600 173.870 ;
      LAYER M4 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V3 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M3 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V2 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M2 ;
        RECT 66.320 173.300 66.520 174.000 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V1 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M1 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER M6 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V5 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M5 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V4 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V6 ;
        RECT 21.400 173.510 21.760 173.870 ;
      LAYER M4 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V3 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M3 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V2 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M2 ;
        RECT 21.480 173.300 21.680 174.000 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V1 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M1 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER M6 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V5 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M5 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V4 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V6 ;
        RECT 28.545 173.510 28.905 173.870 ;
      LAYER M4 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V3 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M3 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V2 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M2 ;
        RECT 28.625 173.300 28.825 174.000 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V1 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M1 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER M6 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V5 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M5 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V4 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V6 ;
        RECT 24.395 173.510 24.755 173.870 ;
      LAYER M4 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V3 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M3 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V2 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M2 ;
        RECT 24.475 173.300 24.675 174.000 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V1 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M1 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER M6 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V5 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M5 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V4 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V6 ;
        RECT 17.995 173.510 18.355 173.870 ;
      LAYER M4 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V3 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M3 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V2 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M2 ;
        RECT 18.075 173.300 18.275 174.000 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V1 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M1 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER M6 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V5 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M5 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V4 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V6 ;
        RECT 13.620 173.510 13.980 173.870 ;
      LAYER M4 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V3 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M3 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V2 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M2 ;
        RECT 13.700 173.300 13.900 174.000 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V1 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M1 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER M6 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V5 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M5 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V4 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V6 ;
        RECT 51.035 173.510 51.395 173.870 ;
      LAYER M4 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V3 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M3 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V2 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M2 ;
        RECT 51.115 173.300 51.315 174.000 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V1 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M1 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER M6 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V5 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M5 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V4 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.435 110.315 69.660 113.895 ;
        RECT 69.435 105.235 69.660 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.855 ;
        RECT 69.300 152.430 70.000 152.730 ;
        RECT 69.640 115.135 70.000 154.220 ;
        RECT 69.300 153.920 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.435 110.315 69.660 113.895 ;
        RECT 69.435 105.235 69.660 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 150.095 69.870 150.295 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.415 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.435 110.315 69.660 113.895 ;
        RECT 69.435 105.235 69.660 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 116.210 69.730 153.550 ;
        RECT 69.300 116.345 69.865 153.425 ;
        RECT 69.300 116.340 69.860 153.430 ;
        RECT 69.300 116.330 69.850 153.440 ;
        RECT 69.300 116.320 69.840 153.450 ;
        RECT 69.300 116.310 69.830 153.460 ;
        RECT 69.300 116.300 69.820 153.470 ;
        RECT 69.300 116.290 69.810 153.480 ;
        RECT 69.300 116.280 69.800 153.490 ;
        RECT 69.300 116.270 69.790 153.500 ;
        RECT 69.300 116.260 69.780 153.510 ;
        RECT 69.300 116.250 69.770 153.520 ;
        RECT 69.300 116.240 69.760 153.530 ;
        RECT 69.300 116.230 69.750 153.540 ;
        RECT 69.300 116.220 69.740 153.550 ;
  END 
END PLBI24S

MACRO PLBI24N
  CLASS  PAD ;
  FOREIGN PLBI24N 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V6 ;
        RECT 9.520 173.510 9.880 173.870 ;
      LAYER M4 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V3 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M3 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V2 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M2 ;
        RECT 9.600 173.300 9.800 174.000 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V1 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M1 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER M6 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V5 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M5 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V4 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V6 ;
        RECT 66.240 173.510 66.600 173.870 ;
      LAYER M4 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V3 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M3 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V2 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M2 ;
        RECT 66.320 173.300 66.520 174.000 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V1 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M1 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER M6 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V5 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M5 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V4 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V6 ;
        RECT 21.400 173.510 21.760 173.870 ;
      LAYER M4 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V3 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M3 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V2 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M2 ;
        RECT 21.480 173.300 21.680 174.000 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V1 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M1 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER M6 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V5 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M5 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V4 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V6 ;
        RECT 28.545 173.510 28.905 173.870 ;
      LAYER M4 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V3 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M3 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V2 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M2 ;
        RECT 28.625 173.300 28.825 174.000 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V1 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M1 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER M6 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V5 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M5 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V4 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V6 ;
        RECT 24.395 173.510 24.755 173.870 ;
      LAYER M4 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V3 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M3 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V2 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M2 ;
        RECT 24.475 173.300 24.675 174.000 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V1 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M1 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER M6 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V5 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M5 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V4 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V6 ;
        RECT 17.995 173.510 18.355 173.870 ;
      LAYER M4 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V3 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M3 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V2 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M2 ;
        RECT 18.075 173.300 18.275 174.000 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V1 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M1 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER M6 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V5 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M5 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V4 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V6 ;
        RECT 13.620 173.510 13.980 173.870 ;
      LAYER M4 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V3 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M3 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V2 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M2 ;
        RECT 13.700 173.300 13.900 174.000 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V1 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M1 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER M6 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V5 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M5 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V4 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V6 ;
        RECT 51.035 173.510 51.395 173.870 ;
      LAYER M4 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V3 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M3 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V2 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M2 ;
        RECT 51.115 173.300 51.315 174.000 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V1 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M1 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER M6 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V5 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M5 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V4 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.435 110.315 69.660 113.895 ;
        RECT 69.435 105.235 69.660 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.855 ;
        RECT 69.300 152.430 70.000 152.730 ;
        RECT 69.640 115.135 70.000 154.220 ;
        RECT 69.300 153.920 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.435 110.315 69.660 113.895 ;
        RECT 69.435 105.235 69.660 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 150.095 69.870 150.295 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.415 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.435 110.315 69.660 113.895 ;
        RECT 69.435 105.235 69.660 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 116.210 69.730 153.550 ;
        RECT 69.300 116.345 69.865 153.425 ;
        RECT 69.300 116.340 69.860 153.430 ;
        RECT 69.300 116.330 69.850 153.440 ;
        RECT 69.300 116.320 69.840 153.450 ;
        RECT 69.300 116.310 69.830 153.460 ;
        RECT 69.300 116.300 69.820 153.470 ;
        RECT 69.300 116.290 69.810 153.480 ;
        RECT 69.300 116.280 69.800 153.490 ;
        RECT 69.300 116.270 69.790 153.500 ;
        RECT 69.300 116.260 69.780 153.510 ;
        RECT 69.300 116.250 69.770 153.520 ;
        RECT 69.300 116.240 69.760 153.530 ;
        RECT 69.300 116.230 69.750 153.540 ;
        RECT 69.300 116.220 69.740 153.550 ;
  END 
END PLBI24N

MACRO PLBI24F
  CLASS  PAD ;
  FOREIGN PLBI24F 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V6 ;
        RECT 9.520 173.510 9.880 173.870 ;
      LAYER M4 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V3 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M3 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V2 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M2 ;
        RECT 9.600 173.300 9.800 174.000 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V1 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M1 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER M6 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V5 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M5 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V4 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V6 ;
        RECT 66.240 173.510 66.600 173.870 ;
      LAYER M4 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V3 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M3 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V2 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M2 ;
        RECT 66.320 173.300 66.520 174.000 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V1 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M1 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER M6 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V5 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M5 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V4 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V6 ;
        RECT 21.400 173.510 21.760 173.870 ;
      LAYER M4 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V3 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M3 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V2 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M2 ;
        RECT 21.480 173.300 21.680 174.000 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V1 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M1 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER M6 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V5 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M5 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V4 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V6 ;
        RECT 28.545 173.510 28.905 173.870 ;
      LAYER M4 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V3 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M3 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V2 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M2 ;
        RECT 28.625 173.300 28.825 174.000 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V1 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M1 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER M6 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V5 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M5 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V4 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V6 ;
        RECT 24.395 173.510 24.755 173.870 ;
      LAYER M4 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V3 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M3 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V2 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M2 ;
        RECT 24.475 173.300 24.675 174.000 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V1 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M1 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER M6 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V5 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M5 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V4 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V6 ;
        RECT 17.995 173.510 18.355 173.870 ;
      LAYER M4 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V3 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M3 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V2 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M2 ;
        RECT 18.075 173.300 18.275 174.000 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V1 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M1 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER M6 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V5 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M5 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V4 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V6 ;
        RECT 13.620 173.510 13.980 173.870 ;
      LAYER M4 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V3 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M3 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V2 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M2 ;
        RECT 13.700 173.300 13.900 174.000 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V1 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M1 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER M6 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V5 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M5 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V4 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V6 ;
        RECT 51.035 173.510 51.395 173.870 ;
      LAYER M4 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V3 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M3 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V2 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M2 ;
        RECT 51.115 173.300 51.315 174.000 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V1 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M1 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER M6 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V5 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M5 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V4 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.435 110.315 69.660 113.895 ;
        RECT 69.435 105.235 69.660 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.855 ;
        RECT 69.300 152.430 70.000 152.730 ;
        RECT 69.640 115.135 70.000 154.220 ;
        RECT 69.300 153.920 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.435 110.315 69.660 113.895 ;
        RECT 69.435 105.235 69.660 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 150.095 69.870 150.295 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.415 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.435 110.315 69.660 113.895 ;
        RECT 69.435 105.235 69.660 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 116.210 69.730 153.550 ;
        RECT 69.300 116.345 69.865 153.425 ;
        RECT 69.300 116.340 69.860 153.430 ;
        RECT 69.300 116.330 69.850 153.440 ;
        RECT 69.300 116.320 69.840 153.450 ;
        RECT 69.300 116.310 69.830 153.460 ;
        RECT 69.300 116.300 69.820 153.470 ;
        RECT 69.300 116.290 69.810 153.480 ;
        RECT 69.300 116.280 69.800 153.490 ;
        RECT 69.300 116.270 69.790 153.500 ;
        RECT 69.300 116.260 69.780 153.510 ;
        RECT 69.300 116.250 69.770 153.520 ;
        RECT 69.300 116.240 69.760 153.530 ;
        RECT 69.300 116.230 69.750 153.540 ;
        RECT 69.300 116.220 69.740 153.550 ;
  END 
END PLBI24F

MACRO PLBI16S
  CLASS  PAD ;
  FOREIGN PLBI16S 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V6 ;
        RECT 9.520 173.510 9.880 173.870 ;
      LAYER M4 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V3 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M3 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V2 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M2 ;
        RECT 9.600 173.300 9.800 174.000 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V1 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M1 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER M6 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V5 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M5 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V4 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V6 ;
        RECT 66.240 173.510 66.600 173.870 ;
      LAYER M4 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V3 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M3 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V2 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M2 ;
        RECT 66.320 173.300 66.520 174.000 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V1 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M1 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER M6 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V5 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M5 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V4 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V6 ;
        RECT 21.400 173.510 21.760 173.870 ;
      LAYER M4 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V3 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M3 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V2 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M2 ;
        RECT 21.480 173.300 21.680 174.000 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V1 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M1 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER M6 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V5 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M5 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V4 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V6 ;
        RECT 28.545 173.510 28.905 173.870 ;
      LAYER M4 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V3 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M3 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V2 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M2 ;
        RECT 28.625 173.300 28.825 174.000 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V1 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M1 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER M6 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V5 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M5 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V4 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V6 ;
        RECT 24.395 173.510 24.755 173.870 ;
      LAYER M4 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V3 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M3 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V2 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M2 ;
        RECT 24.475 173.300 24.675 174.000 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V1 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M1 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER M6 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V5 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M5 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V4 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V6 ;
        RECT 17.995 173.510 18.355 173.870 ;
      LAYER M4 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V3 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M3 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V2 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M2 ;
        RECT 18.075 173.300 18.275 174.000 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V1 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M1 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER M6 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V5 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M5 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V4 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V6 ;
        RECT 13.620 173.510 13.980 173.870 ;
      LAYER M4 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V3 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M3 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V2 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M2 ;
        RECT 13.700 173.300 13.900 174.000 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V1 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M1 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER M6 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V5 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M5 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V4 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V6 ;
        RECT 51.035 173.510 51.395 173.870 ;
      LAYER M4 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V3 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M3 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V2 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M2 ;
        RECT 51.115 173.300 51.315 174.000 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V1 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M1 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER M6 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V5 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M5 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V4 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.405 110.315 69.640 113.895 ;
        RECT 69.405 105.235 69.640 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.855 ;
        RECT 69.300 152.430 70.000 152.730 ;
        RECT 69.640 115.135 70.000 154.220 ;
        RECT 69.300 153.920 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.405 110.315 69.640 113.895 ;
        RECT 69.405 105.235 69.640 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 150.095 69.870 150.295 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.415 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.405 110.315 69.640 113.895 ;
        RECT 69.405 105.235 69.640 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 116.210 69.730 153.550 ;
        RECT 69.300 116.345 69.865 153.425 ;
        RECT 69.300 116.340 69.860 153.430 ;
        RECT 69.300 116.330 69.850 153.440 ;
        RECT 69.300 116.320 69.840 153.450 ;
        RECT 69.300 116.310 69.830 153.460 ;
        RECT 69.300 116.300 69.820 153.470 ;
        RECT 69.300 116.290 69.810 153.480 ;
        RECT 69.300 116.280 69.800 153.490 ;
        RECT 69.300 116.270 69.790 153.500 ;
        RECT 69.300 116.260 69.780 153.510 ;
        RECT 69.300 116.250 69.770 153.520 ;
        RECT 69.300 116.240 69.760 153.530 ;
        RECT 69.300 116.230 69.750 153.540 ;
        RECT 69.300 116.220 69.740 153.550 ;
  END 
END PLBI16S

MACRO PLBI16N
  CLASS  PAD ;
  FOREIGN PLBI16N 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V6 ;
        RECT 9.520 173.510 9.880 173.870 ;
      LAYER M4 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V3 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M3 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V2 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M2 ;
        RECT 9.600 173.300 9.800 174.000 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V1 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M1 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER M6 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V5 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M5 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V4 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V6 ;
        RECT 66.240 173.510 66.600 173.870 ;
      LAYER M4 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V3 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M3 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V2 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M2 ;
        RECT 66.320 173.300 66.520 174.000 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V1 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M1 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER M6 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V5 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M5 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V4 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V6 ;
        RECT 21.400 173.510 21.760 173.870 ;
      LAYER M4 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V3 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M3 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V2 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M2 ;
        RECT 21.480 173.300 21.680 174.000 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V1 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M1 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER M6 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V5 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M5 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V4 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V6 ;
        RECT 28.545 173.510 28.905 173.870 ;
      LAYER M4 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V3 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M3 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V2 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M2 ;
        RECT 28.625 173.300 28.825 174.000 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V1 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M1 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER M6 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V5 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M5 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V4 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V6 ;
        RECT 24.395 173.510 24.755 173.870 ;
      LAYER M4 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V3 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M3 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V2 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M2 ;
        RECT 24.475 173.300 24.675 174.000 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V1 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M1 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER M6 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V5 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M5 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V4 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V6 ;
        RECT 17.995 173.510 18.355 173.870 ;
      LAYER M4 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V3 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M3 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V2 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M2 ;
        RECT 18.075 173.300 18.275 174.000 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V1 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M1 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER M6 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V5 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M5 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V4 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V6 ;
        RECT 13.620 173.510 13.980 173.870 ;
      LAYER M4 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V3 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M3 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V2 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M2 ;
        RECT 13.700 173.300 13.900 174.000 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V1 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M1 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER M6 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V5 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M5 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V4 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V6 ;
        RECT 51.035 173.510 51.395 173.870 ;
      LAYER M4 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V3 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M3 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V2 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M2 ;
        RECT 51.115 173.300 51.315 174.000 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V1 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M1 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER M6 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V5 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M5 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V4 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.405 110.315 69.640 113.895 ;
        RECT 69.405 105.235 69.640 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.855 ;
        RECT 69.300 152.430 70.000 152.730 ;
        RECT 69.640 115.135 70.000 154.220 ;
        RECT 69.300 153.920 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.405 110.315 69.640 113.895 ;
        RECT 69.405 105.235 69.640 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 150.095 69.870 150.295 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.415 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.405 110.315 69.640 113.895 ;
        RECT 69.405 105.235 69.640 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 116.210 69.730 153.550 ;
        RECT 69.300 116.345 69.865 153.425 ;
        RECT 69.300 116.340 69.860 153.430 ;
        RECT 69.300 116.330 69.850 153.440 ;
        RECT 69.300 116.320 69.840 153.450 ;
        RECT 69.300 116.310 69.830 153.460 ;
        RECT 69.300 116.300 69.820 153.470 ;
        RECT 69.300 116.290 69.810 153.480 ;
        RECT 69.300 116.280 69.800 153.490 ;
        RECT 69.300 116.270 69.790 153.500 ;
        RECT 69.300 116.260 69.780 153.510 ;
        RECT 69.300 116.250 69.770 153.520 ;
        RECT 69.300 116.240 69.760 153.530 ;
        RECT 69.300 116.230 69.750 153.540 ;
        RECT 69.300 116.220 69.740 153.550 ;
  END 
END PLBI16N

MACRO PLBI16F
  CLASS  PAD ;
  FOREIGN PLBI16F 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V6 ;
        RECT 9.520 173.510 9.880 173.870 ;
      LAYER M4 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V3 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M3 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V2 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M2 ;
        RECT 9.600 173.300 9.800 174.000 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V1 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M1 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER M6 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V5 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M5 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V4 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V6 ;
        RECT 66.240 173.510 66.600 173.870 ;
      LAYER M4 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V3 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M3 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V2 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M2 ;
        RECT 66.320 173.300 66.520 174.000 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V1 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M1 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER M6 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V5 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M5 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V4 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V6 ;
        RECT 21.400 173.510 21.760 173.870 ;
      LAYER M4 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V3 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M3 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V2 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M2 ;
        RECT 21.480 173.300 21.680 174.000 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V1 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M1 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER M6 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V5 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M5 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V4 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V6 ;
        RECT 28.545 173.510 28.905 173.870 ;
      LAYER M4 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V3 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M3 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V2 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M2 ;
        RECT 28.625 173.300 28.825 174.000 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V1 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M1 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER M6 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V5 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M5 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V4 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V6 ;
        RECT 24.395 173.510 24.755 173.870 ;
      LAYER M4 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V3 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M3 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V2 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M2 ;
        RECT 24.475 173.300 24.675 174.000 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V1 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M1 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER M6 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V5 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M5 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V4 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V6 ;
        RECT 17.995 173.510 18.355 173.870 ;
      LAYER M4 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V3 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M3 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V2 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M2 ;
        RECT 18.075 173.300 18.275 174.000 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V1 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M1 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER M6 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V5 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M5 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V4 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V6 ;
        RECT 13.620 173.510 13.980 173.870 ;
      LAYER M4 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V3 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M3 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V2 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M2 ;
        RECT 13.700 173.300 13.900 174.000 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V1 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M1 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER M6 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V5 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M5 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V4 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V6 ;
        RECT 51.035 173.510 51.395 173.870 ;
      LAYER M4 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V3 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M3 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V2 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M2 ;
        RECT 51.115 173.300 51.315 174.000 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V1 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M1 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER M6 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V5 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M5 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V4 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.405 110.315 69.640 113.895 ;
        RECT 69.405 105.235 69.640 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.855 ;
        RECT 69.300 152.430 70.000 152.730 ;
        RECT 69.640 115.135 70.000 154.220 ;
        RECT 69.300 153.920 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.405 110.315 69.640 113.895 ;
        RECT 69.405 105.235 69.640 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 150.095 69.870 150.295 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.415 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.405 110.315 69.640 113.895 ;
        RECT 69.405 105.235 69.640 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 116.210 69.730 153.550 ;
        RECT 69.300 116.345 69.865 153.425 ;
        RECT 69.300 116.340 69.860 153.430 ;
        RECT 69.300 116.330 69.850 153.440 ;
        RECT 69.300 116.320 69.840 153.450 ;
        RECT 69.300 116.310 69.830 153.460 ;
        RECT 69.300 116.300 69.820 153.470 ;
        RECT 69.300 116.290 69.810 153.480 ;
        RECT 69.300 116.280 69.800 153.490 ;
        RECT 69.300 116.270 69.790 153.500 ;
        RECT 69.300 116.260 69.780 153.510 ;
        RECT 69.300 116.250 69.770 153.520 ;
        RECT 69.300 116.240 69.760 153.530 ;
        RECT 69.300 116.230 69.750 153.540 ;
        RECT 69.300 116.220 69.740 153.550 ;
  END 
END PLBI16F

MACRO PLBI8S
  CLASS  PAD ;
  FOREIGN PLBI8S 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V6 ;
        RECT 9.520 173.510 9.880 173.870 ;
      LAYER M4 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V3 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M3 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V2 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M2 ;
        RECT 9.600 173.300 9.800 174.000 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V1 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M1 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER M6 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V5 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M5 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V4 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V6 ;
        RECT 66.240 173.510 66.600 173.870 ;
      LAYER M4 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V3 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M3 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V2 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M2 ;
        RECT 66.320 173.300 66.520 174.000 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V1 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M1 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER M6 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V5 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M5 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V4 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V6 ;
        RECT 21.400 173.510 21.760 173.870 ;
      LAYER M4 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V3 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M3 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V2 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M2 ;
        RECT 21.480 173.300 21.680 174.000 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V1 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M1 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER M6 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V5 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M5 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V4 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V6 ;
        RECT 28.545 173.510 28.905 173.870 ;
      LAYER M4 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V3 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M3 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V2 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M2 ;
        RECT 28.625 173.300 28.825 174.000 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V1 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M1 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER M6 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V5 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M5 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V4 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V6 ;
        RECT 24.395 173.510 24.755 173.870 ;
      LAYER M4 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V3 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M3 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V2 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M2 ;
        RECT 24.475 173.300 24.675 174.000 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V1 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M1 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER M6 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V5 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M5 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V4 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V6 ;
        RECT 17.995 173.510 18.355 173.870 ;
      LAYER M4 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V3 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M3 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V2 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M2 ;
        RECT 18.075 173.300 18.275 174.000 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V1 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M1 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER M6 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V5 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M5 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V4 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V6 ;
        RECT 13.620 173.510 13.980 173.870 ;
      LAYER M4 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V3 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M3 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V2 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M2 ;
        RECT 13.700 173.300 13.900 174.000 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V1 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M1 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER M6 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V5 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M5 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V4 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V6 ;
        RECT 51.035 173.510 51.395 173.870 ;
      LAYER M4 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V3 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M3 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V2 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M2 ;
        RECT 51.115 173.300 51.315 174.000 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V1 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M1 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER M6 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V5 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M5 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V4 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.430 110.315 69.665 113.895 ;
        RECT 69.430 105.235 69.665 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.855 ;
        RECT 69.300 152.430 70.000 152.730 ;
        RECT 69.640 115.135 70.000 154.220 ;
        RECT 69.300 153.920 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.430 110.315 69.665 113.895 ;
        RECT 69.430 105.235 69.665 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 150.095 69.870 150.295 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.415 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.430 110.315 69.665 113.895 ;
        RECT 69.430 105.235 69.665 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 116.210 69.730 153.550 ;
        RECT 69.300 116.345 69.865 153.425 ;
        RECT 69.300 116.340 69.860 153.430 ;
        RECT 69.300 116.330 69.850 153.440 ;
        RECT 69.300 116.320 69.840 153.450 ;
        RECT 69.300 116.310 69.830 153.460 ;
        RECT 69.300 116.300 69.820 153.470 ;
        RECT 69.300 116.290 69.810 153.480 ;
        RECT 69.300 116.280 69.800 153.490 ;
        RECT 69.300 116.270 69.790 153.500 ;
        RECT 69.300 116.260 69.780 153.510 ;
        RECT 69.300 116.250 69.770 153.520 ;
        RECT 69.300 116.240 69.760 153.530 ;
        RECT 69.300 116.230 69.750 153.540 ;
        RECT 69.300 116.220 69.740 153.550 ;
  END 
END PLBI8S

MACRO PLBI8N
  CLASS  PAD ;
  FOREIGN PLBI8N 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V6 ;
        RECT 9.520 173.510 9.880 173.870 ;
      LAYER M4 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V3 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M3 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V2 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M2 ;
        RECT 9.600 173.300 9.800 174.000 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V1 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M1 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER M6 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V5 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M5 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V4 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V6 ;
        RECT 66.240 173.510 66.600 173.870 ;
      LAYER M4 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V3 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M3 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V2 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M2 ;
        RECT 66.320 173.300 66.520 174.000 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V1 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M1 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER M6 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V5 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M5 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V4 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V6 ;
        RECT 21.400 173.510 21.760 173.870 ;
      LAYER M4 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V3 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M3 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V2 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M2 ;
        RECT 21.480 173.300 21.680 174.000 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V1 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M1 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER M6 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V5 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M5 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V4 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V6 ;
        RECT 28.545 173.510 28.905 173.870 ;
      LAYER M4 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V3 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M3 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V2 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M2 ;
        RECT 28.625 173.300 28.825 174.000 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V1 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M1 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER M6 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V5 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M5 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V4 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V6 ;
        RECT 24.395 173.510 24.755 173.870 ;
      LAYER M4 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V3 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M3 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V2 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M2 ;
        RECT 24.475 173.300 24.675 174.000 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V1 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M1 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER M6 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V5 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M5 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V4 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V6 ;
        RECT 17.995 173.510 18.355 173.870 ;
      LAYER M4 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V3 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M3 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V2 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M2 ;
        RECT 18.075 173.300 18.275 174.000 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V1 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M1 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER M6 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V5 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M5 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V4 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V6 ;
        RECT 13.620 173.510 13.980 173.870 ;
      LAYER M4 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V3 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M3 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V2 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M2 ;
        RECT 13.700 173.300 13.900 174.000 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V1 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M1 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER M6 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V5 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M5 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V4 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V6 ;
        RECT 51.035 173.510 51.395 173.870 ;
      LAYER M4 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V3 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M3 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V2 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M2 ;
        RECT 51.115 173.300 51.315 174.000 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V1 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M1 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER M6 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V5 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M5 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V4 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.430 110.315 69.665 113.895 ;
        RECT 69.430 105.235 69.665 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.855 ;
        RECT 69.300 152.430 70.000 152.730 ;
        RECT 69.640 115.135 70.000 154.220 ;
        RECT 69.300 153.920 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.430 110.315 69.665 113.895 ;
        RECT 69.430 105.235 69.665 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 150.095 69.870 150.295 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.415 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.430 110.315 69.665 113.895 ;
        RECT 69.430 105.235 69.665 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 116.210 69.730 153.550 ;
        RECT 69.300 116.345 69.865 153.425 ;
        RECT 69.300 116.340 69.860 153.430 ;
        RECT 69.300 116.330 69.850 153.440 ;
        RECT 69.300 116.320 69.840 153.450 ;
        RECT 69.300 116.310 69.830 153.460 ;
        RECT 69.300 116.300 69.820 153.470 ;
        RECT 69.300 116.290 69.810 153.480 ;
        RECT 69.300 116.280 69.800 153.490 ;
        RECT 69.300 116.270 69.790 153.500 ;
        RECT 69.300 116.260 69.780 153.510 ;
        RECT 69.300 116.250 69.770 153.520 ;
        RECT 69.300 116.240 69.760 153.530 ;
        RECT 69.300 116.230 69.750 153.540 ;
        RECT 69.300 116.220 69.740 153.550 ;
  END 
END PLBI8N

MACRO PLBI8F
  CLASS  PAD ;
  FOREIGN PLBI8F 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V6 ;
        RECT 9.520 173.510 9.880 173.870 ;
      LAYER M4 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V3 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M3 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V2 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M2 ;
        RECT 9.600 173.300 9.800 174.000 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V1 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M1 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER M6 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V5 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M5 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V4 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V6 ;
        RECT 66.240 173.510 66.600 173.870 ;
      LAYER M4 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V3 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M3 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V2 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M2 ;
        RECT 66.320 173.300 66.520 174.000 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V1 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M1 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER M6 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V5 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M5 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V4 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V6 ;
        RECT 21.400 173.510 21.760 173.870 ;
      LAYER M4 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V3 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M3 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V2 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M2 ;
        RECT 21.480 173.300 21.680 174.000 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V1 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M1 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER M6 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V5 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M5 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V4 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V6 ;
        RECT 28.545 173.510 28.905 173.870 ;
      LAYER M4 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V3 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M3 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V2 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M2 ;
        RECT 28.625 173.300 28.825 174.000 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V1 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M1 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER M6 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V5 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M5 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V4 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V6 ;
        RECT 24.395 173.510 24.755 173.870 ;
      LAYER M4 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V3 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M3 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V2 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M2 ;
        RECT 24.475 173.300 24.675 174.000 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V1 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M1 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER M6 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V5 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M5 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V4 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V6 ;
        RECT 17.995 173.510 18.355 173.870 ;
      LAYER M4 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V3 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M3 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V2 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M2 ;
        RECT 18.075 173.300 18.275 174.000 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V1 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M1 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER M6 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V5 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M5 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V4 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V6 ;
        RECT 13.620 173.510 13.980 173.870 ;
      LAYER M4 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V3 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M3 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V2 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M2 ;
        RECT 13.700 173.300 13.900 174.000 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V1 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M1 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER M6 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V5 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M5 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V4 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V6 ;
        RECT 51.035 173.510 51.395 173.870 ;
      LAYER M4 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V3 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M3 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V2 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M2 ;
        RECT 51.115 173.300 51.315 174.000 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V1 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M1 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER M6 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V5 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M5 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V4 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.430 110.315 69.665 113.895 ;
        RECT 69.430 105.235 69.665 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.855 ;
        RECT 69.300 152.430 70.000 152.730 ;
        RECT 69.640 115.135 70.000 154.220 ;
        RECT 69.300 153.920 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.430 110.315 69.665 113.895 ;
        RECT 69.430 105.235 69.665 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 150.095 69.870 150.295 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.415 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.430 110.315 69.665 113.895 ;
        RECT 69.430 105.235 69.665 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 116.210 69.730 153.550 ;
        RECT 69.300 116.345 69.865 153.425 ;
        RECT 69.300 116.340 69.860 153.430 ;
        RECT 69.300 116.330 69.850 153.440 ;
        RECT 69.300 116.320 69.840 153.450 ;
        RECT 69.300 116.310 69.830 153.460 ;
        RECT 69.300 116.300 69.820 153.470 ;
        RECT 69.300 116.290 69.810 153.480 ;
        RECT 69.300 116.280 69.800 153.490 ;
        RECT 69.300 116.270 69.790 153.500 ;
        RECT 69.300 116.260 69.780 153.510 ;
        RECT 69.300 116.250 69.770 153.520 ;
        RECT 69.300 116.240 69.760 153.530 ;
        RECT 69.300 116.230 69.750 153.540 ;
        RECT 69.300 116.220 69.740 153.550 ;
  END 
END PLBI8F

MACRO PLBI4S
  CLASS  PAD ;
  FOREIGN PLBI4S 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V6 ;
        RECT 9.520 173.510 9.880 173.870 ;
      LAYER M4 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V3 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M3 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V2 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M2 ;
        RECT 9.600 173.300 9.800 174.000 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V1 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M1 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER M6 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V5 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M5 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V4 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V6 ;
        RECT 66.240 173.510 66.600 173.870 ;
      LAYER M4 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V3 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M3 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V2 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M2 ;
        RECT 66.320 173.300 66.520 174.000 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V1 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M1 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER M6 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V5 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M5 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V4 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V6 ;
        RECT 21.400 173.510 21.760 173.870 ;
      LAYER M4 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V3 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M3 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V2 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M2 ;
        RECT 21.480 173.300 21.680 174.000 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V1 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M1 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER M6 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V5 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M5 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V4 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V6 ;
        RECT 28.545 173.510 28.905 173.870 ;
      LAYER M4 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V3 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M3 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V2 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M2 ;
        RECT 28.625 173.300 28.825 174.000 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V1 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M1 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER M6 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V5 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M5 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V4 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V6 ;
        RECT 24.395 173.510 24.755 173.870 ;
      LAYER M4 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V3 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M3 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V2 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M2 ;
        RECT 24.475 173.300 24.675 174.000 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V1 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M1 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER M6 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V5 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M5 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V4 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V6 ;
        RECT 17.995 173.510 18.355 173.870 ;
      LAYER M4 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V3 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M3 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V2 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M2 ;
        RECT 18.075 173.300 18.275 174.000 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V1 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M1 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER M6 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V5 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M5 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V4 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V6 ;
        RECT 13.620 173.510 13.980 173.870 ;
      LAYER M4 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V3 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M3 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V2 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M2 ;
        RECT 13.700 173.300 13.900 174.000 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V1 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M1 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER M6 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V5 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M5 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V4 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V6 ;
        RECT 51.035 173.510 51.395 173.870 ;
      LAYER M4 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V3 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M3 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V2 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M2 ;
        RECT 51.115 173.300 51.315 174.000 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V1 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M1 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER M6 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V5 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M5 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V4 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.415 110.315 69.680 113.895 ;
        RECT 69.415 105.235 69.680 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.855 ;
        RECT 69.300 152.430 70.000 152.730 ;
        RECT 69.640 115.135 70.000 154.220 ;
        RECT 69.300 153.920 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.415 110.315 69.680 113.895 ;
        RECT 69.415 105.235 69.680 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 150.095 69.870 150.295 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.415 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.415 110.315 69.680 113.895 ;
        RECT 69.415 105.235 69.680 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 116.210 69.730 153.550 ;
        RECT 69.300 116.345 69.865 153.425 ;
        RECT 69.300 116.340 69.860 153.430 ;
        RECT 69.300 116.330 69.850 153.440 ;
        RECT 69.300 116.320 69.840 153.450 ;
        RECT 69.300 116.310 69.830 153.460 ;
        RECT 69.300 116.300 69.820 153.470 ;
        RECT 69.300 116.290 69.810 153.480 ;
        RECT 69.300 116.280 69.800 153.490 ;
        RECT 69.300 116.270 69.790 153.500 ;
        RECT 69.300 116.260 69.780 153.510 ;
        RECT 69.300 116.250 69.770 153.520 ;
        RECT 69.300 116.240 69.760 153.530 ;
        RECT 69.300 116.230 69.750 153.540 ;
        RECT 69.300 116.220 69.740 153.550 ;
  END 
END PLBI4S

MACRO PLBI4N
  CLASS  PAD ;
  FOREIGN PLBI4N 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V6 ;
        RECT 9.520 173.510 9.880 173.870 ;
      LAYER M4 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V3 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M3 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V2 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M2 ;
        RECT 9.600 173.300 9.800 174.000 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V1 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M1 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER M6 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V5 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M5 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V4 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V6 ;
        RECT 66.240 173.510 66.600 173.870 ;
      LAYER M4 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V3 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M3 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V2 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M2 ;
        RECT 66.320 173.300 66.520 174.000 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V1 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M1 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER M6 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V5 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M5 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V4 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V6 ;
        RECT 21.400 173.510 21.760 173.870 ;
      LAYER M4 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V3 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M3 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V2 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M2 ;
        RECT 21.480 173.300 21.680 174.000 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V1 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M1 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER M6 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V5 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M5 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V4 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V6 ;
        RECT 28.545 173.510 28.905 173.870 ;
      LAYER M4 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V3 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M3 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V2 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M2 ;
        RECT 28.625 173.300 28.825 174.000 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V1 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M1 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER M6 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V5 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M5 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V4 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V6 ;
        RECT 24.395 173.510 24.755 173.870 ;
      LAYER M4 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V3 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M3 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V2 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M2 ;
        RECT 24.475 173.300 24.675 174.000 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V1 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M1 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER M6 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V5 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M5 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V4 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V6 ;
        RECT 17.995 173.510 18.355 173.870 ;
      LAYER M4 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V3 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M3 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V2 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M2 ;
        RECT 18.075 173.300 18.275 174.000 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V1 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M1 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER M6 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V5 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M5 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V4 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V6 ;
        RECT 13.620 173.510 13.980 173.870 ;
      LAYER M4 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V3 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M3 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V2 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M2 ;
        RECT 13.700 173.300 13.900 174.000 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V1 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M1 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER M6 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V5 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M5 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V4 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V6 ;
        RECT 51.035 173.510 51.395 173.870 ;
      LAYER M4 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V3 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M3 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V2 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M2 ;
        RECT 51.115 173.300 51.315 174.000 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V1 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M1 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER M6 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V5 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M5 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V4 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.415 110.315 69.680 113.895 ;
        RECT 69.415 105.235 69.680 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.855 ;
        RECT 69.300 152.430 70.000 152.730 ;
        RECT 69.640 115.135 70.000 154.220 ;
        RECT 69.300 153.920 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.415 110.315 69.680 113.895 ;
        RECT 69.415 105.235 69.680 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 150.095 69.870 150.295 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.415 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.415 110.315 69.680 113.895 ;
        RECT 69.415 105.235 69.680 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 116.210 69.730 153.550 ;
        RECT 69.300 116.345 69.865 153.425 ;
        RECT 69.300 116.340 69.860 153.430 ;
        RECT 69.300 116.330 69.850 153.440 ;
        RECT 69.300 116.320 69.840 153.450 ;
        RECT 69.300 116.310 69.830 153.460 ;
        RECT 69.300 116.300 69.820 153.470 ;
        RECT 69.300 116.290 69.810 153.480 ;
        RECT 69.300 116.280 69.800 153.490 ;
        RECT 69.300 116.270 69.790 153.500 ;
        RECT 69.300 116.260 69.780 153.510 ;
        RECT 69.300 116.250 69.770 153.520 ;
        RECT 69.300 116.240 69.760 153.530 ;
        RECT 69.300 116.230 69.750 153.540 ;
        RECT 69.300 116.220 69.740 153.550 ;
  END 
END PLBI4N

MACRO PLBI4F
  CLASS  PAD ;
  FOREIGN PLBI4F 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V6 ;
        RECT 9.520 173.510 9.880 173.870 ;
      LAYER M4 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V3 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M3 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V2 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M2 ;
        RECT 9.600 173.300 9.800 174.000 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V1 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M1 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER M6 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V5 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M5 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V4 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V6 ;
        RECT 66.240 173.510 66.600 173.870 ;
      LAYER M4 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V3 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M3 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V2 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M2 ;
        RECT 66.320 173.300 66.520 174.000 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V1 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M1 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER M6 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V5 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M5 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V4 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V6 ;
        RECT 21.400 173.510 21.760 173.870 ;
      LAYER M4 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V3 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M3 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V2 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M2 ;
        RECT 21.480 173.300 21.680 174.000 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V1 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M1 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER M6 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V5 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M5 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V4 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V6 ;
        RECT 28.545 173.510 28.905 173.870 ;
      LAYER M4 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V3 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M3 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V2 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M2 ;
        RECT 28.625 173.300 28.825 174.000 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V1 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M1 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER M6 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V5 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M5 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V4 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V6 ;
        RECT 24.395 173.510 24.755 173.870 ;
      LAYER M4 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V3 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M3 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V2 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M2 ;
        RECT 24.475 173.300 24.675 174.000 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V1 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M1 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER M6 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V5 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M5 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V4 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V6 ;
        RECT 17.995 173.510 18.355 173.870 ;
      LAYER M4 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V3 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M3 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V2 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M2 ;
        RECT 18.075 173.300 18.275 174.000 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V1 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M1 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER M6 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V5 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M5 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V4 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V6 ;
        RECT 13.620 173.510 13.980 173.870 ;
      LAYER M4 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V3 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M3 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V2 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M2 ;
        RECT 13.700 173.300 13.900 174.000 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V1 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M1 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER M6 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V5 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M5 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V4 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V6 ;
        RECT 51.035 173.510 51.395 173.870 ;
      LAYER M4 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V3 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M3 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V2 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M2 ;
        RECT 51.115 173.300 51.315 174.000 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V1 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M1 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER M6 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V5 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M5 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V4 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.415 110.315 69.680 113.895 ;
        RECT 69.415 105.235 69.680 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.855 ;
        RECT 69.300 152.430 70.000 152.730 ;
        RECT 69.640 115.135 70.000 154.220 ;
        RECT 69.300 153.920 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.415 110.315 69.680 113.895 ;
        RECT 69.415 105.235 69.680 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 150.095 69.870 150.295 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.415 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.415 110.315 69.680 113.895 ;
        RECT 69.415 105.235 69.680 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 116.210 69.730 153.550 ;
        RECT 69.300 116.345 69.865 153.425 ;
        RECT 69.300 116.340 69.860 153.430 ;
        RECT 69.300 116.330 69.850 153.440 ;
        RECT 69.300 116.320 69.840 153.450 ;
        RECT 69.300 116.310 69.830 153.460 ;
        RECT 69.300 116.300 69.820 153.470 ;
        RECT 69.300 116.290 69.810 153.480 ;
        RECT 69.300 116.280 69.800 153.490 ;
        RECT 69.300 116.270 69.790 153.500 ;
        RECT 69.300 116.260 69.780 153.510 ;
        RECT 69.300 116.250 69.770 153.520 ;
        RECT 69.300 116.240 69.760 153.530 ;
        RECT 69.300 116.230 69.750 153.540 ;
        RECT 69.300 116.220 69.740 153.550 ;
  END 
END PLBI4F

MACRO PLBI2S
  CLASS  PAD ;
  FOREIGN PLBI2S 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V6 ;
        RECT 9.520 173.510 9.880 173.870 ;
      LAYER M4 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V3 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M3 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V2 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M2 ;
        RECT 9.600 173.300 9.800 174.000 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V1 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M1 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER M6 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V5 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M5 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V4 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V6 ;
        RECT 66.240 173.510 66.600 173.870 ;
      LAYER M4 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V3 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M3 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V2 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M2 ;
        RECT 66.320 173.300 66.520 174.000 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V1 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M1 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER M6 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V5 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M5 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V4 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V6 ;
        RECT 21.400 173.510 21.760 173.870 ;
      LAYER M4 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V3 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M3 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V2 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M2 ;
        RECT 21.480 173.300 21.680 174.000 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V1 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M1 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER M6 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V5 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M5 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V4 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V6 ;
        RECT 28.545 173.510 28.905 173.870 ;
      LAYER M4 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V3 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M3 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V2 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M2 ;
        RECT 28.625 173.300 28.825 174.000 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V1 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M1 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER M6 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V5 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M5 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V4 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V6 ;
        RECT 24.395 173.510 24.755 173.870 ;
      LAYER M4 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V3 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M3 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V2 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M2 ;
        RECT 24.475 173.300 24.675 174.000 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V1 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M1 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER M6 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V5 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M5 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V4 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V6 ;
        RECT 17.995 173.510 18.355 173.870 ;
      LAYER M4 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V3 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M3 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V2 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M2 ;
        RECT 18.075 173.300 18.275 174.000 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V1 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M1 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER M6 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V5 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M5 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V4 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V6 ;
        RECT 13.620 173.510 13.980 173.870 ;
      LAYER M4 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V3 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M3 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V2 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M2 ;
        RECT 13.700 173.300 13.900 174.000 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V1 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M1 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER M6 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V5 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M5 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V4 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V6 ;
        RECT 51.035 173.510 51.395 173.870 ;
      LAYER M4 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V3 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M3 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V2 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M2 ;
        RECT 51.115 173.300 51.315 174.000 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V1 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M1 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER M6 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V5 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M5 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V4 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.430 110.315 69.630 113.895 ;
        RECT 69.430 105.215 69.630 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.855 ;
        RECT 69.300 152.430 70.000 152.730 ;
        RECT 69.640 115.135 70.000 154.220 ;
        RECT 69.300 153.920 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.430 110.315 69.630 113.895 ;
        RECT 69.430 105.215 69.630 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 150.095 69.870 150.295 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.415 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.430 110.315 69.630 113.895 ;
        RECT 69.430 105.215 69.630 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 116.210 69.730 153.550 ;
        RECT 69.300 116.345 69.865 153.425 ;
        RECT 69.300 116.340 69.860 153.430 ;
        RECT 69.300 116.330 69.850 153.440 ;
        RECT 69.300 116.320 69.840 153.450 ;
        RECT 69.300 116.310 69.830 153.460 ;
        RECT 69.300 116.300 69.820 153.470 ;
        RECT 69.300 116.290 69.810 153.480 ;
        RECT 69.300 116.280 69.800 153.490 ;
        RECT 69.300 116.270 69.790 153.500 ;
        RECT 69.300 116.260 69.780 153.510 ;
        RECT 69.300 116.250 69.770 153.520 ;
        RECT 69.300 116.240 69.760 153.530 ;
        RECT 69.300 116.230 69.750 153.540 ;
        RECT 69.300 116.220 69.740 153.550 ;
  END 
END PLBI2S

MACRO PLBI2N
  CLASS  PAD ;
  FOREIGN PLBI2N 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V6 ;
        RECT 9.520 173.510 9.880 173.870 ;
      LAYER M4 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V3 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M3 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V2 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M2 ;
        RECT 9.600 173.300 9.800 174.000 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V1 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M1 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER M6 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V5 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M5 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V4 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V6 ;
        RECT 66.240 173.510 66.600 173.870 ;
      LAYER M4 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V3 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M3 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V2 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M2 ;
        RECT 66.320 173.300 66.520 174.000 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V1 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M1 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER M6 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V5 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M5 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V4 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V6 ;
        RECT 21.400 173.510 21.760 173.870 ;
      LAYER M4 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V3 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M3 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V2 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M2 ;
        RECT 21.480 173.300 21.680 174.000 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V1 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M1 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER M6 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V5 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M5 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V4 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V6 ;
        RECT 28.545 173.510 28.905 173.870 ;
      LAYER M4 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V3 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M3 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V2 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M2 ;
        RECT 28.625 173.300 28.825 174.000 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V1 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M1 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER M6 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V5 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M5 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V4 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V6 ;
        RECT 24.395 173.510 24.755 173.870 ;
      LAYER M4 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V3 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M3 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V2 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M2 ;
        RECT 24.475 173.300 24.675 174.000 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V1 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M1 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER M6 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V5 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M5 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V4 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V6 ;
        RECT 17.995 173.510 18.355 173.870 ;
      LAYER M4 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V3 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M3 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V2 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M2 ;
        RECT 18.075 173.300 18.275 174.000 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V1 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M1 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER M6 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V5 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M5 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V4 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V6 ;
        RECT 13.620 173.510 13.980 173.870 ;
      LAYER M4 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V3 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M3 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V2 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M2 ;
        RECT 13.700 173.300 13.900 174.000 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V1 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M1 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER M6 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V5 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M5 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V4 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V6 ;
        RECT 51.035 173.510 51.395 173.870 ;
      LAYER M4 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V3 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M3 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V2 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M2 ;
        RECT 51.115 173.300 51.315 174.000 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V1 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M1 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER M6 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V5 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M5 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V4 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.430 110.315 69.630 113.895 ;
        RECT 69.430 105.215 69.630 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.855 ;
        RECT 69.300 152.430 70.000 152.730 ;
        RECT 69.640 115.135 70.000 154.220 ;
        RECT 69.300 153.920 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.430 110.315 69.630 113.895 ;
        RECT 69.430 105.215 69.630 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 150.095 69.870 150.295 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.415 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.430 110.315 69.630 113.895 ;
        RECT 69.430 105.215 69.630 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 116.210 69.730 153.550 ;
        RECT 69.300 116.345 69.865 153.425 ;
        RECT 69.300 116.340 69.860 153.430 ;
        RECT 69.300 116.330 69.850 153.440 ;
        RECT 69.300 116.320 69.840 153.450 ;
        RECT 69.300 116.310 69.830 153.460 ;
        RECT 69.300 116.300 69.820 153.470 ;
        RECT 69.300 116.290 69.810 153.480 ;
        RECT 69.300 116.280 69.800 153.490 ;
        RECT 69.300 116.270 69.790 153.500 ;
        RECT 69.300 116.260 69.780 153.510 ;
        RECT 69.300 116.250 69.770 153.520 ;
        RECT 69.300 116.240 69.760 153.530 ;
        RECT 69.300 116.230 69.750 153.540 ;
        RECT 69.300 116.220 69.740 153.550 ;
  END 
END PLBI2N

MACRO PLBI2F
  CLASS  PAD ;
  FOREIGN PLBI2F 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 174.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M7 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M4 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M3 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M2 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M6 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
      LAYER M5 ;
        RECT 3.000 0.665 67.000 0.700 ;
        RECT 3.010 0.660 66.995 0.700 ;
        RECT 3.010 0.655 66.985 0.700 ;
        RECT 3.020 0.650 66.985 0.700 ;
        RECT 3.020 0.645 66.975 0.700 ;
        RECT 3.030 0.640 66.975 0.700 ;
        RECT 3.030 0.635 66.965 0.700 ;
        RECT 3.040 0.630 66.965 0.700 ;
        RECT 3.040 0.625 66.955 0.700 ;
        RECT 3.050 0.620 66.955 0.700 ;
        RECT 3.050 0.615 66.945 0.700 ;
        RECT 3.060 0.610 66.945 0.700 ;
        RECT 3.060 0.605 66.935 0.700 ;
        RECT 3.070 0.600 66.935 0.700 ;
        RECT 3.070 0.595 66.925 0.700 ;
        RECT 3.080 0.590 66.925 0.700 ;
        RECT 3.080 0.585 66.915 0.700 ;
        RECT 3.090 0.580 66.915 0.700 ;
        RECT 3.090 0.575 66.905 0.700 ;
        RECT 3.100 0.570 66.905 0.700 ;
        RECT 3.100 0.565 66.895 0.700 ;
        RECT 3.110 0.560 66.895 0.700 ;
        RECT 3.110 0.555 66.885 0.700 ;
        RECT 3.120 0.550 66.885 0.700 ;
        RECT 3.120 0.545 66.875 0.700 ;
        RECT 3.130 0.540 66.875 0.700 ;
        RECT 3.130 0.535 66.865 0.700 ;
        RECT 3.140 0.530 66.865 0.700 ;
        RECT 3.140 0.525 66.855 0.700 ;
        RECT 3.150 0.520 66.855 0.700 ;
        RECT 3.150 0.515 66.845 0.700 ;
        RECT 3.160 0.510 66.845 0.700 ;
        RECT 3.160 0.505 66.835 0.700 ;
        RECT 3.170 0.500 66.835 0.700 ;
        RECT 3.170 0.495 66.825 0.700 ;
        RECT 3.180 0.490 66.825 0.700 ;
        RECT 3.180 0.485 66.815 0.700 ;
        RECT 3.190 0.480 66.815 0.700 ;
        RECT 3.190 0.475 66.805 0.700 ;
        RECT 3.200 0.470 66.805 0.700 ;
        RECT 3.200 0.465 66.795 0.700 ;
        RECT 3.210 0.460 66.795 0.700 ;
        RECT 3.210 0.455 66.785 0.700 ;
        RECT 3.220 0.450 66.785 0.700 ;
        RECT 3.220 0.445 66.775 0.700 ;
        RECT 3.230 0.440 66.775 0.700 ;
        RECT 3.230 0.435 66.765 0.700 ;
        RECT 3.240 0.430 66.765 0.700 ;
        RECT 3.240 0.425 66.755 0.700 ;
        RECT 3.250 0.420 66.755 0.700 ;
        RECT 3.250 0.415 66.745 0.700 ;
        RECT 3.260 0.410 66.745 0.700 ;
        RECT 3.260 0.405 66.735 0.700 ;
        RECT 3.270 0.400 66.735 0.700 ;
        RECT 3.270 0.395 66.725 0.700 ;
        RECT 3.280 0.390 66.725 0.700 ;
        RECT 3.280 0.385 66.715 0.700 ;
        RECT 3.290 0.380 66.715 0.700 ;
        RECT 3.290 0.375 66.705 0.700 ;
        RECT 3.300 0.370 66.705 0.700 ;
        RECT 3.300 0.365 66.695 0.700 ;
        RECT 3.310 0.360 66.695 0.700 ;
        RECT 3.310 0.355 66.685 0.700 ;
        RECT 3.320 0.350 66.685 0.700 ;
        RECT 3.320 0.345 66.675 0.700 ;
        RECT 3.330 0.340 66.675 0.700 ;
        RECT 3.330 0.335 66.665 0.700 ;
        RECT 3.340 0.330 66.665 0.700 ;
        RECT 3.340 0.325 66.655 0.700 ;
        RECT 3.350 0.320 66.655 0.700 ;
        RECT 3.350 0.315 66.645 0.700 ;
        RECT 3.360 0.310 66.645 0.700 ;
        RECT 3.360 0.305 66.635 0.700 ;
        RECT 3.370 0.300 66.635 0.700 ;
        RECT 3.370 0.295 66.625 0.700 ;
        RECT 3.380 0.290 66.625 0.700 ;
        RECT 3.380 0.285 66.615 0.700 ;
        RECT 3.390 0.280 66.615 0.700 ;
        RECT 3.390 0.275 66.605 0.700 ;
        RECT 3.400 0.270 66.605 0.700 ;
        RECT 3.400 0.265 66.595 0.700 ;
        RECT 3.410 0.260 66.595 0.700 ;
        RECT 3.410 0.255 66.585 0.700 ;
        RECT 3.420 0.250 66.585 0.700 ;
        RECT 3.420 0.245 66.575 0.700 ;
        RECT 3.430 0.240 66.575 0.700 ;
        RECT 3.430 0.235 66.565 0.700 ;
        RECT 3.440 0.230 66.565 0.700 ;
        RECT 3.440 0.225 66.555 0.700 ;
        RECT 3.450 0.220 66.555 0.700 ;
        RECT 3.450 0.215 66.545 0.700 ;
        RECT 3.460 0.210 66.545 0.700 ;
        RECT 3.460 0.205 66.535 0.700 ;
        RECT 3.470 0.200 66.535 0.700 ;
        RECT 3.470 0.195 66.525 0.700 ;
        RECT 3.480 0.190 66.525 0.700 ;
        RECT 3.480 0.185 66.515 0.700 ;
        RECT 3.490 0.180 66.515 0.700 ;
        RECT 3.490 0.175 66.505 0.700 ;
        RECT 3.500 0.170 66.505 0.700 ;
        RECT 3.500 0.165 66.495 0.700 ;
        RECT 3.510 0.160 66.495 0.700 ;
        RECT 3.510 0.155 66.485 0.700 ;
        RECT 3.520 0.150 66.485 0.700 ;
        RECT 3.520 0.145 66.475 0.700 ;
        RECT 3.530 0.140 66.475 0.700 ;
        RECT 3.530 0.135 66.465 0.700 ;
        RECT 3.540 0.130 66.465 0.700 ;
        RECT 3.540 0.125 66.455 0.700 ;
        RECT 3.550 0.120 66.455 0.700 ;
        RECT 3.550 0.115 66.445 0.700 ;
        RECT 3.560 0.110 66.445 0.700 ;
        RECT 3.560 0.105 66.435 0.700 ;
        RECT 3.570 0.100 66.435 0.700 ;
        RECT 3.570 0.095 66.425 0.700 ;
        RECT 3.580 0.090 66.425 0.700 ;
        RECT 3.580 0.085 66.415 0.700 ;
        RECT 3.590 0.080 66.415 0.700 ;
        RECT 3.590 0.075 66.405 0.700 ;
        RECT 3.600 0.070 66.405 0.700 ;
        RECT 3.600 0.065 66.395 0.700 ;
        RECT 3.610 0.060 66.395 0.700 ;
        RECT 3.610 0.055 66.385 0.700 ;
        RECT 3.620 0.050 66.385 0.700 ;
        RECT 3.620 0.045 66.375 0.700 ;
        RECT 3.630 0.040 66.375 0.700 ;
        RECT 3.630 0.035 66.365 0.700 ;
        RECT 3.640 0.030 66.365 0.700 ;
        RECT 3.640 0.025 66.355 0.700 ;
        RECT 3.650 0.020 66.355 0.700 ;
        RECT 3.650 0.015 66.345 0.700 ;
        RECT 3.660 0.010 66.345 0.700 ;
        RECT 3.660 0.005 66.335 0.700 ;
        RECT 3.665 0.000 66.335 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V6 ;
        RECT 9.520 173.510 9.880 173.870 ;
      LAYER M4 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V3 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M3 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V2 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M2 ;
        RECT 9.600 173.300 9.800 174.000 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V1 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M1 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER M6 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V5 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
      LAYER M5 ;
        RECT 9.200 173.380 10.200 174.000 ;
      LAYER V4 ;
        RECT 9.400 173.800 9.590 173.990 ;
        RECT 9.400 173.390 9.590 173.580 ;
        RECT 9.810 173.800 10.000 173.990 ;
        RECT 9.810 173.390 10.000 173.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M7 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V6 ;
        RECT 66.240 173.510 66.600 173.870 ;
      LAYER M4 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V3 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M3 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V2 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M2 ;
        RECT 66.320 173.300 66.520 174.000 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V1 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M1 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER M6 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V5 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
      LAYER M5 ;
        RECT 65.920 173.380 66.920 174.000 ;
      LAYER V4 ;
        RECT 66.120 173.800 66.310 173.990 ;
        RECT 66.120 173.390 66.310 173.580 ;
        RECT 66.530 173.800 66.720 173.990 ;
        RECT 66.530 173.390 66.720 173.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V6 ;
        RECT 21.400 173.510 21.760 173.870 ;
      LAYER M4 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V3 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M3 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V2 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M2 ;
        RECT 21.480 173.300 21.680 174.000 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V1 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M1 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER M6 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V5 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
      LAYER M5 ;
        RECT 21.080 173.380 22.080 174.000 ;
      LAYER V4 ;
        RECT 21.280 173.800 21.470 173.990 ;
        RECT 21.280 173.390 21.470 173.580 ;
        RECT 21.690 173.800 21.880 173.990 ;
        RECT 21.690 173.390 21.880 173.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V6 ;
        RECT 28.545 173.510 28.905 173.870 ;
      LAYER M4 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V3 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M3 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V2 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M2 ;
        RECT 28.625 173.300 28.825 174.000 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V1 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M1 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER M6 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V5 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
      LAYER M5 ;
        RECT 28.225 173.380 29.225 174.000 ;
      LAYER V4 ;
        RECT 28.425 173.800 28.615 173.990 ;
        RECT 28.425 173.390 28.615 173.580 ;
        RECT 28.835 173.800 29.025 173.990 ;
        RECT 28.835 173.390 29.025 173.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V6 ;
        RECT 24.395 173.510 24.755 173.870 ;
      LAYER M4 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V3 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M3 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V2 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M2 ;
        RECT 24.475 173.300 24.675 174.000 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V1 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M1 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER M6 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V5 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
      LAYER M5 ;
        RECT 24.075 173.380 25.075 174.000 ;
      LAYER V4 ;
        RECT 24.275 173.800 24.465 173.990 ;
        RECT 24.275 173.390 24.465 173.580 ;
        RECT 24.685 173.800 24.875 173.990 ;
        RECT 24.685 173.390 24.875 173.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V6 ;
        RECT 17.995 173.510 18.355 173.870 ;
      LAYER M4 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V3 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M3 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V2 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M2 ;
        RECT 18.075 173.300 18.275 174.000 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V1 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M1 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER M6 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V5 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
      LAYER M5 ;
        RECT 17.675 173.380 18.675 174.000 ;
      LAYER V4 ;
        RECT 17.875 173.800 18.065 173.990 ;
        RECT 17.875 173.390 18.065 173.580 ;
        RECT 18.285 173.800 18.475 173.990 ;
        RECT 18.285 173.390 18.475 173.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V6 ;
        RECT 13.620 173.510 13.980 173.870 ;
      LAYER M4 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V3 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M3 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V2 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M2 ;
        RECT 13.700 173.300 13.900 174.000 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V1 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M1 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER M6 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V5 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
      LAYER M5 ;
        RECT 13.300 173.380 14.300 174.000 ;
      LAYER V4 ;
        RECT 13.500 173.800 13.690 173.990 ;
        RECT 13.500 173.390 13.690 173.580 ;
        RECT 13.910 173.800 14.100 173.990 ;
        RECT 13.910 173.390 14.100 173.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M7 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V6 ;
        RECT 51.035 173.510 51.395 173.870 ;
      LAYER M4 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V3 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M3 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V2 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M2 ;
        RECT 51.115 173.300 51.315 174.000 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V1 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M1 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER M6 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V5 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
      LAYER M5 ;
        RECT 50.715 173.380 51.715 174.000 ;
      LAYER V4 ;
        RECT 50.915 173.800 51.105 173.990 ;
        RECT 50.915 173.390 51.105 173.580 ;
        RECT 51.325 173.800 51.515 173.990 ;
        RECT 51.325 173.390 51.515 173.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.430 110.315 69.630 113.895 ;
        RECT 69.430 105.215 69.630 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
      LAYER M1 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 115.135 0.700 154.220 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 70.000 0.700 108.815 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 115.135 70.000 115.855 ;
        RECT 69.300 152.430 70.000 152.730 ;
        RECT 69.640 115.135 70.000 154.220 ;
        RECT 69.300 153.920 70.000 154.220 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 70.000 70.000 108.815 ;
      LAYER M3 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.280 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.430 110.315 69.630 113.895 ;
        RECT 69.430 105.215 69.630 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 150.095 69.870 150.295 ;
      LAYER M6 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 137.395 0.700 147.565 ;
        RECT 0.000 127.100 0.700 134.395 ;
        RECT 0.000 121.860 0.700 124.100 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 97.700 0.700 108.815 ;
        RECT 0.000 86.640 0.700 94.700 ;
        RECT 0.000 75.630 0.700 83.640 ;
        RECT 0.000 70.000 0.700 72.630 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 137.395 70.000 147.565 ;
        RECT 69.300 127.100 70.000 134.395 ;
        RECT 69.300 121.860 70.000 124.100 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 97.700 70.000 108.815 ;
        RECT 69.300 86.640 70.000 94.700 ;
        RECT 69.300 75.630 70.000 83.640 ;
        RECT 69.300 70.000 70.000 72.630 ;
      LAYER M5 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M7 ;
        RECT 0.000 171.175 0.700 172.780 ;
        RECT 0.000 162.720 0.700 170.715 ;
        RECT 0.000 155.725 0.700 161.220 ;
        RECT 0.000 150.480 0.700 154.220 ;
        RECT 0.000 143.340 0.700 147.565 ;
        RECT 0.000 131.850 0.700 140.340 ;
        RECT 0.000 121.860 0.700 128.850 ;
        RECT 0.000 115.135 0.700 119.705 ;
        RECT 0.000 110.315 0.700 113.895 ;
        RECT 0.000 103.280 0.700 108.815 ;
        RECT 0.000 92.280 0.700 100.280 ;
        RECT 0.000 81.280 0.700 89.280 ;
        RECT 0.000 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.300 171.175 70.000 172.780 ;
        RECT 69.300 162.720 70.000 170.715 ;
        RECT 69.300 155.725 70.000 161.220 ;
        RECT 69.300 150.480 70.000 154.220 ;
        RECT 69.300 143.340 70.000 147.565 ;
        RECT 69.300 131.850 70.000 140.340 ;
        RECT 69.300 121.860 70.000 128.850 ;
        RECT 69.300 115.135 70.000 119.705 ;
        RECT 69.300 110.315 70.000 113.895 ;
        RECT 69.300 103.280 70.000 108.815 ;
        RECT 69.300 92.280 70.000 100.280 ;
        RECT 69.300 81.280 70.000 89.280 ;
        RECT 69.300 70.000 70.000 78.280 ;
      LAYER M2 ;
        RECT 0.160 171.175 0.700 172.780 ;
        RECT 0.160 162.720 0.700 170.465 ;
        RECT 0.160 155.725 0.700 161.220 ;
        RECT 0.160 150.720 0.700 154.220 ;
        RECT 0.160 115.135 0.700 119.705 ;
        RECT 0.160 110.315 0.700 113.895 ;
        RECT 0.160 105.215 0.700 108.815 ;
        RECT 0.160 92.280 0.700 100.415 ;
        RECT 0.160 81.280 0.700 89.280 ;
        RECT 0.160 70.000 0.700 78.280 ;
        RECT 1.100 1.100 68.900 172.900 ;
        RECT 69.430 110.315 69.630 113.895 ;
        RECT 69.430 105.215 69.630 108.815 ;
        RECT 69.300 171.175 69.840 172.780 ;
        RECT 69.300 162.720 69.840 170.465 ;
        RECT 69.300 92.280 69.840 100.280 ;
        RECT 69.300 81.280 69.840 89.280 ;
        RECT 69.300 70.000 69.840 78.280 ;
        RECT 69.300 155.725 69.850 161.220 ;
        RECT 69.300 116.210 69.730 153.550 ;
        RECT 69.300 116.345 69.865 153.425 ;
        RECT 69.300 116.340 69.860 153.430 ;
        RECT 69.300 116.330 69.850 153.440 ;
        RECT 69.300 116.320 69.840 153.450 ;
        RECT 69.300 116.310 69.830 153.460 ;
        RECT 69.300 116.300 69.820 153.470 ;
        RECT 69.300 116.290 69.810 153.480 ;
        RECT 69.300 116.280 69.800 153.490 ;
        RECT 69.300 116.270 69.790 153.500 ;
        RECT 69.300 116.260 69.780 153.510 ;
        RECT 69.300 116.250 69.770 153.520 ;
        RECT 69.300 116.240 69.760 153.530 ;
        RECT 69.300 116.230 69.750 153.540 ;
        RECT 69.300 116.220 69.740 153.550 ;
  END 
END PLBI2F

END LIBRARY
