`timescale 1ns/10ps
`celldefine
module AND2CLKHD1XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2CLKHD2XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2CLKHD3XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2CLKHD4XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2HD1XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2HD1XSPGHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2HD2XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2HD2XSPGHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2HDLXHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2HDMXHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2HDUXHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND3HD1XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (Z, A, B, C);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND3HD2XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (Z, A, B, C);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND3HDLXHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (Z, A, B, C);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND3HDMXHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (Z, A, B, C);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND4HD1XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (Z, A, B, C, D);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND4HD2XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (Z, A, B, C, D);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND4HDLXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (Z, A, B, C, D);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND4HDMXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (Z, A, B, C, D);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI211HD1XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I0_out, A, B);
   or  (I2_out, I0_out, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI211HD2XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I0_out, A, B);
   or  (I2_out, I0_out, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI211HDLXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I0_out, A, B);
   or  (I2_out, I0_out, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI211HDMXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I0_out, A, B);
   or  (I2_out, I0_out, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI21B2HD1XHT (Z, AN, BN, C);
input  AN ;
input  BN ;
input  C ;
output Z ;

   or  (I0_out, AN, BN);
   not (I1_out, I0_out);
   or  (I2_out, I1_out, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI21B2HD2XHT (Z, AN, BN, C);
input  AN ;
input  BN ;
input  C ;
output Z ;

   or  (I0_out, AN, BN);
   not (I1_out, I0_out);
   or  (I2_out, I1_out, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI21B2HDLXHT (Z, AN, BN, C);
input  AN ;
input  BN ;
input  C ;
output Z ;

   or  (I0_out, AN, BN);
   not (I1_out, I0_out);
   or  (I2_out, I1_out, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI21B2HDMXHT (Z, AN, BN, C);
input  AN ;
input  BN ;
input  C ;
output Z ;

   or  (I0_out, AN, BN);
   not (I1_out, I0_out);
   or  (I2_out, I1_out, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI21HD1XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I0_out, A, B);
   or  (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI21HD2XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I0_out, A, B);
   or  (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI21HDLXHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I0_out, A, B);
   or  (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI21HDMXHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I0_out, A, B);
   or  (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI21HDUXHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I0_out, A, B);
   or  (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI221HD1XHT (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   and (I0_out, A, B);
   and (I1_out, C, D);
   or  (I3_out, I0_out, I1_out, E);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI221HD2XHT (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   and (I0_out, A, B);
   and (I1_out, C, D);
   or  (I3_out, I0_out, I1_out, E);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI221HDLXHT (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   and (I0_out, A, B);
   and (I1_out, C, D);
   or  (I3_out, I0_out, I1_out, E);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI221HDMXHT (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   and (I0_out, A, B);
   and (I1_out, C, D);
   or  (I3_out, I0_out, I1_out, E);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI222HD1XHT (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   and (I0_out, E, F);
   and (I1_out, A, B);
   and (I3_out, C, D);
   or  (I4_out, I0_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && E == 1'b0 && F == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI222HD2XHT (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   and (I0_out, E, F);
   and (I1_out, A, B);
   and (I3_out, C, D);
   or  (I4_out, I0_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && E == 1'b0 && F == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI222HDLXHT (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   and (I0_out, E, F);
   and (I1_out, A, B);
   and (I3_out, C, D);
   or  (I4_out, I0_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && E == 1'b0 && F == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI222HDMXHT (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   and (I0_out, E, F);
   and (I1_out, A, B);
   and (I3_out, C, D);
   or  (I4_out, I0_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && E == 1'b0 && F == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI22B2HD1XHT (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, AN, BN);
   not (I1_out, I0_out);
   and (I2_out, C, D);
   or  (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (AN *> Z) = (0, 0);
     ifnone (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (BN *> Z) = (0, 0);
     ifnone (BN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI22B2HD2XHT (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, AN, BN);
   not (I1_out, I0_out);
   and (I2_out, C, D);
   or  (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (AN *> Z) = (0, 0);
     ifnone (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (BN *> Z) = (0, 0);
     ifnone (BN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI22B2HDLXHT (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, AN, BN);
   not (I1_out, I0_out);
   and (I2_out, C, D);
   or  (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (AN *> Z) = (0, 0);
     ifnone (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (BN *> Z) = (0, 0);
     ifnone (BN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI22B2HDMXHT (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, AN, BN);
   not (I1_out, I0_out);
   and (I2_out, C, D);
   or  (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (AN *> Z) = (0, 0);
     ifnone (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (BN *> Z) = (0, 0);
     ifnone (BN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI22HD1XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I0_out, C, D);
   and (I1_out, A, B);
   or  (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI22HD2XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I0_out, A, B);
   and (I1_out, C, D);
   or  (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI22HDLXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I0_out, C, D);
   and (I1_out, A, B);
   or  (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI22HDMXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I0_out, C, D);
   and (I1_out, A, B);
   or  (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI22HDUXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I0_out, C, D);
   and (I1_out, A, B);
   or  (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI31HD1XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I1_out, A, B, C);
   or  (I2_out, I1_out, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI31HD2XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I1_out, A, B, C);
   or  (I2_out, I1_out, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI31HDLXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I1_out, A, B, C);
   or  (I2_out, I1_out, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI31HDMXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I1_out, A, B, C);
   or  (I2_out, I1_out, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI32HD1XHT (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   and (I0_out, D, E);
   and (I2_out, A, B, C);
   or  (I3_out, I0_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI32HD2XHT (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   and (I1_out, A, B, C);
   and (I2_out, D, E);
   or  (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI32HDLXHT (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   and (I0_out, D, E);
   and (I2_out, A, B, C);
   or  (I3_out, I0_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI32HDMXHT (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   and (I0_out, D, E);
   and (I2_out, A, B, C);
   or  (I3_out, I0_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI33HD1XHT (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   and (I1_out, D, E, F);
   and (I3_out, A, B, C);
   or  (I4_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI33HD2XHT (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   and (I1_out, A, B, C);
   and (I3_out, D, E, F);
   or  (I4_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI33HDLXHT (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   and (I1_out, D, E, F);
   and (I3_out, A, B, C);
   or  (I4_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI33HDMXHT (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   and (I1_out, D, E, F);
   and (I3_out, A, B, C);
   or  (I4_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD10XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD12XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD14XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD16XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD1XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD20XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD2XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD30XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD3XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD40XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD4XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD5XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD6XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD7XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD80XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD8XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHDLXHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHDMXHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHDUXHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD12XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD16XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD1XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD20XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD2XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD3XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD4XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD5XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD6XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD7XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD8XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD8XSPGHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHDLXHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHDMXHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHDUXHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD12XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD16XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD1XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD20XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD2XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD3XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD4XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD5XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD6XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD7XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD8XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHDLXHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHDMXHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHDUXHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL1HD1XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL1HDMXHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL1HDMXSPGHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL2HD1XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL2HDMXHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL2HDMXSPGHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL3HD1XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL3HDMXHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL4HD1XHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL4HDMXHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL4HDMXSPGHT (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FAHD1XHT (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // path delays
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (0, 0);
     ifnone (A *> CO) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (0, 0);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (0, 0);
     ifnone (B *> CO) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (0, 0);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (0, 0);
     ifnone (CI *> CO) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (0, 0);
     ifnone (CI *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FAHD2XHT (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // path delays
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (0, 0);
     ifnone (A *> CO) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (0, 0);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (0, 0);
     ifnone (B *> CO) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (0, 0);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (0, 0);
     ifnone (CI *> CO) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (0, 0);
     ifnone (CI *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FAHDLXHT (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // path delays
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (0, 0);
     ifnone (A *> CO) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (0, 0);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (0, 0);
     ifnone (B *> CO) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (0, 0);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (0, 0);
     ifnone (CI *> CO) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (0, 0);
     ifnone (CI *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FAHDMXHT (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // path delays
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (0, 0);
     ifnone (A *> CO) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (0, 0);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (0, 0);
     ifnone (B *> CO) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (0, 0);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (0, 0);
     ifnone (CI *> CO) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (0, 0);
     ifnone (CI *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FAHDUXHT (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // path delays
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (0, 0);
     ifnone (A *> CO) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (0, 0);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (0, 0);
     ifnone (B *> CO) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (0, 0);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (0, 0);
     ifnone (CI *> CO) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (0, 0);
     ifnone (CI *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FAHHD1XHT (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // path delays
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (0, 0);
     ifnone (A *> CO) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (0, 0);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (0, 0);
     ifnone (B *> CO) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (0, 0);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (0, 0);
     ifnone (CI *> CO) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (0, 0);
     ifnone (CI *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FAHHD2XHT (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // path delays
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (0, 0);
     ifnone (A *> CO) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (0, 0);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (0, 0);
     ifnone (B *> CO) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (0, 0);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (0, 0);
     ifnone (CI *> CO) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (0, 0);
     ifnone (CI *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FAHHDLXHT (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // path delays
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (0, 0);
     ifnone (A *> CO) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (0, 0);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (0, 0);
     ifnone (B *> CO) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (0, 0);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (0, 0);
     ifnone (CI *> CO) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (0, 0);
     ifnone (CI *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FAHHDMXHT (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // path delays
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (0, 0);
     ifnone (A *> CO) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (0, 0);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (0, 0);
     ifnone (B *> CO) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (0, 0);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (0, 0);
     ifnone (CI *> CO) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (0, 0);
     ifnone (CI *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDCRHD1XHT (Q, QN, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, 1'b1, dly_RN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDCRHD2XHT (Q, QN, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, 1'b1, dly_RN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDCRHDLXHT (Q, QN, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, 1'b1, dly_RN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDCRHDMXHT (Q, QN, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, 1'b1, dly_RN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDHD1XHT (Q, QN, CK, D);
input  CK ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDHD1XSPGHT (Q, QN, CK, D);
input  CK ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDHD2XHT (Q, QN, CK, D);
input  CK ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDHDLXHT (Q, QN, CK, D);
input  CK ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDHDMXHT (Q, QN, CK, D);
input  CK ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDHQHD1XHT (Q, CK, D);
input  CK ;
input  D ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDHQHD2XHT (Q, CK, D);
input  CK ;
input  D ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDHQHD3XHT (Q, CK, D);
input  CK ;
input  D ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDHQHDMXHT (Q, CK, D);
input  CK ;
input  D ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNHD1XHT (Q, QN, CKN, D);
input  CKN ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     $setuphold(negedge CKN, negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNHD2XHT (Q, QN, CKN, D);
input  CKN ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     $setuphold(negedge CKN, negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNHDLXHT (Q, QN, CKN, D);
input  CKN ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     $setuphold(negedge CKN, negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNHDMXHT (Q, QN, CKN, D);
input  CKN ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     $setuphold(negedge CKN, negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNRHD1XHT (Q, QN, CKN, D, RN);
input  CKN ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNRHD2XHT (Q, QN, CKN, D, RN);
input  CKN ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNRHDLXHT (Q, QN, CKN, D, RN);
input  CKN ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNRHDMXHT (Q, QN, CKN, D, RN);
input  CKN ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNSHD1XHT (Q, QN, CKN, D, SN);
input  CKN ;
input  D ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNSHD2XHT (Q, QN, CKN, D, SN);
input  CKN ;
input  D ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNSHDLXHT (Q, QN, CKN, D, SN);
input  CKN ;
input  D ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNSHDMXHT (Q, QN, CKN, D, SN);
input  CKN ;
input  D ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNSRHD1XHT (Q, QN, CKN, D, RN, SN);
input  CKN ;
input  D ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge CKN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNSRHD2XHT (Q, QN, CKN, D, RN, SN);
input  CKN ;
input  D ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge CKN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNSRHDLXHT (Q, QN, CKN, D, RN, SN);
input  CKN ;
input  D ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge CKN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNSRHDMXHT (Q, QN, CKN, D, RN, SN);
input  CKN ;
input  D ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge CKN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQHD1XHT (Q, CK, D);
input  CK ;
input  D ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQHD2XHT (Q, CK, D);
input  CK ;
input  D ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQHDLXHT (Q, CK, D);
input  CK ;
input  D ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQHDMXHT (Q, CK, D);
input  CK ;
input  D ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQRHD1XHT (Q, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQRHD2XHT (Q, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQRHDLXHT (Q, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQRHDMXHT (Q, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQSHD1XHT (Q, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQSHD2XHT (Q, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQSHDLXHT (Q, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQSHDMXHT (Q, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQSRHD1XHT (Q, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        and _i1 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQSRHD2XHT (Q, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        and _i1 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQSRHDLXHT (Q, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        and _i1 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQSRHDMXHT (Q, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        and _i1 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDRHD1XHT (Q, QN, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDRHD2XHT (Q, QN, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDRHDLXHT (Q, QN, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDRHDMXHT (Q, QN, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDRHQHD1XHT (Q, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDRHQHD2XHT (Q, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDRHQHD3XHT (Q, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDRHQHDMXHT (Q, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSHD1XHT (Q, QN, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSHD2XHT (Q, QN, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSHDLXHT (Q, QN, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSHDMXHT (Q, QN, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSHQHD1XHT (Q, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSHQHD2XHT (Q, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSHQHD3XHT (Q, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSHQHDMXHT (Q, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSRHD1XHT (Q, QN, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSRHD2XHT (Q, QN, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSRHDLXHT (Q, QN, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSRHDMXHT (Q, QN, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSRHQHD1XHT (Q, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        and _i1 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSRHQHD2XHT (Q, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        and _i1 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSRHQHD3XHT (Q, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        and _i1 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSRHQHDMXHT (Q, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        and _i1 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDCRHD1XHT (Q, QN, CK, D, E, RN);
input  CK ;
input  D ;
input  E ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, dly_RN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\E&RN ,E,RN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK &&& \E&RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDCRHD2XHT (Q, QN, CK, D, E, RN);
input  CK ;
input  D ;
input  E ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, dly_RN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\E&RN ,E,RN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK &&& \E&RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDCRHDLXHT (Q, QN, CK, D, E, RN);
input  CK ;
input  D ;
input  E ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, dly_RN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\E&RN ,E,RN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK &&& \E&RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDCRHDMXHT (Q, QN, CK, D, E, RN);
input  CK ;
input  D ;
input  E ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, dly_RN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\E&RN ,E,RN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK &&& \E&RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDHD1XHT (Q, QN, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDHD2XHT (Q, QN, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDHDLXHT (Q, QN, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDHDMXHT (Q, QN, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDHQHD1XHT (Q, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDHQHD2XHT (Q, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDHQHD3XHT (Q, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDHQHDMXHT (Q, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDQHD1XHT (Q, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDQHD2XHT (Q, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDQHDLXHT (Q, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDQHDMXHT (Q, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDCRHD1XHT (Q, QN, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, 1'b1, dly_RN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\RN&~TE ,RN,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDCRHD2XHT (Q, QN, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, 1'b1, dly_RN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\RN&~TE ,RN,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDCRHDLXHT (Q, QN, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, 1'b1, dly_RN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\RN&~TE ,RN,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDCRHDMXHT (Q, QN, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, 1'b1, dly_RN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\RN&~TE ,RN,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDHD1XHT (Q, QN, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDHD1XSPGHT (Q, QN, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDHD2XHT (Q, QN, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDHDLXHT (Q, QN, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDHDMXHT (Q, QN, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDHQHD1XHT (Q, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDHQHD2XHT (Q, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDHQHD3XHT (Q, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDHQHDMXHT (Q, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNHD1XHT (Q, QN, CKN, D, TE, TI);
input  CKN ;
input  D ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNHD2XHT (Q, QN, CKN, D, TE, TI);
input  CKN ;
input  D ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNHDLXHT (Q, QN, CKN, D, TE, TI);
input  CKN ;
input  D ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNHDMXHT (Q, QN, CKN, D, TE, TI);
input  CKN ;
input  D ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNRHD1XHT (Q, QN, CKN, D, RN, TE, TI);
input  CKN ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&~TE ,RN,n1);
        and _i4 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN, posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNRHD2XHT (Q, QN, CKN, D, RN, TE, TI);
input  CKN ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&~TE ,RN,n1);
        and _i4 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN, posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNRHDLXHT (Q, QN, CKN, D, RN, TE, TI);
input  CKN ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&~TE ,RN,n1);
        and _i4 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN, posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNRHDMXHT (Q, QN, CKN, D, RN, TE, TI);
input  CKN ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&~TE ,RN,n1);
        and _i4 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN, posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNSHD1XHT (Q, QN, CKN, D, SN, TE, TI);
input  CKN ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\SN&~TE ,SN,n1);
        and _i4 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN, posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNSHD2XHT (Q, QN, CKN, D, SN, TE, TI);
input  CKN ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\SN&~TE ,SN,n1);
        and _i4 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN, posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNSHDLXHT (Q, QN, CKN, D, SN, TE, TI);
input  CKN ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\SN&~TE ,SN,n1);
        and _i4 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN, posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNSHDMXHT (Q, QN, CKN, D, SN, TE, TI);
input  CKN ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\SN&~TE ,SN,n1);
        and _i4 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN, posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNSRHD1XHT (Q, QN, CKN, D, RN, SN, TE, TI);
input  CKN ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&SN ,RN,SN);
        and _i4 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i5 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge CKN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNSRHD2XHT (Q, QN, CKN, D, RN, SN, TE, TI);
input  CKN ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&SN ,RN,SN);
        and _i4 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i5 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge CKN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNSRHDLXHT (Q, QN, CKN, D, RN, SN, TE, TI);
input  CKN ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&SN ,RN,SN);
        and _i4 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i5 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge CKN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNSRHDMXHT (Q, QN, CKN, D, RN, SN, TE, TI);
input  CKN ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&SN ,RN,SN);
        and _i4 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i5 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge CKN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQHD1XHT (Q, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQHD2XHT (Q, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQHDLXHT (Q, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQHDMXHT (Q, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQRHD1XHT (Q, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&~TE ,RN,n1);
        and _i3 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQRHD2XHT (Q, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&~TE ,RN,n1);
        and _i3 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQRHDLXHT (Q, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&~TE ,RN,n1);
        and _i3 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQRHDMXHT (Q, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&~TE ,RN,n1);
        and _i3 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQSHD1XHT (Q, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\SN&~TE ,SN,n1);
        and _i3 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQSHD2XHT (Q, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\SN&~TE ,SN,n1);
        and _i3 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQSHDLXHT (Q, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\SN&~TE ,SN,n1);
        and _i3 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQSHDMXHT (Q, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\SN&~TE ,SN,n1);
        and _i3 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQSRHD1XHT (Q, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&SN ,RN,SN);
        and _i3 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i4 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQSRHD2XHT (Q, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&SN ,RN,SN);
        and _i3 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i4 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQSRHDLXHT (Q, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&SN ,RN,SN);
        and _i3 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i4 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQSRHDMXHT (Q, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&SN ,RN,SN);
        and _i3 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i4 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDRHD1XHT (Q, QN, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&~TE ,RN,n1);
        and _i4 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDRHD2XHT (Q, QN, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&~TE ,RN,n1);
        and _i4 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDRHDLXHT (Q, QN, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&~TE ,RN,n1);
        and _i4 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDRHDMXHT (Q, QN, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&~TE ,RN,n1);
        and _i4 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDRHQHD1XHT (Q, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&~TE ,RN,n1);
        and _i3 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDRHQHD2XHT (Q, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&~TE ,RN,n1);
        and _i3 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDRHQHD3XHT (Q, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&~TE ,RN,n1);
        and _i3 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDRHQHDMXHT (Q, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&~TE ,RN,n1);
        and _i3 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSHD1XHT (Q, QN, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\SN&~TE ,SN,n1);
        and _i4 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSHD2XHT (Q, QN, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\SN&~TE ,SN,n1);
        and _i4 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSHDLXHT (Q, QN, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\SN&~TE ,SN,n1);
        and _i4 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSHDMXHT (Q, QN, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\SN&~TE ,SN,n1);
        and _i4 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSHQHD1XHT (Q, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\SN&~TE ,SN,n1);
        and _i3 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSHQHD2XHT (Q, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\SN&~TE ,SN,n1);
        and _i3 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSHQHD3XHT (Q, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\SN&~TE ,SN,n1);
        and _i3 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSHQHDMXHT (Q, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\SN&~TE ,SN,n1);
        and _i3 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSRHD1XHT (Q, QN, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&SN ,RN,SN);
        and _i4 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i5 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSRHD2XHT (Q, QN, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&SN ,RN,SN);
        and _i4 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i5 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSRHDLXHT (Q, QN, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&SN ,RN,SN);
        and _i4 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i5 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSRHDMXHT (Q, QN, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&SN ,RN,SN);
        and _i4 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i5 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSRHQHD1XHT (Q, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&SN ,RN,SN);
        and _i3 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i4 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSRHQHD2XHT (Q, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&SN ,RN,SN);
        and _i3 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i4 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSRHQHD3XHT (Q, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&SN ,RN,SN);
        and _i3 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i4 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSRHQHDMXHT (Q, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&SN ,RN,SN);
        and _i3 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i4 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDCRHD1XHT (Q, QN, CK, D, E, RN, TE, TI);
input  CK ;
input  D ;
input  E ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, dly_RN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\RN&~TE ,RN,\~TE );
        and _i4 (\E&RN&~TE ,E,\RN&~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& \~TE , negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& \~TE , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDCRHD2XHT (Q, QN, CK, D, E, RN, TE, TI);
input  CK ;
input  D ;
input  E ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, dly_RN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\RN&~TE ,RN,\~TE );
        and _i4 (\E&RN&~TE ,E,\RN&~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& \~TE , negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& \~TE , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDCRHDLXHT (Q, QN, CK, D, E, RN, TE, TI);
input  CK ;
input  D ;
input  E ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, dly_RN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\RN&~TE ,RN,\~TE );
        and _i4 (\E&RN&~TE ,E,\RN&~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& \~TE , negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& \~TE , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDCRHDMXHT (Q, QN, CK, D, E, RN, TE, TI);
input  CK ;
input  D ;
input  E ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, dly_RN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\RN&~TE ,RN,\~TE );
        and _i4 (\E&RN&~TE ,E,\RN&~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& \~TE , negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& \~TE , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDHD1XHT (Q, QN, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDHD2XHT (Q, QN, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDHDLXHT (Q, QN, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDHDMXHT (Q, QN, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDHQHD1XHT (Q, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
        and _i2 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDHQHD2XHT (Q, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
        and _i2 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDHQHD3XHT (Q, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
        and _i2 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDHQHDMXHT (Q, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
        and _i2 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDQHD1XHT (Q, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
        and _i2 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDQHD2XHT (Q, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
        and _i2 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDQHDLXHT (Q, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
        and _i2 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDQHDMXHT (Q, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
        and _i2 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module HAHD1XHT (CO, S, A, B);
input  A ;
input  B ;
output CO ;
output S ;

   and (CO, A, B);
   xor (S, A, B);

   specify
     // path delays
     (A *> CO) = (0, 0);
     if (B == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b1)
       (A *> S) = (0, 0);
     (B *> CO) = (0, 0);
     if (A == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b1)
       (B *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module HAHD2XHT (CO, S, A, B);
input  A ;
input  B ;
output CO ;
output S ;

   and (CO, A, B);
   xor (S, A, B);

   specify
     // path delays
     (A *> CO) = (0, 0);
     if (B == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b1)
       (A *> S) = (0, 0);
     (B *> CO) = (0, 0);
     if (A == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b1)
       (B *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module HAHDLXHT (CO, S, A, B);
input  A ;
input  B ;
output CO ;
output S ;

   and (CO, A, B);
   xor (S, A, B);

   specify
     // path delays
     (A *> CO) = (0, 0);
     if (B == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b1)
       (A *> S) = (0, 0);
     (B *> CO) = (0, 0);
     if (A == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b1)
       (B *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module HAHDMXHT (CO, S, A, B);
input  A ;
input  B ;
output CO ;
output S ;

   and (CO, A, B);
   xor (S, A, B);

   specify
     // path delays
     (A *> CO) = (0, 0);
     if (B == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b1)
       (A *> S) = (0, 0);
     (B *> CO) = (0, 0);
     if (A == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b1)
       (B *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module HOLDHDHT (Z);
inout  Z ;

   not (weak1,weak0) _i0(Z,DUMMY);
   not _i1 (DUMMY,Z);


endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD10XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD12XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD14XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD16XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD1XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD20XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD2XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD30XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD3XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD40XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD4XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD5XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD6XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD7XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD80XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD8XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHDLXHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHDMXHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHDUXHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD12XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD16XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD1XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD1XSPGHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD20XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD2XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD3XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD4XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD5XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD6XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD7XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD8XHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHDLXHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHDMXHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHDPXHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHDUXHT (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD12XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD16XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD1XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD20XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD2XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD3XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD4XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD5XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD6XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD7XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD8XHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHDLXHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHDMXHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHDUXHT (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATHD1XHT (Q, QN, D, G);
input  D ;
input  G ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G, 1'b1, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     $setuphold(negedge G, negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $width(posedge G, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATHD1XSPGHT (Q, QN, D, G);
input  D ;
input  G ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G, 1'b1, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     $setuphold(negedge G, negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $width(posedge G, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATHD2XHT (Q, QN, D, G);
input  D ;
input  G ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G, 1'b1, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     $setuphold(negedge G, negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $width(posedge G, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATHDLXHT (Q, QN, D, G);
input  D ;
input  G ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G, 1'b1, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     $setuphold(negedge G, negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $width(posedge G, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATHDMXHT (Q, QN, D, G);
input  D ;
input  G ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G, 1'b1, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     $setuphold(negedge G, negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $width(posedge G, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNHD1XHT (Q, QN, D, GN);
input  D ;
input  GN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN, 1'b1, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     $setuphold(posedge GN, negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $width(negedge GN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNHD2XHT (Q, QN, D, GN);
input  D ;
input  GN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN, 1'b1, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     $setuphold(posedge GN, negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $width(negedge GN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNHDLXHT (Q, QN, D, GN);
input  D ;
input  GN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN, 1'b1, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     $setuphold(posedge GN, negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $width(negedge GN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNHDMXHT (Q, QN, D, GN);
input  D ;
input  GN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN, 1'b1, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     $setuphold(posedge GN, negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $width(negedge GN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNRHD1XHT (Q, QN, D, GN, RN);
input  D ;
input  GN ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN, 1'b1,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge GN &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge RN, 0, 0, NOTIFIER, , , dly_GN, dly_RN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNRHD2XHT (Q, QN, D, GN, RN);
input  D ;
input  GN ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN, 1'b1,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge GN &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge RN, 0, 0, NOTIFIER, , , dly_GN, dly_RN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNRHDLXHT (Q, QN, D, GN, RN);
input  D ;
input  GN ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN, 1'b1,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge GN &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge RN, 0, 0, NOTIFIER, , , dly_GN, dly_RN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNRHDMXHT (Q, QN, D, GN, RN);
input  D ;
input  GN ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN, 1'b1,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge GN &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge RN, 0, 0, NOTIFIER, , , dly_GN, dly_RN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNSHD1XHT (Q, QN, D, GN, SN);
input  D ;
input  GN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN,dly_SN, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge GN &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge SN, 0, 0, NOTIFIER, , , dly_GN, dly_SN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNSHD2XHT (Q, QN, D, GN, SN);
input  D ;
input  GN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN,dly_SN, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge GN &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge SN, 0, 0, NOTIFIER, , , dly_GN, dly_SN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNSHDLXHT (Q, QN, D, GN, SN);
input  D ;
input  GN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN,dly_SN, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge GN &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge SN, 0, 0, NOTIFIER, , , dly_GN, dly_SN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNSHDMXHT (Q, QN, D, GN, SN);
input  D ;
input  GN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN,dly_SN, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge GN &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge SN, 0, 0, NOTIFIER, , , dly_GN, dly_SN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNSRHD1XHT (Q, QN, D, GN, RN, SN);
input  D ;
input  GN ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN,dly_SN,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge GN &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_GN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge GN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_GN, dly_SN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNSRHD2XHT (Q, QN, D, GN, RN, SN);
input  D ;
input  GN ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN,dly_SN,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge GN &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_GN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge GN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_GN, dly_SN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNSRHDLXHT (Q, QN, D, GN, RN, SN);
input  D ;
input  GN ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN,dly_SN,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge GN &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_GN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge GN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_GN, dly_SN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNSRHDMXHT (Q, QN, D, GN, RN, SN);
input  D ;
input  GN ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN,dly_SN,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge GN &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_GN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge GN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_GN, dly_SN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATRHD1XHT (Q, QN, D, G, RN);
input  D ;
input  G ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G, 1'b1, dly_RN,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge G &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge RN, 0, 0, NOTIFIER, , , dly_G, dly_RN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATRHD2XHT (Q, QN, D, G, RN);
input  D ;
input  G ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G, 1'b1, dly_RN,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge G &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge RN, 0, 0, NOTIFIER, , , dly_G, dly_RN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATRHDLXHT (Q, QN, D, G, RN);
input  D ;
input  G ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G, 1'b1, dly_RN,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge G &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge RN, 0, 0, NOTIFIER, , , dly_G, dly_RN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATRHDMXHT (Q, QN, D, G, RN);
input  D ;
input  G ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G, 1'b1, dly_RN,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge G &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge RN, 0, 0, NOTIFIER, , , dly_G, dly_RN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATSHD1XHT (Q, QN, D, G, SN);
input  D ;
input  G ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G,dly_SN, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge G &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge SN, 0, 0, NOTIFIER, , , dly_G, dly_SN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATSHD2XHT (Q, QN, D, G, SN);
input  D ;
input  G ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G,dly_SN, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge G &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge SN, 0, 0, NOTIFIER, , , dly_G, dly_SN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATSHDLXHT (Q, QN, D, G, SN);
input  D ;
input  G ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G,dly_SN, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge G &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge SN, 0, 0, NOTIFIER, , , dly_G, dly_SN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATSHDMXHT (Q, QN, D, G, SN);
input  D ;
input  G ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G,dly_SN, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge G &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge SN, 0, 0, NOTIFIER, , , dly_G, dly_SN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATSRHD1XHT (Q, QN, D, G, RN, SN);
input  D ;
input  G ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G,dly_SN,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge G &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_G, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge G &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_G, dly_SN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATSRHD2XHT (Q, QN, D, G, RN, SN);
input  D ;
input  G ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G,dly_SN,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge G &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_G, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge G &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_G, dly_SN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATSRHDLXHT (Q, QN, D, G, RN, SN);
input  D ;
input  G ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G,dly_SN,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge G &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_G, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge G &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_G, dly_SN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATSRHDMXHT (Q, QN, D, G, RN, SN);
input  D ;
input  G ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G,dly_SN,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge G &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_G, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge G &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_G, dly_SN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATTSHD1XHT (Q, D, E, G);
input  D ;
input  E ;
input  G ;
output Q ;
reg NOTIFIER ;
        ip_latchsr _i0 (_n1, dly_D, dly_G, 1'b1, 1'b1, NOTIFIER);
        bufif1 _i1 (Q, _n1, E);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (E *> Q) = (0, 0, 0, 0, 0, 0);
     (G *> Q) = (0, 0);
     $setuphold(negedge G, negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $width(posedge G, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATTSHD2XHT (Q, D, E, G);
input  D ;
input  E ;
input  G ;
output Q ;
reg NOTIFIER ;
        ip_latchsr _i0 (_n1, dly_D, dly_G, 1'b1, 1'b1, NOTIFIER);
        bufif1 _i1 (Q, _n1, E);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (E *> Q) = (0, 0, 0, 0, 0, 0);
     (G *> Q) = (0, 0);
     $setuphold(negedge G, negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $width(posedge G, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATTSHDLXHT (Q, D, E, G);
input  D ;
input  E ;
input  G ;
output Q ;
reg NOTIFIER ;
        ip_latchsr _i0 (_n1, dly_D, dly_G, 1'b1, 1'b1, NOTIFIER);
        bufif1 _i1 (Q, _n1, E);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (E *> Q) = (0, 0, 0, 0, 0, 0);
     (G *> Q) = (0, 0);
     $setuphold(negedge G, negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $width(posedge G, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATTSHDMXHT (Q, D, E, G);
input  D ;
input  E ;
input  G ;
output Q ;
reg NOTIFIER ;
        ip_latchsr _i0 (_n1, dly_D, dly_G, 1'b1, 1'b1, NOTIFIER);
        bufif1 _i1 (Q, _n1, E);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (E *> Q) = (0, 0, 0, 0, 0, 0);
     (G *> Q) = (0, 0);
     $setuphold(negedge G, negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $width(posedge G, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2CLKHD1XHT (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2CLKHD2XHT (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2CLKHD3XHT (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2CLKHD4XHT (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2HD1XHT (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2HD1XSPGHT (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2HD2XHT (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2HD3XHT (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2HDLXHT (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2HDMXHT (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2HDUXHT (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX4HD1XHT (Z, A, B, C, D, S0, S1);
input  A ;
input  B ;
input  C ;
input  D ;
input  S0 ;
input  S1 ;
output Z ;

   udp_mux2 (I0_out, C, D, S0);
   udp_mux2 (I1_out, A, B, S0);
   udp_mux2 (Z, I1_out, I0_out, S1);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     ifnone (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX4HD2XHT (Z, A, B, C, D, S0, S1);
input  A ;
input  B ;
input  C ;
input  D ;
input  S0 ;
input  S1 ;
output Z ;

   udp_mux2 (I0_out, C, D, S0);
   udp_mux2 (I1_out, A, B, S0);
   udp_mux2 (Z, I1_out, I0_out, S1);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     ifnone (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX4HDLXHT (Z, A, B, C, D, S0, S1);
input  A ;
input  B ;
input  C ;
input  D ;
input  S0 ;
input  S1 ;
output Z ;

   udp_mux2 (I0_out, C, D, S0);
   udp_mux2 (I1_out, A, B, S0);
   udp_mux2 (Z, I1_out, I0_out, S1);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     ifnone (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX4HDMXHT (Z, A, B, C, D, S0, S1);
input  A ;
input  B ;
input  C ;
input  D ;
input  S0 ;
input  S1 ;
output Z ;

   udp_mux2 (I0_out, C, D, S0);
   udp_mux2 (I1_out, A, B, S0);
   udp_mux2 (Z, I1_out, I0_out, S1);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     ifnone (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUXI2HD1XHT (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (I0_out, A, B, S0);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUXI2HD2XHT (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (I0_out, A, B, S0);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUXI2HD3XHT (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (I0_out, A, B, S0);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUXI2HDLXHT (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (I0_out, A, B, S0);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUXI2HDMXHT (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (I0_out, A, B, S0);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUXI4HD1XHT (Z, A, B, C, D, S0, S1);
input  A ;
input  B ;
input  C ;
input  D ;
input  S0 ;
input  S1 ;
output Z ;

   udp_mux2 (I0_out, C, D, S0);
   udp_mux2 (I1_out, A, B, S0);
   udp_mux2 (I2_out, I1_out, I0_out, S1);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     ifnone (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUXI4HD2XHT (Z, A, B, C, D, S0, S1);
input  A ;
input  B ;
input  C ;
input  D ;
input  S0 ;
input  S1 ;
output Z ;

   udp_mux2 (I0_out, C, D, S0);
   udp_mux2 (I1_out, A, B, S0);
   udp_mux2 (I2_out, I1_out, I0_out, S1);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     ifnone (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUXI4HDLXHT (Z, A, B, C, D, S0, S1);
input  A ;
input  B ;
input  C ;
input  D ;
input  S0 ;
input  S1 ;
output Z ;

   udp_mux2 (I0_out, C, D, S0);
   udp_mux2 (I1_out, A, B, S0);
   udp_mux2 (I2_out, I1_out, I0_out, S1);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     ifnone (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUXI4HDMXHT (Z, A, B, C, D, S0, S1);
input  A ;
input  B ;
input  C ;
input  D ;
input  S0 ;
input  S1 ;
output Z ;

   udp_mux2 (I0_out, C, D, S0);
   udp_mux2 (I1_out, A, B, S0);
   udp_mux2 (I2_out, I1_out, I0_out, S1);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     ifnone (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2B1HD1XHT (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   and (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2B1HD2XHT (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   and (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2B1HDLXHT (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   and (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2B1HDMXHT (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   and (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2B1HDUXHT (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   and (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2HD1XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2HD1XSPGHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2HD2XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2HD2XSPGHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2HD3XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2HDLXHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2HDMXHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2HDUXHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3B1HD1XHT (Z, AN, B, C);
input  AN ;
input  B ;
input  C ;
output Z ;

   not (I0_out, AN);
   and (I2_out, I0_out, B, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3B1HD2XHT (Z, AN, B, C);
input  AN ;
input  B ;
input  C ;
output Z ;

   not (I0_out, AN);
   and (I2_out, I0_out, B, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3B1HDLXHT (Z, AN, B, C);
input  AN ;
input  B ;
input  C ;
output Z ;

   not (I0_out, AN);
   and (I2_out, I0_out, B, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3B1HDMXHT (Z, AN, B, C);
input  AN ;
input  B ;
input  C ;
output Z ;

   not (I0_out, AN);
   and (I2_out, I0_out, B, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3HD1XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3HD2XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3HD3XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3HDLXHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3HDMXHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4B1HD1XHT (Z, AN, B, C, D);
input  AN ;
input  B ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   and (I3_out, I0_out, B, C, D);
   not (Z, I3_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4B1HD2XHT (Z, AN, B, C, D);
input  AN ;
input  B ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   and (I3_out, I0_out, B, C, D);
   not (Z, I3_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4B1HDLXHT (Z, AN, B, C, D);
input  AN ;
input  B ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   and (I3_out, I0_out, B, C, D);
   not (Z, I3_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4B1HDMXHT (Z, AN, B, C, D);
input  AN ;
input  B ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   and (I3_out, I0_out, B, C, D);
   not (Z, I3_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4B2HD1XHT (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   not (I0_out, BN);
   not (I1_out, AN);
   and (I4_out, I0_out, I1_out, C, D);
   not (Z, I4_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4B2HD2XHT (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   not (I0_out, BN);
   not (I1_out, AN);
   and (I4_out, I0_out, I1_out, C, D);
   not (Z, I4_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4B2HDLXHT (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   not (I1_out, BN);
   and (I4_out, I0_out, I1_out, C, D);
   not (Z, I4_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4B2HDMXHT (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   not (I1_out, BN);
   and (I4_out, I0_out, I1_out, C, D);
   not (Z, I4_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4HD1XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4HD2XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4HD3XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4HDLXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4HDMXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2B1HD1XHT (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   or  (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2B1HD2XHT (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   or  (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2B1HDLXHT (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   or  (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2B1HDMXHT (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   or  (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2B1HDUXHT (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   or  (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2HD1XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2HD1XSPGHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2HD2XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2HD2XSPGHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2HD3XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2HDLXHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2HDMXHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2HDUXHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR3B1HD1XHT (Z, AN, B, C);
input  AN ;
input  B ;
input  C ;
output Z ;

   not (I0_out, AN);
   or  (I2_out, I0_out, B, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR3B1HD2XHT (Z, AN, B, C);
input  AN ;
input  B ;
input  C ;
output Z ;

   not (I0_out, AN);
   or  (I2_out, I0_out, B, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR3B1HDLXHT (Z, AN, B, C);
input  AN ;
input  B ;
input  C ;
output Z ;

   not (I0_out, AN);
   or  (I2_out, I0_out, B, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR3B1HDMXHT (Z, AN, B, C);
input  AN ;
input  B ;
input  C ;
output Z ;

   not (I0_out, AN);
   or  (I2_out, I0_out, B, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR3HD1XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR3HD2XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR3HD3XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR3HDLXHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR3HDMXHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4B1HD1XHT (Z, AN, B, C, D);
input  AN ;
input  B ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   or  (I3_out, I0_out, B, C, D);
   not (Z, I3_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4B1HD2XHT (Z, AN, B, C, D);
input  AN ;
input  B ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   or  (I3_out, I0_out, B, C, D);
   not (Z, I3_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4B1HDLXHT (Z, AN, B, C, D);
input  AN ;
input  B ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   or  (I3_out, I0_out, B, C, D);
   not (Z, I3_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4B1HDMXHT (Z, AN, B, C, D);
input  AN ;
input  B ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   or  (I3_out, I0_out, B, C, D);
   not (Z, I3_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4B2HD1XHT (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   not (I0_out, BN);
   not (I1_out, AN);
   or  (I4_out, I0_out, I1_out, C, D);
   not (Z, I4_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4B2HD2XHT (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   not (I0_out, BN);
   not (I1_out, AN);
   or  (I4_out, I0_out, I1_out, C, D);
   not (Z, I4_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4B2HDLXHT (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   not (I0_out, BN);
   not (I1_out, AN);
   or  (I4_out, I0_out, I1_out, C, D);
   not (Z, I4_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4B2HDMXHT (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   not (I0_out, BN);
   not (I1_out, AN);
   or  (I4_out, I0_out, I1_out, C, D);
   not (Z, I4_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4HD1XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4HD2XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4HD3XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4HDLXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4HDMXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI211HD1XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, A, B);
   and (I2_out, I0_out, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI211HD2XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, A, B);
   and (I2_out, I0_out, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI211HDLXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, A, B);
   and (I2_out, I0_out, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI211HDMXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, A, B);
   and (I2_out, I0_out, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI21B2HD1XHT (Z, AN, BN, C);
input  AN ;
input  BN ;
input  C ;
output Z ;

   and (I0_out, AN, BN);
   not (I1_out, I0_out);
   and (I2_out, I1_out, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI21B2HD2XHT (Z, AN, BN, C);
input  AN ;
input  BN ;
input  C ;
output Z ;

   and (I0_out, AN, BN);
   not (I1_out, I0_out);
   and (I2_out, I1_out, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI21B2HDLXHT (Z, AN, BN, C);
input  AN ;
input  BN ;
input  C ;
output Z ;

   and (I0_out, AN, BN);
   not (I1_out, I0_out);
   and (I2_out, I1_out, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI21B2HDMXHT (Z, AN, BN, C);
input  AN ;
input  BN ;
input  C ;
output Z ;

   and (I0_out, AN, BN);
   not (I1_out, I0_out);
   and (I2_out, I1_out, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI21HD1XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I0_out, A, B);
   and (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI21HD2XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I0_out, A, B);
   and (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI21HDLXHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I0_out, A, B);
   and (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI21HDMXHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I0_out, A, B);
   and (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI21HDUXHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I0_out, A, B);
   and (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI221HD1XHT (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   or  (I0_out, A, B);
   or  (I1_out, C, D);
   and (I3_out, I0_out, I1_out, E);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI221HD2XHT (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   or  (I0_out, A, B);
   or  (I1_out, C, D);
   and (I3_out, I0_out, I1_out, E);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI221HDLXHT (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   or  (I0_out, A, B);
   or  (I1_out, C, D);
   and (I3_out, I0_out, I1_out, E);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI221HDMXHT (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   or  (I0_out, A, B);
   or  (I1_out, C, D);
   and (I3_out, I0_out, I1_out, E);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI222HD1XHT (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   or  (I0_out, A, B);
   or  (I1_out, E, F);
   or  (I3_out, C, D);
   and (I4_out, I0_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && E == 1'b1 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI222HD2XHT (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   or  (I0_out, A, B);
   or  (I1_out, C, D);
   or  (I3_out, E, F);
   and (I4_out, I0_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && E == 1'b1 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI222HDLXHT (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   or  (I0_out, A, B);
   or  (I1_out, E, F);
   or  (I3_out, C, D);
   and (I4_out, I0_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && E == 1'b1 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI222HDMXHT (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   or  (I0_out, A, B);
   or  (I1_out, E, F);
   or  (I3_out, C, D);
   and (I4_out, I0_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && E == 1'b1 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI22B2HD1XHT (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   and (I0_out, AN, BN);
   not (I1_out, I0_out);
   or  (I2_out, C, D);
   and (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (AN *> Z) = (0, 0);
     ifnone (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (BN *> Z) = (0, 0);
     ifnone (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI22B2HD2XHT (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   and (I0_out, AN, BN);
   not (I1_out, I0_out);
   or  (I2_out, C, D);
   and (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (AN *> Z) = (0, 0);
     ifnone (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (BN *> Z) = (0, 0);
     ifnone (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI22B2HDLXHT (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   and (I0_out, AN, BN);
   not (I1_out, I0_out);
   or  (I2_out, C, D);
   and (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (AN *> Z) = (0, 0);
     ifnone (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (BN *> Z) = (0, 0);
     ifnone (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI22B2HDMXHT (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   and (I0_out, AN, BN);
   not (I1_out, I0_out);
   or  (I2_out, C, D);
   and (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (AN *> Z) = (0, 0);
     ifnone (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (BN *> Z) = (0, 0);
     ifnone (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI22HD1XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, C, D);
   or  (I1_out, A, B);
   and (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI22HD2XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, A, B);
   or  (I1_out, C, D);
   and (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI22HDLXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, C, D);
   or  (I1_out, A, B);
   and (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI22HDMXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, C, D);
   or  (I1_out, A, B);
   and (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI22HDUXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, C, D);
   or  (I1_out, A, B);
   and (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI31HD1XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I1_out, A, B, C);
   and (I2_out, I1_out, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI31HD2XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I1_out, A, B, C);
   and (I2_out, I1_out, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI31HDLXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I1_out, A, B, C);
   and (I2_out, I1_out, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI31HDMXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I1_out, A, B, C);
   and (I2_out, I1_out, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI32HD1XHT (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   or  (I1_out, A, B, C);
   or  (I2_out, D, E);
   and (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI32HD2XHT (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   or  (I1_out, A, B, C);
   or  (I2_out, D, E);
   and (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI32HDLXHT (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   or  (I0_out, D, E);
   or  (I2_out, A, B, C);
   and (I3_out, I0_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI32HDMXHT (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   or  (I0_out, D, E);
   or  (I2_out, A, B, C);
   and (I3_out, I0_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI33HD1XHT (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   or  (I1_out, A, B, C);
   or  (I3_out, D, E, F);
   and (I4_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI33HD2XHT (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   or  (I1_out, A, B, C);
   or  (I3_out, D, E, F);
   and (I4_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI33HDLXHT (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   or  (I1_out, D, E, F);
   or  (I3_out, A, B, C);
   and (I4_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI33HDMXHT (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   or  (I1_out, D, E, F);
   or  (I3_out, A, B, C);
   and (I4_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR2HD1XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR2HD1XSPGHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR2HD2XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR2HD2XSPGHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR2HDLXHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR2HDMXHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR2HDUXHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR3HD1XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (Z, A, B, C);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR3HD2XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (Z, A, B, C);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR3HDLXHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (Z, A, B, C);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR3HDMXHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (Z, A, B, C);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR4HD1XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (Z, A, B, C, D);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR4HD2XHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (Z, A, B, C, D);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR4HDLXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (Z, A, B, C, D);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR4HDMXHT (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (Z, A, B, C, D);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module PULLDHDHT (Z, EN);
        output Z;
        input  EN;
        bufif0 _i0 (Z, 1'b0, EN);
        specify

                (EN => Z) = (0,0,0,0,0,0);
        endspecify
endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module PULLUHDHT (Z, E);
        output Z;
        input  E;
        bufif1 _i0 (Z, 1'b1, E);
        specify

                (E => Z) = (0,0,0,0,0,0);
        endspecify
endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RSLATHD1XHT (Q, QN, R, S);
input  R ;
input  S ;
output Q ;
output QN ;
reg NOTIFIER ;
        rslat _i0 (q,dly_R,dly_S,NOTIFIER);
        rslatn _i1 (qn,dly_R,dly_S,NOTIFIER);
        buf _i2 (QN,qn);
        buf _i3 (Q,q);
   specify
     // path delays
     (R *> Q) = (0, 0);
     (R *> QN) = (0, 0);
     (S *> Q) = (0, 0);
     (S *> QN) = (0, 0);
     $setuphold(negedge S, negedge R, 0, 0, NOTIFIER, , , dly_S, dly_R);
     $setuphold(negedge R, negedge S, 0, 0, NOTIFIER, , , dly_R, dly_S);
     $width(posedge R, 0, 0, NOTIFIER);
     $width(posedge S, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RSLATHD2XHT (Q, QN, R, S);
input  R ;
input  S ;
output Q ;
output QN ;
reg NOTIFIER ;
        rslat _i0 (q,dly_R,dly_S,NOTIFIER);
        rslatn _i1 (qn,dly_R,dly_S,NOTIFIER);
        buf _i2 (QN,qn);
        buf _i3 (Q,q);
   specify
     // path delays
     (R *> Q) = (0, 0);
     (R *> QN) = (0, 0);
     (S *> Q) = (0, 0);
     (S *> QN) = (0, 0);
     $setuphold(negedge S, negedge R, 0, 0, NOTIFIER, , , dly_S, dly_R);
     $setuphold(negedge R, negedge S, 0, 0, NOTIFIER, , , dly_R, dly_S);
     $width(posedge R, 0, 0, NOTIFIER);
     $width(posedge S, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RSLATHDLXHT (Q, QN, R, S);
input  R ;
input  S ;
output Q ;
output QN ;
reg NOTIFIER ;
        rslat _i0 (q,dly_R,dly_S,NOTIFIER);
        rslatn _i1 (qn,dly_R,dly_S,NOTIFIER);
        buf _i2 (QN,qn);
        buf _i3 (Q,q);
   specify
     // path delays
     (R *> Q) = (0, 0);
     (R *> QN) = (0, 0);
     (S *> Q) = (0, 0);
     (S *> QN) = (0, 0);
     $setuphold(negedge S, negedge R, 0, 0, NOTIFIER, , , dly_S, dly_R);
     $setuphold(negedge R, negedge S, 0, 0, NOTIFIER, , , dly_R, dly_S);
     $width(posedge R, 0, 0, NOTIFIER);
     $width(posedge S, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RSLATHDMXHT (Q, QN, R, S);
input  R ;
input  S ;
output Q ;
output QN ;
reg NOTIFIER ;
        rslat _i0 (q,dly_R,dly_S,NOTIFIER);
        rslatn _i1 (qn,dly_R,dly_S,NOTIFIER);
        buf _i2 (QN,qn);
        buf _i3 (Q,q);
   specify
     // path delays
     (R *> Q) = (0, 0);
     (R *> QN) = (0, 0);
     (S *> Q) = (0, 0);
     (S *> QN) = (0, 0);
     $setuphold(negedge S, negedge R, 0, 0, NOTIFIER, , , dly_S, dly_R);
     $setuphold(negedge R, negedge S, 0, 0, NOTIFIER, , , dly_R, dly_S);
     $width(posedge R, 0, 0, NOTIFIER);
     $width(posedge S, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RSLATNHD1XHT (Q, QN, RN, SN);
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        rsblat _i0 (q,dly_RN,dly_SN,NOTIFIER);
        rsblatn _i1 (qn,dly_RN,dly_SN,NOTIFIER);
        buf _i2 (QN,qn);
        buf _i3 (Q,q);
   specify
     // path delays
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge SN, posedge RN, 0, 0, NOTIFIER, , , dly_SN, dly_RN);
     $setuphold(posedge RN, posedge SN, 0, 0, NOTIFIER, , , dly_RN, dly_SN);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RSLATNHD2XHT (Q, QN, RN, SN);
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        rsblat _i0 (q,dly_RN,dly_SN,NOTIFIER);
        rsblatn _i1 (qn,dly_RN,dly_SN,NOTIFIER);
        buf _i2 (QN,qn);
        buf _i3 (Q,q);
   specify
     // path delays
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge SN, posedge RN, 0, 0, NOTIFIER, , , dly_SN, dly_RN);
     $setuphold(posedge RN, posedge SN, 0, 0, NOTIFIER, , , dly_RN, dly_SN);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RSLATNHDLXHT (Q, QN, RN, SN);
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        rsblat _i0 (q,dly_RN,dly_SN,NOTIFIER);
        rsblatn _i1 (qn,dly_RN,dly_SN,NOTIFIER);
        buf _i2 (QN,qn);
        buf _i3 (Q,q);
   specify
     // path delays
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge SN, posedge RN, 0, 0, NOTIFIER, , , dly_SN, dly_RN);
     $setuphold(posedge RN, posedge SN, 0, 0, NOTIFIER, , , dly_RN, dly_SN);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RSLATNHDMXHT (Q, QN, RN, SN);
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        rsblat _i0 (q,dly_RN,dly_SN,NOTIFIER);
        rsblatn _i1 (qn,dly_RN,dly_SN,NOTIFIER);
        buf _i2 (QN,qn);
        buf _i3 (Q,q);
   specify
     // path delays
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge SN, posedge RN, 0, 0, NOTIFIER, , , dly_SN, dly_RN);
     $setuphold(posedge RN, posedge SN, 0, 0, NOTIFIER, , , dly_RN, dly_SN);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module TIEHHDHT (Z);
output Z ;

   buf (Z, 1'B1);


endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module TIELHDHT (Z);
output Z ;

   buf (Z, 1'B0);


endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR2HD1XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR2HD2XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR2HD3XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR2HDLXHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR2HDMXHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR3HD1XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR3HD2XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR3HD3XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR3HDLXHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR3HDMXHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR2CLKHD1XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (Z, A, B);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR2CLKHD2XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (Z, A, B);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR2CLKHD3XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (Z, A, B);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR2CLKHD4XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (Z, A, B);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR2HD1XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (Z, A, B);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR2HD2XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (Z, A, B);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR2HD3XHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (Z, A, B);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR2HDLXHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (Z, A, B);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR2HDMXHT (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (Z, A, B);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR3HD1XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (Z, I0_out, C);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR3HD2XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (Z, I0_out, C);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR3HD3XHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (Z, I0_out, C);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR3HDLXHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (Z, I0_out, C);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR3HDMXHT (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (Z, I0_out, C);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVODHD8XHT (Z0, Z1, Z2, Z3, Z4, Z5, Z6, Z7, A);
	output Z0;
	output Z1;
	output Z2;
	output Z3;
	output Z4;
	output Z5;
	output Z6;
	output Z7;
	input  A;
	pmos _i0 (Z0, 1'b0, A);
	pmos _i1 (Z1, 1'b0, A);
	pmos _i2 (Z2, 1'b0, A);
	pmos _i3 (Z3, 1'b0, A);
	pmos _i4 (Z4, 1'b0, A);
	pmos _i5 (Z5, 1'b0, A);
	pmos _i6 (Z6, 1'b0, A);
	pmos _i7 (Z7, 1'b0, A);
	specify
	(A *> Z0) = (0,0,0,0,0,0);
	(A *> Z1) = (0,0,0,0,0,0);
	(A *> Z2) = (0,0,0,0,0,0);
	(A *> Z3) = (0,0,0,0,0,0);
	(A *> Z4) = (0,0,0,0,0,0);
	(A *> Z5) = (0,0,0,0,0,0);
	(A *> Z6) = (0,0,0,0,0,0);
	(A *> Z7) = (0,0,0,0,0,0);
	endspecify
endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2ODHDHT (Z, A, B);
	output Z;
	input  A;
	input  B;
	and _i0 (_n1,A,B);
	nmos _i1 (Z, 1'b0, _n1);
	specify
	(A *> Z) = (0,0,0,0,0,0);
	(B *> Z) = (0,0,0,0,0,0);
	endspecify
endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3ODHDHT (Z, A, B, C);
	output Z;
	input  A;
	input  B;
	input  C;
	and _i0 (_n1,C,A,B);
	nmos _i1 (Z, 1'b0, _n1);
	specify
	(A *> Z) = (0,0,0,0,0,0);
	(B *> Z) = (0,0,0,0,0,0);
	(C *> Z) = (0,0,0,0,0,0);
	endspecify
endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR2ODHDHT (Z, A, B);
	output Z;
	input  A;
	input  B;
	nor _i0 (_n1,A,B);
	nmos _i1 (Z, 1'b0, _n1);
	specify
	(A *> Z) = (0,0,0,0,0,0);
	(B *> Z) = (0,0,0,0,0,0);
	endspecify
endmodule
`endcelldefine

primitive p_mux21 (q, data1, data0, dselect);
    output q;
    input data1, data0, dselect;

// FUNCTION :  TWO TO ONE MULTIPLEXER
table
//data1 data0 dselect :   q
	0     0       ?   :   0 ;
	1     1       ?   :   1 ;

	0     ?       1   :   0 ;
	1     ?       1   :   1 ;

	?     0       0   :   0 ;
	?     1       0   :   1 ;
endtable
endprimitive

primitive ip_latchsr (Q, D, G, SB, RB, NOTIFIER);
   output Q;  
   input  D, G, SB, RB, NOTIFIER;
   reg    Q;

   table

// D  G  SB   RB  NOT  : Qt : Qt+1
//
   1  1   1   1   ?   : ?  :  1  ; // 
   0  1   1   1   ?   : ?  :  0  ; // 
   1  *   1   1   ?   : 1  :  1  ; // reduce pessimism
   0  *   1   1   ?   : 0  :  0  ; // reduce pessimism
   *  0   1   1   ?   : ?  :  -  ; // no changes when in switches
   ?  ?   0   ?   ?   : ?  :  1  ; // set output
   ?  0   (?1)   ?   ?   : 1  :  1  ; // cover all transistions on SB
   1  ?   (?1)   ?   ?   : 1  :  1  ; // cover all transistions on SB
   ?  ?   1   0   ?   : ?  :  0  ; // reset output
   ?  0   1   (?1)   ?   : 0  :  0  ; // cover all transistions on RB
   0  ?   1   (?1)   ?   : 0  :  0  ; // cover all transistions on RB
   ?  ?   ?   ?   *   : ?  :  x  ; // any notifier changed

   endtable
endprimitive // ip_latchsr


primitive ip_latchnsr (Q, D, GB, SB, RB, NOTIFIER);
   output Q;  
   input  D, GB, SB, RB, NOTIFIER;
   reg    Q;

   table

// D  GB  SB   RB  NOT  : Qt : Qt+1
//
   1  0   1   1   ?   : ?  :  1  ; //
   0  0   1   1   ?   : ?  :  0  ; //
   1  *   1   1   ?   : 1  :  1  ; // reduce pessimism
   0  *   1   1   ?   : 0  :  0  ; // reduce pessimism
   *  1   1   1   ?   : ?  :  -  ; // no changes when in switches
   ?  ?   0   ?   ?   : ?  :  1  ; // set output
   ?  1   (?1)   ?   ?   : 1  :  1  ; // cover all transistions on SB
   1  ?   (?1)   ?   ?   : 1  :  1  ; // cover all transistions on SB
   ?  ?   1   0   ?   : ?  :  0  ; // reset output
   ?  1   1   (?1)   ?   : 0  :  0  ; // cover all transistions on RB
   0  ?   1   (?1)   ?   : 0  :  0  ; // cover all transistions on RB
   ?  ?   ?   ?   *   : ?  :  x  ; // any notifier changed

   endtable
endprimitive // ip_latchnsr

primitive ip_ffsdsr (Q, D, CP, RB, SB, TE, TI, NOTIFIER);
    output Q;  reg    Q;
    input D, CP, RB, SB, TE, TI,NOTIFIER;
    table
    //  D   CP      RB   SB   TE   TI   No  :   Qt  :   Qt+1
        1 (01) 1 1 0 ? ? : ? : 1;  // clocked data 1
        ? (01) 1 1 1 1 ? : ? : 1;  // clocked scan in 1
        0 (01) 1 1 0 ? ? : ? : 0;  // clocked data 0
        ? (01) 1 1 1 0 ? : ? : 0;  // clocked scan in 0
        ? ? 0 1 ? ? ? : ? : 0;  // asynchronous clear
        ? ? ? 0 ? ? ? : ? : 1;  // asynchronous set
        ? (?0) ? ? ? ? ? : ? : -;  //ignore falling clock
        ? (1x) ? ? ? ? ? : ? : -;  //ignore falling clock
        * ? ? ? ? ? ? : ? : -;  // ignore data edges
        ? ? ? ? ? * ? : ? : -;  // ignore scan in edges
        ? ? ? ? * ? ? : ? : -;  // ignore scan enable edges
	1 (x1) 1 1 0 ? ? : 1 : 1;  // reducing pessimism
        ? (x1) 1 1 1 1 ? : 1 : 1;  // reducing pessimism
        0 (x1) 1 1 0 ? ? : 0 : 0;
        ? (x1) 1 1 1 0 ? : 0 : 0;
        1 (0x) 1 1 0 ? ? : 1 : 1;
        ? (0x) 1 1 1 1 ? : 1 : 1;
        0 (0x) 1 1 0 ? ? : 0 : 0;
        ? (0x) 1 1 1 0 ? : 0 : 0;
        ? ? (?1) 1 ? ? ? : ? : -;  // ignore the edges on
        ? ? ? (?1) ? ? ? : ? : -;  // set and clear

        ? ? ? ? ? ? * : ? : x;
    endtable
endprimitive

primitive ip_ffsdnsr (Q, D, CPB, RB, SB, TE, TI, NOTIFIER);
    output Q;  reg    Q;
    input D, CPB, RB, SB, TE, TI,NOTIFIER;
    table
    //  D   CPB    RB   SB   TE   TI   No  :   Qt  :   Qt+1
        1 (10) 1 1 0 ? ? : ? : 1;  // clocked data 1
        ? (10) 1 1 1 1 ? : ? : 1;  // clocked scan in 1
        0 (10) 1 1 0 ? ? : ? : 0;  // clocked data 0
        ? (10) 1 1 1 0 ? : ? : 0;  // clocked scan in 0
        ? ? 0 1 ? ? ? : ? : 0;  // asynchronous clear
        ? ? ? 0 ? ? ? : ? : 1;  // asynchronous set
        ? (?1) ? ? ? ? ? : ? : -;  //ignore rising clock
        ? (0x) ? ? ? ? ? : ? : -;  //ignore rising clock
        * ? ? ? ? ? ? : ? : -;  // ignore data edges
        ? ? ? ? ? * ? : ? : -;  // ignore scan in edges
        ? ? ? ? * ? ? : ? : -;  // ignore scan enable edges
	1 (x0) 1 1 0 ? ? : 1 : 1;  // reducing pessimism
        ? (x0) 1 1 1 1 ? : 1 : 1;  // reducing pessimism
        0 (x0) 1 1 0 ? ? : 0 : 0;
        ? (x0) 1 1 1 0 ? : 0 : 0;
        1 (1x) 1 1 0 ? ? : 1 : 1;
        ? (1x) 1 1 1 1 ? : 1 : 1;
        0 (1x) 1 1 0 ? ? : 0 : 0;
        ? (1x) 1 1 1 0 ? : 0 : 0;
        ? ? (?1) 1 ? ? ? : ? : -;  // ignore the edges on
        ? ? ? (?1) ? ? ? : ? : -;  // set and clear

        ? ? ? ? ? ? * : ? : x;
    endtable
endprimitive

primitive ip_ffsedcr (Q, D, CP, E, RB, TE, TI, NOTIFIER);
    output Q;  reg    Q;
    input D, CP, E, RB, TE, TI,NOTIFIER;
    table
    //  D   CP   E   RB   TE   TI   No  :   Qt  :   Qt+1
        1 (01) 1 1 0 ? ? : ? : 1;  // clocked data 1
        0 (01) 1 ? 0 ? ? : ? : 0;  // clocked data 0
	? (01) 0 ? 0 ? ? : 0 : 0;  // data disabled
	? (01) 0 1 0 ? ? : 1 : 1;  // data disabled
        ? (01) ? 0 0 ? ? : ? : 0;  // synchronous clear
        ? (01) ? ? 1 1 ? : ? : 1;  // clocked scan in 1
        ? (01) ? ? 1 0 ? : ? : 0;  // clocked scan in 0

        1 (x1) 1 1 0 ? ? : 1 : 1;  // reducing pessimism
        ? (x1) 0 1 0 ? ? : 1 : 1;  // reducing pessimism
        ? (x1) ? ? 1 1 ? : 1 : 1;
        0 (x1) 1 ? 0 ? ? : 0 : 0;
        ? (x1) 0 ? 0 ? ? : 0 : 0;
        ? (x1) ? 0 0 ? ? : 0 : 0;
        ? (x1) ? ? 1 0 ? : 0 : 0;
	1 (0x) 1 1 0 ? ? : 1 : 1;
	? (0x) 0 1 0 ? ? : 1 : 1;
	? (0x) ? ? 1 1 ? : 1 : 1;  
        0 (0x) 1 ? 0 ? ? : 0 : 0;
        ? (0x) 0 ? 0 ? ? : 0 : 0;
        ? (0x) ? 0 0 ? ? : 0 : 0;
        ? (0x) ? ? 1 0 ? : 0 : 0;

        ? (?0) ? ? ? ? ? : ? : -;  //ignore falling clock
        ? (1x) ? ? ? ? ? : ? : -;  //ignore falling clock
        * ? ? ? ? ? ? : ? : -;  // ignore data edges
        ? ? ? ? ? * ? : ? : -;  // ignore scan in edges
        ? ? ? ? * ? ? : ? : -;  // ignore scan enable edges
        ? ? * ? ? ? ? : ? : -;  // ignore enable edges
        ? ? ? * ? ? ? : ? : -;  // ignore clear edges

        ? ? ? ? ? ? * : ? : x;
    endtable
endprimitive

primitive ip_ffsjksr (Q, J, K, CP, RB, SB, TE, TI, NOTIFIER);
    output Q;  reg    Q;
    input J, K, CP, RB, SB, TE, TI,NOTIFIER;
    table
    //  J   K   CP   RB   SB   TE   TI   No  :   Qt  :   Qt+1
        1 0 (01) 1 1 0 ? ? : 0 : 1;  // clocked data 1
        1 0 (01) 1 1 0 ? ? : 1 : 1;  // clocked data 1
        0 1 (01) 1 1 0 ? ? : ? : 0;  // clocked data 0
        0 ? (01) 1 1 0 ? ? : 0 : 0;
        ? 0 (01) 1 1 0 ? ? : 1 : 1;
	1 ? (01) 1 1 0 ? ? : 0 : 1;  // J=1, K=1, toggle
	? 1 (01) 1 1 0 ? ? : 1 : 0;
        ? ? (01) 1 1 1 1 ? : ? : 1;  // clocked scan in 1
        ? ? (01) 1 1 1 0 ? : ? : 0;  // clocked scan in 0

        1 0 (x1) 1 1 0 ? ? : 1 : 1;  // reducing pessimism
        ? 0 (x1) 1 1 0 ? ? : 1 : 1;  // reducing pessimism
        ? ? (x1) 1 1 1 1 ? : 1 : 1;  // reducing pessimism
        0 1 (x1) 1 1 0 ? ? : 0 : 0;
        0 ? (x1) 1 1 0 ? ? : 0 : 0;
        ? ? (x1) 1 1 1 0 ? : 0 : 0;
        1 0 (0x) 1 1 0 ? ? : 1 : 1;
        ? 0 (0x) 1 1 0 ? ? : 1 : 1;
        ? ? (0x) 1 1 1 1 ? : 1 : 1;
        0 1 (0x) 1 1 0 ? ? : 0 : 0;
        0 ? (0x) 1 1 0 ? ? : 0 : 0;
        ? ? (0x) 1 1 1 0 ? : 0 : 0;

        ? ? ? 0 1 ? ? ? : ? : 0;  // asynchronous clear
        ? ? ? ? 0 ? ? ? : ? : 1;  // asynchronous set

        ? ? (?0) ? ? ? ? ? : ? : -;  //ignore falling clock
        ? ? (1x) ? ? ? ? ? : ? : -;  //ignore falling clock
        * ? ? ? ? ? ? ? : ? : -;  // ignore J edges
        ? * ? ? ? ? ? ? : ? : -;  // ignore K edges
        ? ? ? ? ? ? * ? : ? : -;  // ignore scan in edges
        ? ? ? ? ? * ? ? : ? : -;  // ignore scan enable edges

        ? ? ? (?1) 1 ? ? ? : ? : -;  // ignore the edges on
        ? ? ? ? (?1) ? ? ? : ? : -;  // set and clear

        ? ? ? ? ? ? ? * : ? : x;
    endtable
endprimitive

primitive rslat (Q, R, S, NOTIFIER);
    output Q;
    input  R, S, NOTIFIER;
    reg    Q;
    table
    //  R   S   NOT : Qt : Qt+1
        (?0) 0   ?   : ?  :  -  ; // no change
         0  (?0) ?   : ?  :  -  ; // no change
         1   ?   ?   : ?  :  0  ; // reset
        (?0) 1   ?   : ?  :  1  ; // set
         0  (?1) ?   : ?  :  1  ; // set
        (?0) x   ?   : 1  :  1  ; // reduced pessimism
         0  (?x) ?   : 1  :  1  ; // reduced pessimism
        (?x) 0   ?   : 0  :  0  ; // reduced pessimism
         x  (?0) ?   : 0  :  0  ; // reduced pessimism
         ?   ?   *   : ?  :  x  ; // any NOTIFIER changed
    endtable
endprimitive

primitive rslatn (QN, R, S, NOTIFIER);
    output QN;
    input  R, S, NOTIFIER;
    reg    QN;
    table
    //  R   S   NOT : Qt : Qt+1
        (?0) 0   ?   : ?  :  -  ; // no change
         0  (?0) ?   : ?  :  -  ; // no change
        (?1) 0   ?   : ?  :  1  ; // reset
         1  (?0) ?   : ?  :  1  ; // reset
         ?   1   ?   : ?  :  0  ; // set
        (?0) x   ?   : 0  :  0  ; // reduced pessimism
         0  (?x) ?   : 0  :  0  ; // reduced pessimism
        (?x) 0   ?   : 1  :  1  ; // reduced pessimism
         x  (?0) ?   : 1  :  1  ; // reduced pessimism
         ?   ?   *   : ?  :  x  ; // any NOTIFIER changed
    endtable
endprimitive

primitive rsblat (Q, RN, SN, NOTIFIER);
    output Q;
    input  RN, SN, NOTIFIER;
    reg    Q;
    table
    //  RN  SN  NOT : Qt : Qt+1
        (?1) 1   ?   : ?  :  -  ; // no change
         1  (?1) ?   : ?  :  -  ; // no change
        (?0) 1   ?   : ?  :  0  ; // reset
         0  (?1) ?   : ?  :  0  ; // reset
         ?   0   ?   : ?  :  1  ; // unused state
        (?1) x   ?   : 1  :  1  ; // reduced pessimism
         1  (?x) ?   : 1  :  1  ; // reduced pessimism
        (?x) 1   ?   : 0  :  0  ; // reduced pessimism
         x  (?1) ?   : 0  :  0  ; // reduced pessimism
         ?   ?   *   : ?  :  x  ; // any NOTIFIER changed
    endtable
endprimitive

primitive rsblatn (QN, RN, SN, NOTIFIER);
    output QN;
    input  RN, SN, NOTIFIER;
    reg    QN;
    table
    //  RN  SN  NOT : Qt : Qt+1
        (?1) 1   ?   : ?  :  -  ; // no change
         1  (?1) ?   : ?  :  -  ; // no change
         0   ?   ?   : ?  :  1  ; // reset
        (?1) 0   ?   : ?  :  0  ; // set
         1  (?0) ?   : ?  :  0  ; // set
        (?1) x   ?   : 0  :  0  ; // reduced pessimism
         1  (?x) ?   : 0  :  0  ; // reduced pessimism
        (?x) 1   ?   : 1  :  1  ; // reduced pessimism
         x  (?1) ?   : 1  :  1  ; // reduced pessimism
         ?   ?   *   : ?  :  x  ; // any NOTIFIER changed
    endtable
endprimitive

primitive udp_mux2 (out, in0, in1, sel);
   output out;
   input  in0, in1, sel;

   table

// sel in0 in1 :  out
//
    1  ?  0 :  1 ;
    0  ?  0 :  0 ;
    ?  1  1 :  1 ;
    ?  0  1 :  0 ;
    0  0  x :  0 ;
    1  1  x :  1 ;

   endtable
endprimitive // udp_mux2
