VERSION 5.3.1 ;

LAYER M1
    ANTENNACUMAREARATIO  600 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 600 ) ( 0.249 600 ) ( 0.251 2300.4 ) ( 1 2600 ) ) ;
END M1

LAYER V1
    ANTENNACUMAREARATIO  20 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.249 20 ) ( 0.25 92.59 ) ( 1 160 ) ) ;
END V1

LAYER M2
    ANTENNACUMAREARATIO  600 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 600 ) ( 0.249 600 ) ( 0.25 2300.4 ) ( 1 2600 ) ) ;
END M2

LAYER V2
    ANTENNACUMAREARATIO  20 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.249 20 ) ( 0.25 92.59 ) ( 1 160 ) ) ;
END V2

LAYER M3
    ANTENNACUMAREARATIO  600 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 600 ) ( 0.249 600 ) ( 0.25  2300.4 ) ( 1 2600 ) ) ;
END M3

LAYER V3
    ANTENNACUMAREARATIO  20 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.249 20 ) ( 0.25 92.59 ) ( 1 160 ) ) ;
END V3

LAYER M4
    ANTENNACUMAREARATIO  600 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 600 ) ( 0.249 600 ) ( 0.25  2300.4 ) ( 1 2600 ) ) ;
END M4

LAYER V4
    ANTENNACUMAREARATIO  20 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.249 20 ) ( 0.25 92.59 ) ( 1 160 ) ) ;
END V4

LAYER M5
    ANTENNACUMAREARATIO  600 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 600 ) ( 0.249 600 ) ( 0.25  2300.4 ) ( 1 2600 ) ) ;
END M5

LAYER V5
    ANTENNACUMAREARATIO  20 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.249 20 ) ( 0.25 92.59 ) ( 1 160 ) ) ;
END V5

LAYER M6
    ANTENNACUMAREARATIO  600 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 600 ) ( 0.249 600 ) ( 0.25  2300.4 ) ( 1 2600 ) ) ;
END M6

MACRO AND2CLKHD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.104 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.104 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5865 LAYER M1 ;
  END Z
END AND2CLKHD1X

MACRO AND2CLKHD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1664 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1664 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6747 LAYER M1 ;
  END Z
END AND2CLKHD2X

MACRO AND2CLKHD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.27155 LAYER M1 ;
  END Z
END AND2CLKHD3X

MACRO AND2CLKHD4X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2548 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2548 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.3494 LAYER M1 ;
  END Z
END AND2CLKHD4X

MACRO AND2HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END AND2HD1X

MACRO AND2HD1XSPG
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
    AntennaGateArea  0.0858 LAYER M2 ;
    AntennaGateArea  0.0858 LAYER M3 ;
    AntennaGateArea  0.0858 LAYER M4 ;
    AntennaGateArea  0.0858 LAYER M5 ;
    AntennaGateArea  0.0858 LAYER M6 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
    AntennaGateArea  0.0858 LAYER M2 ;
    AntennaGateArea  0.0858 LAYER M3 ;
    AntennaGateArea  0.0858 LAYER M4 ;
    AntennaGateArea  0.0858 LAYER M5 ;
    AntennaGateArea  0.0858 LAYER M6 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
    AntennaDiffArea  0.72795 LAYER M2 ;
    AntennaDiffArea  0.72795 LAYER M3 ;
    AntennaDiffArea  0.72795 LAYER M4 ;
    AntennaDiffArea  0.72795 LAYER M5 ;
    AntennaDiffArea  0.72795 LAYER M6 ;
  END Z
END AND2HD1XSPG

MACRO AND2HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1547 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1547 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END AND2HD2X

MACRO AND2HD2XSPG
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1547 LAYER M1 ;
    AntennaGateArea  0.1547 LAYER M2 ;
    AntennaGateArea  0.1547 LAYER M3 ;
    AntennaGateArea  0.1547 LAYER M4 ;
    AntennaGateArea  0.1547 LAYER M5 ;
    AntennaGateArea  0.1547 LAYER M6 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1547 LAYER M1 ;
    AntennaGateArea  0.1547 LAYER M2 ;
    AntennaGateArea  0.1547 LAYER M3 ;
    AntennaGateArea  0.1547 LAYER M4 ;
    AntennaGateArea  0.1547 LAYER M5 ;
    AntennaGateArea  0.1547 LAYER M6 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
    AntennaDiffArea  0.8229 LAYER M2 ;
    AntennaDiffArea  0.8229 LAYER M3 ;
    AntennaDiffArea  0.8229 LAYER M4 ;
    AntennaDiffArea  0.8229 LAYER M5 ;
    AntennaDiffArea  0.8229 LAYER M6 ;
  END Z
END AND2HD2XSPG

MACRO AND2HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
END AND2HDLX

MACRO AND2HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END AND2HDMX

MACRO AND2HDUX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.216 LAYER M1 ;
  END Z
END AND2HDUX

MACRO AND3HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0884 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0884 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0884 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END AND3HD1X

MACRO AND3HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8651 LAYER M1 ;
  END Z
END AND3HD2X

MACRO AND3HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
END AND3HDLX

MACRO AND3HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END AND3HDMX

MACRO AND4HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.091 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.091 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.091 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.091 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.74905 LAYER M1 ;
  END Z
END AND4HD1X

MACRO AND4HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1859 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1859 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1859 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1859 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8651 LAYER M1 ;
  END Z
END AND4HD2X

MACRO AND4HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2556 LAYER M1 ;
  END Z
END AND4HDLX

MACRO AND4HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3834 LAYER M1 ;
  END Z
END AND4HDMX

MACRO ANTFIXHD
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.7744 LAYER M1 ;
  END Z
END ANTFIXHD

MACRO AOI211HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END AOI211HD1X

MACRO AOI211HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END AOI211HD2X

MACRO AOI211HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.66735 LAYER M1 ;
  END Z
END AOI211HDLX

MACRO AOI211HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END AOI211HDMX

MACRO AOI21B2HD1X
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
  END C
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.67715 LAYER M1 ;
  END Z
END AOI21B2HD1X

MACRO AOI21B2HD2X
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1209 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.4862 LAYER M1 ;
  END C
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1209 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.9949 LAYER M1 ;
  END Z
END AOI21B2HD2X

MACRO AOI21B2HDLX
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END C
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.31365 LAYER M1 ;
  END Z
END AOI21B2HDLX

MACRO AOI21B2HDMX
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1703 LAYER M1 ;
  END C
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4722 LAYER M1 ;
  END Z
END AOI21B2HDMX

MACRO AOI21HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8328 LAYER M1 ;
  END Z
END AOI21HD1X

MACRO AOI21HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END AOI21HD2X

MACRO AOI21HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.34755 LAYER M1 ;
  END Z
END AOI21HDLX

MACRO AOI21HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1885 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1885 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1703 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5163 LAYER M1 ;
  END Z
END AOI21HDMX

MACRO AOI21HDUX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0754 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2569 LAYER M1 ;
  END Z
END AOI21HDUX

MACRO AOI221HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END AOI221HD1X

MACRO AOI221HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END AOI221HD2X

MACRO AOI221HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8514 LAYER M1 ;
  END Z
END AOI221HDLX

MACRO AOI221HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3861 LAYER M1 ;
  END Z
END AOI221HDMX

MACRO AOI222HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END AOI222HD1X

MACRO AOI222HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END AOI222HD2X

MACRO AOI222HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.693 LAYER M1 ;
  END Z
END AOI222HDLX

MACRO AOI222HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3915 LAYER M1 ;
  END Z
END AOI222HDMX

MACRO AOI22B2HD1X
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.73395 LAYER M1 ;
  END Z
END AOI22B2HD1X

MACRO AOI22B2HD2X
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1209 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1209 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.0725 LAYER M1 ;
  END Z
END AOI22B2HD2X

MACRO AOI22B2HDLX
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3105 LAYER M1 ;
  END Z
END AOI22B2HDLX

MACRO AOI22B2HDMX
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1885 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1885 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.454 LAYER M1 ;
  END Z
END AOI22B2HDMX

MACRO AOI22HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.99265 LAYER M1 ;
  END Z
END AOI22HD1X

MACRO AOI22HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END AOI22HD2X

MACRO AOI22HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.303 LAYER M1 ;
  END Z
END AOI22HDLX

MACRO AOI22HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.44475 LAYER M1 ;
  END Z
END AOI22HDMX

MACRO AOI22HDUX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2772 LAYER M1 ;
  END Z
END AOI22HDUX

MACRO AOI31HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.221 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8412 LAYER M1 ;
  END Z
END AOI31HD1X

MACRO AOI31HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1404 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END AOI31HD2X

MACRO AOI31HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1404 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.47585 LAYER M1 ;
  END Z
END AOI31HDLX

MACRO AOI31HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2119 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2119 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2119 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6502 LAYER M1 ;
  END Z
END AOI31HDMX

MACRO AOI32HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2392 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2392 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8187 LAYER M1 ;
  END Z
END AOI32HD1X

MACRO AOI32HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1326 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1326 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1326 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END AOI32HD2X

MACRO AOI32HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1326 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1326 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1326 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4008 LAYER M1 ;
  END Z
END AOI32HDLX

MACRO AOI32HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1807 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1807 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1807 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1599 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1599 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5472 LAYER M1 ;
  END Z
END AOI32HDMX

MACRO AOI33HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.26105 LAYER M1 ;
  END Z
END AOI33HD1X

MACRO AOI33HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END AOI33HD2X

MACRO AOI33HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.44205 LAYER M1 ;
  END Z
END AOI33HDLX

MACRO AOI33HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.69825 LAYER M1 ;
  END Z
END AOI33HDMX

MACRO BUFCLKHD10X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.689 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.1041 LAYER M1 ;
  END Z
END BUFCLKHD10X

MACRO BUFCLKHD12X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.689 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.90525 LAYER M1 ;
  END Z
END BUFCLKHD12X

MACRO BUFCLKHD14X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.9217 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.6075 LAYER M1 ;
  END Z
END BUFCLKHD14X

MACRO BUFCLKHD16X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.157 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  4.3139 LAYER M1 ;
  END Z
END BUFCLKHD16X

MACRO BUFCLKHD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5934 LAYER M1 ;
  END Z
END BUFCLKHD1X

MACRO BUFCLKHD20X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.521 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  7.3671 LAYER M1 ;
  END Z
END BUFCLKHD20X

MACRO BUFCLKHD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.7045 LAYER M1 ;
  END Z
END BUFCLKHD2X

MACRO BUFCLKHD30X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.6796 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  10.7733 LAYER M1 ;
  END Z
END BUFCLKHD30X

MACRO BUFCLKHD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.35835 LAYER M1 ;
  END Z
END BUFCLKHD3X

MACRO BUFCLKHD40X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  2.236 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  13.962 LAYER M1 ;
  END Z
END BUFCLKHD40X

MACRO BUFCLKHD4X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2236 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.43775 LAYER M1 ;
  END Z
END BUFCLKHD4X

MACRO BUFCLKHD5X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2236 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.0355 LAYER M1 ;
  END Z
END BUFCLKHD5X

MACRO BUFCLKHD6X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.3367 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.78875 LAYER M1 ;
  END Z
END BUFCLKHD6X

MACRO BUFCLKHD7X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.3367 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.1996 LAYER M1 ;
  END Z
END BUFCLKHD7X

MACRO BUFCLKHD80X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  4.5916 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  27.9403 LAYER M1 ;
  END Z
END BUFCLKHD80X

MACRO BUFCLKHD8X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4628 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.0508 LAYER M1 ;
  END Z
END BUFCLKHD8X

MACRO BUFCLKHDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.36225 LAYER M1 ;
  END Z
END BUFCLKHDLX

MACRO BUFCLKHDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4347 LAYER M1 ;
  END Z
END BUFCLKHDMX

MACRO BUFCLKHDUX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.091 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2775 LAYER M1 ;
  END Z
END BUFCLKHDUX

MACRO BUFHD12X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.0972 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  4.9374 LAYER M1 ;
  END Z
END BUFHD12X

MACRO BUFHD16X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.3715 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  6.5832 LAYER M1 ;
  END Z
END BUFHD16X

MACRO BUFHD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END BUFHD1X

MACRO BUFHD20X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.6458 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  8.229 LAYER M1 ;
  END Z
END BUFHD20X

MACRO BUFHD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1846 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END BUFHD2X

MACRO BUFHD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END BUFHD3X

MACRO BUFHD4X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.3653 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.6458 LAYER M1 ;
  END Z
END BUFHD4X

MACRO BUFHD5X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.3653 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.37375 LAYER M1 ;
  END Z
END BUFHD5X

MACRO BUFHD6X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4121 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.4687 LAYER M1 ;
  END Z
END BUFHD6X

MACRO BUFHD7X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.19665 LAYER M1 ;
  END Z
END BUFHD7X

MACRO BUFHD8X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.7306 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.2916 LAYER M1 ;
  END Z
END BUFHD8X

MACRO BUFHD8XSPG
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.7306 LAYER M1 ;
    AntennaGateArea  0.7306 LAYER M2 ;
    AntennaGateArea  0.7306 LAYER M3 ;
    AntennaGateArea  0.7306 LAYER M4 ;
    AntennaGateArea  0.7306 LAYER M5 ;
    AntennaGateArea  0.7306 LAYER M6 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.2916 LAYER M1 ;
    AntennaDiffArea  3.2916 LAYER M2 ;
    AntennaDiffArea  3.2916 LAYER M3 ;
    AntennaDiffArea  3.2916 LAYER M4 ;
    AntennaDiffArea  3.2916 LAYER M5 ;
    AntennaDiffArea  3.2916 LAYER M6 ;
  END Z
END BUFHD8XSPG

MACRO BUFHDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
END BUFHDLX

MACRO BUFHDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END BUFHDMX

MACRO BUFHDUX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0624 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.216 LAYER M1 ;
  END Z
END BUFHDUX

MACRO BUFTSHD12X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.8229 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.6578 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  5.5704 LAYER M1 ;
  END Z
END BUFTSHD12X

MACRO BUFTSHD16X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.6458 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  1.0335 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  7.2162 LAYER M1 ;
  END Z
END BUFTSHD16X

MACRO BUFTSHD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2613 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6694 LAYER M1 ;
  END Z
END BUFTSHD1X

MACRO BUFTSHD20X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.9201 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  1.209 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  8.862 LAYER M1 ;
  END Z
END BUFTSHD20X

MACRO BUFTSHD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1924 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.034 LAYER M1 ;
  END Z
END BUFTSHD2X

MACRO BUFTSHD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.2349 LAYER M1 ;
  END Z
END BUFTSHD3X

MACRO BUFTSHD4X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4368 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.299 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.89385 LAYER M1 ;
  END Z
END BUFTSHD4X

MACRO BUFTSHD5X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4992 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.3432 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.37375 LAYER M1 ;
  END Z
END BUFTSHD5X

MACRO BUFTSHD6X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.3705 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.4687 LAYER M1 ;
  END Z
END BUFTSHD6X

MACRO BUFTSHD7X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.7488 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.442 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.19665 LAYER M1 ;
  END Z
END BUFTSHD7X

MACRO BUFTSHD8X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.8229 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.4186 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.9246 LAYER M1 ;
  END Z
END BUFTSHD8X

MACRO BUFTSHDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1443 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.40365 LAYER M1 ;
  END Z
END BUFTSHDLX

MACRO BUFTSHDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1703 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6072 LAYER M1 ;
  END Z
END BUFTSHDMX

MACRO BUFTSHDUX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0624 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.0884 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2275 LAYER M1 ;
  END Z
END BUFTSHDUX

MACRO DEL1HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.7042 LAYER M1 ;
  END Z
END DEL1HD1X

MACRO DEL1HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END DEL1HDMX

MACRO DEL1HDMXSPG
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
    AntennaGateArea  0.0936 LAYER M2 ;
    AntennaGateArea  0.0936 LAYER M3 ;
    AntennaGateArea  0.0936 LAYER M4 ;
    AntennaGateArea  0.0936 LAYER M5 ;
    AntennaGateArea  0.0936 LAYER M6 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.35835 LAYER M1 ;
    AntennaDiffArea  0.35835 LAYER M2 ;
    AntennaDiffArea  0.35835 LAYER M3 ;
    AntennaDiffArea  0.35835 LAYER M4 ;
    AntennaDiffArea  0.35835 LAYER M5 ;
    AntennaDiffArea  0.35835 LAYER M6 ;
  END Z
END DEL1HDMXSPG

MACRO DEL2HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END DEL2HD1X

MACRO DEL2HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END DEL2HDMX

MACRO DEL2HDMXSPG
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
    AntennaGateArea  0.0936 LAYER M2 ;
    AntennaGateArea  0.0936 LAYER M3 ;
    AntennaGateArea  0.0936 LAYER M4 ;
    AntennaGateArea  0.0936 LAYER M5 ;
    AntennaGateArea  0.0936 LAYER M6 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
    AntennaDiffArea  0.327 LAYER M2 ;
    AntennaDiffArea  0.327 LAYER M3 ;
    AntennaDiffArea  0.327 LAYER M4 ;
    AntennaDiffArea  0.327 LAYER M5 ;
    AntennaDiffArea  0.327 LAYER M6 ;
  END Z
END DEL2HDMXSPG

MACRO DEL3HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END DEL3HD1X

MACRO DEL3HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END DEL3HDMX

MACRO DEL4HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END DEL4HD1X

MACRO DEL4HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END DEL4HDMX

MACRO DEL4HDMXSPG
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
    AntennaGateArea  0.0936 LAYER M2 ;
    AntennaGateArea  0.0936 LAYER M3 ;
    AntennaGateArea  0.0936 LAYER M4 ;
    AntennaGateArea  0.0936 LAYER M5 ;
    AntennaGateArea  0.0936 LAYER M6 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
    AntennaDiffArea  0.327 LAYER M2 ;
    AntennaDiffArea  0.327 LAYER M3 ;
    AntennaDiffArea  0.327 LAYER M4 ;
    AntennaDiffArea  0.327 LAYER M5 ;
    AntennaDiffArea  0.327 LAYER M6 ;
  END Z
END DEL4HDMXSPG

MACRO FAHD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4368 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.3211 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END S
  PIN CI
    #DIRECTION INPUT ;
    AntennaGateArea  0.2886 LAYER M1 ;
  END CI
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5845 LAYER M1 ;
  END CO
END FAHD1X

MACRO FAHD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.4823 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END S
  PIN CI
    #DIRECTION INPUT ;
    AntennaGateArea  0.3939 LAYER M1 ;
  END CI
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END CO
END FAHD2X

MACRO FAHDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.3744 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.3211 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END S
  PIN CI
    #DIRECTION INPUT ;
    AntennaGateArea  0.2626 LAYER M1 ;
  END CI
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.261 LAYER M1 ;
  END CO
END FAHDLX

MACRO FAHDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.3744 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.3211 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.36225 LAYER M1 ;
  END S
  PIN CI
    #DIRECTION INPUT ;
    AntennaGateArea  0.2626 LAYER M1 ;
  END CI
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.38115 LAYER M1 ;
  END CO
END FAHDMX

MACRO FAHDUX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.216 LAYER M1 ;
  END S
  PIN CI
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END CI
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.216 LAYER M1 ;
  END CO
END FAHDUX

MACRO FAHHD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END S
  PIN CI
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END CI
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.73985 LAYER M1 ;
  END CO
END FAHHD1X

MACRO FAHHD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1651 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.3029 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END S
  PIN CI
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END CI
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END CO
END FAHHD2X

MACRO FAHHDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2499 LAYER M1 ;
  END S
  PIN CI
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END CI
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.255 LAYER M1 ;
  END CO
END FAHHDLX

MACRO FAHHDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3741 LAYER M1 ;
  END S
  PIN CI
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END CI
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3855 LAYER M1 ;
  END CO
END FAHHDMX

MACRO FFDCRHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
END FFDCRHD1X

MACRO FFDCRHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1144 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1144 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
END FFDCRHD2X

MACRO FFDCRHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.24 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.052 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.052 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
END FFDCRHDLX

MACRO FFDCRHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.33 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0637 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0637 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
END FFDCRHDMX

MACRO FFDHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
END FFDHD1X

MACRO FFDHD1XSPG
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
    AntennaDiffArea  0.72795 LAYER M2 ;
    AntennaDiffArea  0.72795 LAYER M3 ;
    AntennaDiffArea  0.72795 LAYER M4 ;
    AntennaDiffArea  0.72795 LAYER M5 ;
    AntennaDiffArea  0.72795 LAYER M6 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
    AntennaDiffArea  0.72795 LAYER M2 ;
    AntennaDiffArea  0.72795 LAYER M3 ;
    AntennaDiffArea  0.72795 LAYER M4 ;
    AntennaDiffArea  0.72795 LAYER M5 ;
    AntennaDiffArea  0.72795 LAYER M6 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
    AntennaGateArea  0.117 LAYER M2 ;
    AntennaGateArea  0.117 LAYER M3 ;
    AntennaGateArea  0.117 LAYER M4 ;
    AntennaGateArea  0.117 LAYER M5 ;
    AntennaGateArea  0.117 LAYER M6 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
    AntennaGateArea  0.078 LAYER M2 ;
    AntennaGateArea  0.078 LAYER M3 ;
    AntennaGateArea  0.078 LAYER M4 ;
    AntennaGateArea  0.078 LAYER M5 ;
    AntennaGateArea  0.078 LAYER M6 ;
  END CK
END FFDHD1XSPG

MACRO FFDHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
END FFDHD2X

MACRO FFDHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
END FFDHDLX

MACRO FFDHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
END FFDHDMX

MACRO FFDHQHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
END FFDHQHD1X

MACRO FFDHQHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
END FFDHQHD2X

MACRO FFDHQHD3X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
END FFDHQHD3X

MACRO FFDHQHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
END FFDHQHDMX

MACRO FFDNHD1X
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
END FFDNHD1X

MACRO FFDNHD2X
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
END FFDNHD2X

MACRO FFDNHDLX
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.065 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
END FFDNHDLX

MACRO FFDNHDMX
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
END FFDNHDMX

MACRO FFDNRHD1X
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
END FFDNRHD1X

MACRO FFDNRHD2X
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
END FFDNRHD2X

MACRO FFDNRHDLX
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.065 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
END FFDNRHDLX

MACRO FFDNRHDMX
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
END FFDNRHDMX

MACRO FFDNSHD1X
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFDNSHD1X

MACRO FFDNSHD2X
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3094 LAYER M1 ;
  END SN
END FFDNSHD2X

MACRO FFDNSHDLX
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.065 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFDNSHDLX

MACRO FFDNSHDMX
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFDNSHDMX

MACRO FFDNSRHD1X
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6814 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6168 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFDNSRHD1X

MACRO FFDNSRHD2X
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.338 LAYER M1 ;
  END SN
END FFDNSRHD2X

MACRO FFDNSRHDLX
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.065 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFDNSRHDLX

MACRO FFDNSRHDMX
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFDNSRHDMX

MACRO FFDQHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
END FFDQHD1X

MACRO FFDQHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
END FFDQHD2X

MACRO FFDQHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.27255 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
END FFDQHDLX

MACRO FFDQHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
END FFDQHDMX

MACRO FFDQRHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
END FFDQRHD1X

MACRO FFDQRHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
END FFDQRHD2X

MACRO FFDQRHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
END FFDQRHDLX

MACRO FFDQRHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
END FFDQRHDMX

MACRO FFDQSHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1859 LAYER M1 ;
  END SN
END FFDQSHD1X

MACRO FFDQSHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2405 LAYER M1 ;
  END SN
END FFDQSHD2X

MACRO FFDQSHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFDQSHDLX

MACRO FFDQSHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFDQSHDMX

MACRO FFDQSRHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1859 LAYER M1 ;
  END SN
END FFDQSRHD1X

MACRO FFDQSRHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2405 LAYER M1 ;
  END SN
END FFDQSRHD2X

MACRO FFDQSRHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFDQSRHDLX

MACRO FFDQSRHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFDQSRHDMX

MACRO FFDRHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
END FFDRHD1X

MACRO FFDRHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
END FFDRHD2X

MACRO FFDRHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
END FFDRHDLX

MACRO FFDRHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
END FFDRHDMX

MACRO FFDRHQHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
END FFDRHQHD1X

MACRO FFDRHQHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1755 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1404 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
END FFDRHQHD2X

MACRO FFDRHQHD3X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.5043 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2145 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
END FFDRHQHD3X

MACRO FFDRHQHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
END FFDRHQHDMX

MACRO FFDSHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFDSHD1X

MACRO FFDSHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3094 LAYER M1 ;
  END SN
END FFDSHD2X

MACRO FFDSHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFDSHDLX

MACRO FFDSHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFDSHDMX

MACRO FFDSHQHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2574 LAYER M1 ;
  END SN
END FFDSHQHD1X

MACRO FFDSHQHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.4559 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1755 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3198 LAYER M1 ;
  END SN
END FFDSHQHD2X

MACRO FFDSHQHD3X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2145 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3783 LAYER M1 ;
  END SN
END FFDSHQHD3X

MACRO FFDSHQHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFDSHQHDMX

MACRO FFDSRHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.70515 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.70515 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFDSRHD1X

MACRO FFDSRHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.338 LAYER M1 ;
  END SN
END FFDSRHD2X

MACRO FFDSRHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFDSRHDLX

MACRO FFDSRHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.35835 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.35835 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFDSRHDMX

MACRO FFDSRHQHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
  END SN
END FFDSRHQHD1X

MACRO FFDSRHQHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1755 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1404 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3198 LAYER M1 ;
  END SN
END FFDSRHQHD2X

MACRO FFDSRHQHD3X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2145 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3783 LAYER M1 ;
  END SN
END FFDSRHQHD3X

MACRO FFDSRHQHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3945 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.208 LAYER M1 ;
  END SN
END FFDSRHQHDMX

MACRO FFEDCRHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
END FFEDCRHD1X

MACRO FFEDCRHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
END FFEDCRHD2X

MACRO FFEDCRHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END E
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
END FFEDCRHDLX

MACRO FFEDCRHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3945 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1794 LAYER M1 ;
  END E
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
END FFEDCRHDMX

MACRO FFEDHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.7042 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
END FFEDHD1X

MACRO FFEDHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.2659 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
END FFEDHD2X

MACRO FFEDHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1794 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
END FFEDHDLX

MACRO FFEDHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
END FFEDHDMX

MACRO FFEDHQHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
END FFEDHQHD1X

MACRO FFEDHQHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.234 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.3276 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
END FFEDHQHD2X

MACRO FFEDHQHD3X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2756 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.3692 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
END FFEDHQHD3X

MACRO FFEDHQHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.52095 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
END FFEDHQHDMX

MACRO FFEDQHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
END FFEDQHD1X

MACRO FFEDQHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
END FFEDQHD2X

MACRO FFEDQHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
END FFEDQHDLX

MACRO FFEDQHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1794 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
END FFEDQHDMX

MACRO FFSDCRHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSDCRHD1X

MACRO FFSDCRHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSDCRHD2X

MACRO FFSDCRHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.169 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0689 LAYER M1 ;
  END TI
END FFSDCRHDLX

MACRO FFSDCRHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1144 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1144 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1846 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0689 LAYER M1 ;
  END TI
END FFSDCRHDMX

MACRO FFSDHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDHD1X

MACRO FFSDHD1XSPG
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
    AntennaDiffArea  0.72795 LAYER M2 ;
    AntennaDiffArea  0.72795 LAYER M3 ;
    AntennaDiffArea  0.72795 LAYER M4 ;
    AntennaDiffArea  0.72795 LAYER M5 ;
    AntennaDiffArea  0.72795 LAYER M6 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
    AntennaDiffArea  0.72795 LAYER M2 ;
    AntennaDiffArea  0.72795 LAYER M3 ;
    AntennaDiffArea  0.72795 LAYER M4 ;
    AntennaDiffArea  0.72795 LAYER M5 ;
    AntennaDiffArea  0.72795 LAYER M6 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
    AntennaGateArea  0.156 LAYER M2 ;
    AntennaGateArea  0.156 LAYER M3 ;
    AntennaGateArea  0.156 LAYER M4 ;
    AntennaGateArea  0.156 LAYER M5 ;
    AntennaGateArea  0.156 LAYER M6 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
    AntennaGateArea  0.2366 LAYER M2 ;
    AntennaGateArea  0.2366 LAYER M3 ;
    AntennaGateArea  0.2366 LAYER M4 ;
    AntennaGateArea  0.2366 LAYER M5 ;
    AntennaGateArea  0.2366 LAYER M6 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
    AntennaGateArea  0.078 LAYER M2 ;
    AntennaGateArea  0.078 LAYER M3 ;
    AntennaGateArea  0.078 LAYER M4 ;
    AntennaGateArea  0.078 LAYER M5 ;
    AntennaGateArea  0.078 LAYER M6 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
    AntennaGateArea  0.117 LAYER M2 ;
    AntennaGateArea  0.117 LAYER M3 ;
    AntennaGateArea  0.117 LAYER M4 ;
    AntennaGateArea  0.117 LAYER M5 ;
    AntennaGateArea  0.117 LAYER M6 ;
  END TI
END FFSDHD1XSPG

MACRO FFSDHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDHD2X

MACRO FFSDHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
END FFSDHDLX

MACRO FFSDHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
END FFSDHDMX

MACRO FFSDHQHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDHQHD1X

MACRO FFSDHQHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.234 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2886 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDHQHD2X

MACRO FFSDHQHD3X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2925 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDHQHD3X

MACRO FFSDHQHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4752 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDHQHDMX

MACRO FFSDNHD1X
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDNHD1X

MACRO FFSDNHD2X
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDNHD2X

MACRO FFSDNHDLX
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.065 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
END FFSDNHDLX

MACRO FFSDNHDMX
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
END FFSDNHDMX

MACRO FFSDNRHD1X
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.70515 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDNRHD1X

MACRO FFSDNRHD2X
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDNRHD2X

MACRO FFSDNRHDLX
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.065 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
END FFSDNRHDLX

MACRO FFSDNRHDMX
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
END FFSDNRHDMX

MACRO FFSDNSHD1X
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFSDNSHD1X

MACRO FFSDNSHD2X
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3094 LAYER M1 ;
  END SN
END FFSDNSHD2X

MACRO FFSDNSHDLX
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.065 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFSDNSHDLX

MACRO FFSDNSHDMX
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFSDNSHDMX

MACRO FFSDNSRHD1X
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6814 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6168 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFSDNSRHD1X

MACRO FFSDNSRHD2X
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.338 LAYER M1 ;
  END SN
END FFSDNSRHD2X

MACRO FFSDNSRHDLX
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.065 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFSDNSRHDLX

MACRO FFSDNSRHDMX
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFSDNSRHDMX

MACRO FFSDQHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDQHD1X

MACRO FFSDQHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDQHD2X

MACRO FFSDQHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
END FFSDQHDLX

MACRO FFSDQHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
END FFSDQHDMX

MACRO FFSDQRHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDQRHD1X

MACRO FFSDQRHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDQRHD2X

MACRO FFSDQRHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
END FFSDQRHDLX

MACRO FFSDQRHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
END FFSDQRHDMX

MACRO FFSDQSHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1859 LAYER M1 ;
  END SN
END FFSDQSHD1X

MACRO FFSDQSHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2405 LAYER M1 ;
  END SN
END FFSDQSHD2X

MACRO FFSDQSHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2709 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFSDQSHDLX

MACRO FFSDQSHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFSDQSHDMX

MACRO FFSDQSRHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1859 LAYER M1 ;
  END SN
END FFSDQSRHD1X

MACRO FFSDQSRHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2405 LAYER M1 ;
  END SN
END FFSDQSRHD2X

MACRO FFSDQSRHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFSDQSRHDLX

MACRO FFSDQSRHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFSDQSRHDMX

MACRO FFSDRHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDRHD1X

MACRO FFSDRHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDRHD2X

MACRO FFSDRHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
END FFSDRHDLX

MACRO FFSDRHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
END FFSDRHDMX

MACRO FFSDRHQHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDRHQHD1X

MACRO FFSDRHQHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.234 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1404 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2886 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDRHQHD2X

MACRO FFSDRHQHD3X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2925 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDRHQHD3X

MACRO FFSDRHQHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDRHQHDMX

MACRO FFSDSHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFSDSHD1X

MACRO FFSDSHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3094 LAYER M1 ;
  END SN
END FFSDSHD2X

MACRO FFSDSHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFSDSHDLX

MACRO FFSDSHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFSDSHDMX

MACRO FFSDSHQHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2574 LAYER M1 ;
  END SN
END FFSDSHQHD1X

MACRO FFSDSHQHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.234 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2886 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3198 LAYER M1 ;
  END SN
END FFSDSHQHD2X

MACRO FFSDSHQHD3X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2925 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3783 LAYER M1 ;
  END SN
END FFSDSHQHD3X

MACRO FFSDSHQHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFSDSHQHDMX

MACRO FFSDSRHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.70515 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.70515 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFSDSRHD1X

MACRO FFSDSRHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.338 LAYER M1 ;
  END SN
END FFSDSRHD2X

MACRO FFSDSRHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFSDSRHDLX

MACRO FFSDSRHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFSDSRHDMX

MACRO FFSDSRHQHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
  END SN
END FFSDSRHQHD1X

MACRO FFSDSRHQHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.234 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1404 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2886 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3198 LAYER M1 ;
  END SN
END FFSDSRHQHD2X

MACRO FFSDSRHQHD3X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.49955 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2925 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3783 LAYER M1 ;
  END SN
END FFSDSRHQHD3X

MACRO FFSDSRHQHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.208 LAYER M1 ;
  END SN
END FFSDSRHQHDMX

MACRO FFSEDCRHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSEDCRHD1X

MACRO FFSEDCRHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSEDCRHD2X

MACRO FFSEDCRHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END E
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
END FFSEDCRHDLX

MACRO FFSEDCRHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1794 LAYER M1 ;
  END E
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
END FFSEDCRHDMX

MACRO FFSEDHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDHD1X

MACRO FFSEDHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDHD2X

MACRO FFSEDHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDHDLX

MACRO FFSEDHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.35835 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.35835 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1794 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDHDMX

MACRO FFSEDHQHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDHQHD1X

MACRO FFSEDHQHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDHQHD2X

MACRO FFSEDHQHD3X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDHQHD3X

MACRO FFSEDHQHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.52095 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDHQHDMX

MACRO FFSEDQHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDQHD1X

MACRO FFSEDQHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDQHD2X

MACRO FFSEDQHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDQHDLX

MACRO FFSEDQHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1794 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDQHDMX

MACRO FILLER16HD
END FILLER16HD

MACRO FILLER1HD
END FILLER1HD

MACRO FILLER2HD
END FILLER2HD

MACRO FILLER32HD
END FILLER32HD

MACRO FILLER3HD
END FILLER3HD

MACRO FILLER4HD
END FILLER4HD

MACRO FILLER64HD
END FILLER64HD

MACRO FILLER6HD
END FILLER6HD

MACRO FILLER8HD
END FILLER8HD

MACRO FILLERC16HD
END FILLERC16HD

MACRO FILLERC1HD
END FILLERC1HD

MACRO FILLERC2HD
END FILLERC2HD

MACRO FILLERC32HD
END FILLERC32HD

MACRO FILLERC3HD
END FILLERC3HD

MACRO FILLERC4HD
END FILLERC4HD

MACRO FILLERC64HD
END FILLERC64HD

MACRO FILLERC6HD
END FILLERC6HD

MACRO FILLERC8HD
END FILLERC8HD

MACRO HAHD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1885 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END S
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END CO
END HAHD1X

MACRO HAHD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.3276 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.4108 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END S
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END CO
END HAHD2X

MACRO HAHDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1794 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2574 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END S
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END CO
END HAHDLX

MACRO HAHDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1794 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2574 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END S
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END CO
END HAHDMX

MACRO HOLDHD
  PIN Z
    #DIRECTION INOUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
    AntennaDiffArea  0.32445 LAYER M1 ;
  END Z
END HOLDHD

MACRO INVCLKHD10X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.911 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.09885 LAYER M1 ;
  END Z
END INVCLKHD10X

MACRO INVCLKHD12X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  2.262 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.393 LAYER M1 ;
  END Z
END INVCLKHD12X

MACRO INVCLKHD14X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  2.7807 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  4.3834 LAYER M1 ;
  END Z
END INVCLKHD14X

MACRO INVCLKHD16X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  3.484 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  5.2326 LAYER M1 ;
  END Z
END INVCLKHD16X

MACRO INVCLKHD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2236 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5934 LAYER M1 ;
  END Z
END INVCLKHD1X

MACRO INVCLKHD20X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  4.537 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  6.8066 LAYER M1 ;
  END Z
END INVCLKHD20X

MACRO INVCLKHD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4498 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6747 LAYER M1 ;
  END Z
END INVCLKHD2X

MACRO INVCLKHD30X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.455 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  10.3545 LAYER M1 ;
  END Z
END INVCLKHD30X

MACRO INVCLKHD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.6838 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.2897 LAYER M1 ;
  END Z
END INVCLKHD3X

MACRO INVCLKHD40X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5642 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  14.0082 LAYER M1 ;
  END Z
END INVCLKHD40X

MACRO INVCLKHD4X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.9087 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.3636 LAYER M1 ;
  END Z
END INVCLKHD4X

MACRO INVCLKHD5X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.053 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.8225 LAYER M1 ;
  END Z
END INVCLKHD5X

MACRO INVCLKHD6X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.2324 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.8486 LAYER M1 ;
  END Z
END INVCLKHD6X

MACRO INVCLKHD7X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.417 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.2324 LAYER M1 ;
  END Z
END INVCLKHD7X

MACRO INVCLKHD80X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.1193 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  28.0111 LAYER M1 ;
  END Z
END INVCLKHD80X

MACRO INVCLKHD8X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.638 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.4659 LAYER M1 ;
  END Z
END INVCLKHD8X

MACRO INVCLKHDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.36225 LAYER M1 ;
  END Z
END INVCLKHDLX

MACRO INVCLKHDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4347 LAYER M1 ;
  END Z
END INVCLKHDMX

MACRO INVCLKHDUX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.091 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2775 LAYER M1 ;
  END Z
END INVCLKHDUX

MACRO INVHD12X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  4.9374 LAYER M1 ;
  END Z
END INVHD12X

MACRO INVHD16X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4875 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  6.5832 LAYER M1 ;
  END Z
END INVHD16X

MACRO INVHD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END INVHD1X

MACRO INVHD1XSPG
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
    AntennaGateArea  0.2743 LAYER M2 ;
    AntennaGateArea  0.2743 LAYER M3 ;
    AntennaGateArea  0.2743 LAYER M4 ;
    AntennaGateArea  0.2743 LAYER M5 ;
    AntennaGateArea  0.2743 LAYER M6 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
    AntennaDiffArea  0.72795 LAYER M2 ;
    AntennaDiffArea  0.72795 LAYER M3 ;
    AntennaDiffArea  0.72795 LAYER M4 ;
    AntennaDiffArea  0.72795 LAYER M5 ;
    AntennaDiffArea  0.72795 LAYER M6 ;
  END Z
END INVHD1XSPG

MACRO INVHD20X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  8.862 LAYER M1 ;
  END Z
END INVHD20X

MACRO INVHD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END INVHD2X

MACRO INVHD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.8229 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END INVHD3X

MACRO INVHD4X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.0972 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.6458 LAYER M1 ;
  END Z
END INVHD4X

MACRO INVHD5X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.3715 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.37375 LAYER M1 ;
  END Z
END INVHD5X

MACRO INVHD6X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.6458 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.4687 LAYER M1 ;
  END Z
END INVHD6X

MACRO INVHD7X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.9201 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.19665 LAYER M1 ;
  END Z
END INVHD7X

MACRO INVHD8X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  2.1944 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.2916 LAYER M1 ;
  END Z
END INVHD8X

MACRO INVHDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
END INVHDLX

MACRO INVHDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1404 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END INVHDMX

MACRO INVHDPX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6555 LAYER M1 ;
  END Z
END INVHDPX

MACRO INVHDUX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0624 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2246 LAYER M1 ;
  END Z
END INVHDUX

MACRO INVODHD8X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN Z0
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z0
  PIN Z1
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z1
  PIN Z2
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z2
  PIN Z3
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z3
  PIN Z4
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z4
  PIN Z5
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z5
  PIN Z6
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z6
  PIN Z7
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z7
END INVODHD8X

MACRO INVTSHD12X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.6578 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  5.5704 LAYER M1 ;
  END Z
END INVTSHD12X

MACRO INVTSHD16X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  1.0335 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  7.2162 LAYER M1 ;
  END Z
END INVTSHD16X

MACRO INVTSHD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4459 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2587 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6694 LAYER M1 ;
  END Z
END INVTSHD1X

MACRO INVTSHD20X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  1.209 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  8.862 LAYER M1 ;
  END Z
END INVTSHD20X

MACRO INVTSHD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.8918 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.5174 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.3388 LAYER M1 ;
  END Z
END INVTSHD2X

MACRO INVTSHD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.2349 LAYER M1 ;
  END Z
END INVTSHD3X

MACRO INVTSHD4X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1495 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.299 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.89385 LAYER M1 ;
  END Z
END INVTSHD4X

MACRO INVTSHD5X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1677 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.3432 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.06505 LAYER M1 ;
  END Z
END INVTSHD5X

MACRO INVTSHD6X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1833 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.3705 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.74215 LAYER M1 ;
  END Z
END INVTSHD6X

MACRO INVTSHD7X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.442 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.88195 LAYER M1 ;
  END Z
END INVTSHD7X

MACRO INVTSHD8X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.4186 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.9246 LAYER M1 ;
  END Z
END INVTSHD8X

MACRO INVTSHDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1534 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1456 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4071 LAYER M1 ;
  END Z
END INVTSHDLX

MACRO INVTSHDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2288 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1703 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6072 LAYER M1 ;
  END Z
END INVTSHDMX

MACRO INVTSHDUX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1014 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.0962 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2889 LAYER M1 ;
  END Z
END INVTSHDUX

MACRO LATHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
END LATHD1X

MACRO LATHD1XSPG
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
    AntennaDiffArea  0.72795 LAYER M2 ;
    AntennaDiffArea  0.72795 LAYER M3 ;
    AntennaDiffArea  0.72795 LAYER M4 ;
    AntennaDiffArea  0.72795 LAYER M5 ;
    AntennaDiffArea  0.72795 LAYER M6 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
    AntennaDiffArea  0.72795 LAYER M2 ;
    AntennaDiffArea  0.72795 LAYER M3 ;
    AntennaDiffArea  0.72795 LAYER M4 ;
    AntennaDiffArea  0.72795 LAYER M5 ;
    AntennaDiffArea  0.72795 LAYER M6 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
    AntennaGateArea  0.156 LAYER M2 ;
    AntennaGateArea  0.156 LAYER M3 ;
    AntennaGateArea  0.156 LAYER M4 ;
    AntennaGateArea  0.156 LAYER M5 ;
    AntennaGateArea  0.156 LAYER M6 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
    AntennaGateArea  0.117 LAYER M2 ;
    AntennaGateArea  0.117 LAYER M3 ;
    AntennaGateArea  0.117 LAYER M4 ;
    AntennaGateArea  0.117 LAYER M5 ;
    AntennaGateArea  0.117 LAYER M6 ;
  END G
END LATHD1XSPG

MACRO LATHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2405 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
END LATHD2X

MACRO LATHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2442 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2589 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END G
END LATHDLX

MACRO LATHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END G
END LATHDMX

MACRO LATNHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
END LATNHD1X

MACRO LATNHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2405 LAYER M1 ;
  END D
END LATNHD2X

MACRO LATNHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
END LATNHDLX

MACRO LATNHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
END LATNHDMX

MACRO LATNRHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6396 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2288 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END RN
END LATNRHD1X

MACRO LATNRHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3523 LAYER M1 ;
  END RN
END LATNRHD2X

MACRO LATNRHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2376 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1508 LAYER M1 ;
  END RN
END LATNRHDLX

MACRO LATNRHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.34125 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2132 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2145 LAYER M1 ;
  END RN
END LATNRHDMX

MACRO LATNSHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.67285 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
  END D
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END LATNSHD1X

MACRO LATNSHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1261 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
  END D
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END SN
END LATNSHD2X

MACRO LATNSHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1885 LAYER M1 ;
  END D
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END LATNSHDLX

MACRO LATNSHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.35835 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2262 LAYER M1 ;
  END D
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END LATNSHDMX

MACRO LATNSRHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6168 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6814 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2652 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END SN
END LATNSRHD1X

MACRO LATNSRHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3523 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END SN
END LATNSRHD2X

MACRO LATNSRHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.221 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END LATNSRHDLX

MACRO LATNSRHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2652 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END SN
END LATNSRHDMX

MACRO LATRHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6396 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2288 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END RN
END LATRHD1X

MACRO LATRHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3523 LAYER M1 ;
  END RN
END LATRHD2X

MACRO LATRHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END G
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1508 LAYER M1 ;
  END RN
END LATRHDLX

MACRO LATRHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.34125 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2132 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2145 LAYER M1 ;
  END RN
END LATRHDMX

MACRO LATSHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.67285 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END LATSHD1X

MACRO LATSHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END SN
END LATSHD2X

MACRO LATSHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1885 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END G
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END LATSHDLX

MACRO LATSHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.35835 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2262 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END LATSHDMX

MACRO LATSRHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6168 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6814 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2652 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END SN
END LATSRHD1X

MACRO LATSRHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3523 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END SN
END LATSRHD2X

MACRO LATSRHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END G
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.221 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END LATSRHDLX

MACRO LATSRHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2652 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END SN
END LATSRHDMX

MACRO LATTSHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.3938 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.312 LAYER M1 ;
  END E
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
END LATTSHD1X

MACRO LATTSHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END E
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
END LATTSHD2X

MACRO LATTSHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.32515 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1456 LAYER M1 ;
  END E
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END G
END LATTSHDLX

MACRO LATTSHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4968 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END E
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
END LATTSHDMX

MACRO MUX2CLKHD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5865 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END S0
END MUX2CLKHD1X

MACRO MUX2CLKHD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.69615 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END S0
END MUX2CLKHD2X

MACRO MUX2CLKHD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2197 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2197 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.30605 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.3133 LAYER M1 ;
  END S0
END MUX2CLKHD3X

MACRO MUX2CLKHD4X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.312 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.312 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.3701 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.4056 LAYER M1 ;
  END S0
END MUX2CLKHD4X

MACRO MUX2HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2184 LAYER M1 ;
  END S0
END MUX2HD1X

MACRO MUX2HD1XSPG
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
    AntennaGateArea  0.1248 LAYER M2 ;
    AntennaGateArea  0.1248 LAYER M3 ;
    AntennaGateArea  0.1248 LAYER M4 ;
    AntennaGateArea  0.1248 LAYER M5 ;
    AntennaGateArea  0.1248 LAYER M6 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
    AntennaGateArea  0.1248 LAYER M2 ;
    AntennaGateArea  0.1248 LAYER M3 ;
    AntennaGateArea  0.1248 LAYER M4 ;
    AntennaGateArea  0.1248 LAYER M5 ;
    AntennaGateArea  0.1248 LAYER M6 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
    AntennaDiffArea  0.72795 LAYER M2 ;
    AntennaDiffArea  0.72795 LAYER M3 ;
    AntennaDiffArea  0.72795 LAYER M4 ;
    AntennaDiffArea  0.72795 LAYER M5 ;
    AntennaDiffArea  0.72795 LAYER M6 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2184 LAYER M1 ;
    AntennaGateArea  0.2184 LAYER M2 ;
    AntennaGateArea  0.2184 LAYER M3 ;
    AntennaGateArea  0.2184 LAYER M4 ;
    AntennaGateArea  0.2184 LAYER M5 ;
    AntennaGateArea  0.2184 LAYER M6 ;
  END S0
END MUX2HD1XSPG

MACRO MUX2HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.89675 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.3432 LAYER M1 ;
  END S0
END MUX2HD2X

MACRO MUX2HD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.3679 LAYER M1 ;
  END S0
END MUX2HD3X

MACRO MUX2HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S0
END MUX2HDLX

MACRO MUX2HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S0
END MUX2HDMX

MACRO MUX2HDUX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0624 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0624 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.461 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END S0
END MUX2HDUX

MACRO MUX4HD1X
  PIN S1
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S1
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6814 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END S0
END MUX4HD1X

MACRO MUX4HD2X
  PIN S1
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S1
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END S0
END MUX4HD2X

MACRO MUX4HDLX
  PIN S1
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S1
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END S0
END MUX4HDLX

MACRO MUX4HDMX
  PIN S1
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S1
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END S0
END MUX4HDMX

MACRO MUXI2HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S0
END MUXI2HD1X

MACRO MUXI2HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S0
END MUXI2HD2X

MACRO MUXI2HD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S0
END MUXI2HD3X

MACRO MUXI2HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S0
END MUXI2HDLX

MACRO MUXI2HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S0
END MUXI2HDMX

MACRO MUXI4HD1X
  PIN S1
    #DIRECTION INPUT ;
    AntennaGateArea  0.2184 LAYER M1 ;
  END S1
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END S0
END MUXI4HD1X

MACRO MUXI4HD2X
  PIN S1
    #DIRECTION INPUT ;
    AntennaGateArea  0.3432 LAYER M1 ;
  END S1
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.3198 LAYER M1 ;
  END S0
END MUXI4HD2X

MACRO MUXI4HDLX
  PIN S1
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S1
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END S0
END MUXI4HDLX

MACRO MUXI4HDMX
  PIN S1
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S1
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END S0
END MUXI4HDMX

MACRO NAND2B1HD1X
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.717 LAYER M1 ;
  END Z
END NAND2B1HD1X

MACRO NAND2B1HD2X
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.5044 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1404 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.17 LAYER M1 ;
  END Z
END NAND2B1HD2X

MACRO NAND2B1HDLX
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2439 LAYER M1 ;
  END Z
END NAND2B1HDLX

MACRO NAND2B1HDMX
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1508 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4067 LAYER M1 ;
  END Z
END NAND2B1HDMX

MACRO NAND2B1HDUX
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0624 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.318 LAYER M1 ;
  END Z
END NAND2B1HDUX

MACRO NAND2HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.0438 LAYER M1 ;
  END Z
END NAND2HD1X

MACRO NAND2HD1XSPG
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
    AntennaGateArea  0.2522 LAYER M2 ;
    AntennaGateArea  0.2522 LAYER M3 ;
    AntennaGateArea  0.2522 LAYER M4 ;
    AntennaGateArea  0.2522 LAYER M5 ;
    AntennaGateArea  0.2522 LAYER M6 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
    AntennaGateArea  0.2522 LAYER M2 ;
    AntennaGateArea  0.2522 LAYER M3 ;
    AntennaGateArea  0.2522 LAYER M4 ;
    AntennaGateArea  0.2522 LAYER M5 ;
    AntennaGateArea  0.2522 LAYER M6 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.0186 LAYER M1 ;
    AntennaDiffArea  1.0186 LAYER M2 ;
    AntennaDiffArea  1.0186 LAYER M3 ;
    AntennaDiffArea  1.0186 LAYER M4 ;
    AntennaDiffArea  1.0186 LAYER M5 ;
    AntennaDiffArea  1.0186 LAYER M6 ;
  END Z
END NAND2HD1XSPG

MACRO NAND2HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5044 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.5044 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.17 LAYER M1 ;
  END Z
END NAND2HD2X

MACRO NAND2HD2XSPG
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5044 LAYER M1 ;
    AntennaGateArea  0.5044 LAYER M2 ;
    AntennaGateArea  0.5044 LAYER M3 ;
    AntennaGateArea  0.5044 LAYER M4 ;
    AntennaGateArea  0.5044 LAYER M5 ;
    AntennaGateArea  0.5044 LAYER M6 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.5044 LAYER M1 ;
    AntennaGateArea  0.5044 LAYER M2 ;
    AntennaGateArea  0.5044 LAYER M3 ;
    AntennaGateArea  0.5044 LAYER M4 ;
    AntennaGateArea  0.5044 LAYER M5 ;
    AntennaGateArea  0.5044 LAYER M6 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.17 LAYER M1 ;
    AntennaDiffArea  1.17 LAYER M2 ;
    AntennaDiffArea  1.17 LAYER M3 ;
    AntennaDiffArea  1.17 LAYER M4 ;
    AntennaDiffArea  1.17 LAYER M5 ;
    AntennaDiffArea  1.17 LAYER M6 ;
  END Z
END NAND2HD2XSPG

MACRO NAND2HD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.7566 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.7566 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.205 LAYER M1 ;
  END Z
END NAND2HD3X

MACRO NAND2HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2439 LAYER M1 ;
  END Z
END NAND2HDLX

MACRO NAND2HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1508 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1508 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.42855 LAYER M1 ;
  END Z
END NAND2HDMX

MACRO NAND2HDUX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0676 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0676 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.321 LAYER M1 ;
  END Z
END NAND2HDUX

MACRO NAND2ODHD
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z
END NAND2ODHD

MACRO NAND3B1HD1X
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2288 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2288 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.9548 LAYER M1 ;
  END Z
END NAND3B1HD1X

MACRO NAND3B1HD2X
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NAND3B1HD2X

MACRO NAND3B1HDLX
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4705 LAYER M1 ;
  END Z
END NAND3B1HDLX

MACRO NAND3B1HDMX
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.78895 LAYER M1 ;
  END Z
END NAND3B1HDMX

MACRO NAND3HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2288 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2288 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2288 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.9352 LAYER M1 ;
  END Z
END NAND3HD1X

MACRO NAND3HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NAND3HD2X

MACRO NAND3HD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END NAND3HD3X

MACRO NAND3HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3285 LAYER M1 ;
  END Z
END NAND3HDLX

MACRO NAND3HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.68985 LAYER M1 ;
  END Z
END NAND3HDMX

MACRO NAND3ODHD
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z
END NAND3ODHD

MACRO NAND4B1HD1X
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END NAND4B1HD1X

MACRO NAND4B1HD2X
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NAND4B1HD2X

MACRO NAND4B1HDLX
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.471 LAYER M1 ;
  END Z
END NAND4B1HDLX

MACRO NAND4B1HDMX
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.7329 LAYER M1 ;
  END Z
END NAND4B1HDMX

MACRO NAND4B2HD1X
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END NAND4B2HD1X

MACRO NAND4B2HD2X
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NAND4B2HD2X

MACRO NAND4B2HDLX
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.345 LAYER M1 ;
  END Z
END NAND4B2HDLX

MACRO NAND4B2HDMX
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.7272 LAYER M1 ;
  END Z
END NAND4B2HDMX

MACRO NAND4HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END NAND4HD1X

MACRO NAND4HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NAND4HD2X

MACRO NAND4HD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END NAND4HD3X

MACRO NAND4HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.34785 LAYER M1 ;
  END Z
END NAND4HDLX

MACRO NAND4HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6949 LAYER M1 ;
  END Z
END NAND4HDMX

MACRO NOR2B1HD1X
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.67395 LAYER M1 ;
  END Z
END NOR2B1HD1X

MACRO NOR2B1HD2X
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.4862 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1404 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.9789 LAYER M1 ;
  END Z
END NOR2B1HD2X

MACRO NOR2B1HDLX
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3165 LAYER M1 ;
  END Z
END NOR2B1HDLX

MACRO NOR2B1HDMX
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1703 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4765 LAYER M1 ;
  END Z
END NOR2B1HDMX

MACRO NOR2B1HDUX
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0754 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0624 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2511 LAYER M1 ;
  END Z
END NOR2B1HDUX

MACRO NOR2HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6801 LAYER M1 ;
  END Z
END NOR2HD1X

MACRO NOR2HD1XSPG
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
    AntennaGateArea  0.2431 LAYER M2 ;
    AntennaGateArea  0.2431 LAYER M3 ;
    AntennaGateArea  0.2431 LAYER M4 ;
    AntennaGateArea  0.2431 LAYER M5 ;
    AntennaGateArea  0.2431 LAYER M6 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
    AntennaGateArea  0.2431 LAYER M2 ;
    AntennaGateArea  0.2431 LAYER M3 ;
    AntennaGateArea  0.2431 LAYER M4 ;
    AntennaGateArea  0.2431 LAYER M5 ;
    AntennaGateArea  0.2431 LAYER M6 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6801 LAYER M1 ;
    AntennaDiffArea  0.6801 LAYER M2 ;
    AntennaDiffArea  0.6801 LAYER M3 ;
    AntennaDiffArea  0.6801 LAYER M4 ;
    AntennaDiffArea  0.6801 LAYER M5 ;
    AntennaDiffArea  0.6801 LAYER M6 ;
  END Z
END NOR2HD1XSPG

MACRO NOR2HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4862 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.4862 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.0286 LAYER M1 ;
  END Z
END NOR2HD2X

MACRO NOR2HD2XSPG
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4862 LAYER M1 ;
    AntennaGateArea  0.4862 LAYER M2 ;
    AntennaGateArea  0.4862 LAYER M3 ;
    AntennaGateArea  0.4862 LAYER M4 ;
    AntennaGateArea  0.4862 LAYER M5 ;
    AntennaGateArea  0.4862 LAYER M6 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.4862 LAYER M1 ;
    AntennaGateArea  0.4862 LAYER M2 ;
    AntennaGateArea  0.4862 LAYER M3 ;
    AntennaGateArea  0.4862 LAYER M4 ;
    AntennaGateArea  0.4862 LAYER M5 ;
    AntennaGateArea  0.4862 LAYER M6 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.0286 LAYER M1 ;
    AntennaDiffArea  1.0286 LAYER M2 ;
    AntennaDiffArea  1.0286 LAYER M3 ;
    AntennaDiffArea  1.0286 LAYER M4 ;
    AntennaDiffArea  1.0286 LAYER M5 ;
    AntennaDiffArea  1.0286 LAYER M6 ;
  END Z
END NOR2HD2XSPG

MACRO NOR2HD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.7332 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.7332 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.87255 LAYER M1 ;
  END Z
END NOR2HD3X

MACRO NOR2HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.31365 LAYER M1 ;
  END Z
END NOR2HDLX

MACRO NOR2HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1703 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1703 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4722 LAYER M1 ;
  END Z
END NOR2HDMX

MACRO NOR2HDUX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0754 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0754 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4029 LAYER M1 ;
  END Z
END NOR2HDUX

MACRO NOR3B1HD1X
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.83595 LAYER M1 ;
  END Z
END NOR3B1HD1X

MACRO NOR3B1HD2X
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NOR3B1HD2X

MACRO NOR3B1HDLX
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5943 LAYER M1 ;
  END Z
END NOR3B1HDLX

MACRO NOR3B1HDMX
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.65805 LAYER M1 ;
  END Z
END NOR3B1HDMX

MACRO NOR3HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.83595 LAYER M1 ;
  END Z
END NOR3HD1X

MACRO NOR3HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NOR3HD2X

MACRO NOR3HD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END NOR3HD3X

MACRO NOR3HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4463 LAYER M1 ;
  END Z
END NOR3HDLX

MACRO NOR3HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6723 LAYER M1 ;
  END Z
END NOR3HDMX

MACRO NOR4B1HD1X
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END NOR4B1HD1X

MACRO NOR4B1HD2X
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NOR4B1HD2X

MACRO NOR4B1HDLX
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.62025 LAYER M1 ;
  END Z
END NOR4B1HDLX

MACRO NOR4B1HDMX
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.93295 LAYER M1 ;
  END Z
END NOR4B1HDMX

MACRO NOR4B2HD1X
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.7042 LAYER M1 ;
  END Z
END NOR4B2HD1X

MACRO NOR4B2HD2X
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NOR4B2HD2X

MACRO NOR4B2HDLX
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.49275 LAYER M1 ;
  END Z
END NOR4B2HDLX

MACRO NOR4B2HDMX
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.74085 LAYER M1 ;
  END Z
END NOR4B2HDMX

MACRO NOR4HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END NOR4HD1X

MACRO NOR4HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NOR4HD2X

MACRO NOR4HD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END NOR4HD3X

MACRO NOR4HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.53025 LAYER M1 ;
  END Z
END NOR4HDLX

MACRO NOR4HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.79715 LAYER M1 ;
  END Z
END NOR4HDMX

MACRO OAI211HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1976 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1976 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.999 LAYER M1 ;
  END Z
END OAI211HD1X

MACRO OAI211HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0897 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0897 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OAI211HD2X

MACRO OAI211HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0897 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0897 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4503 LAYER M1 ;
  END Z
END OAI211HDLX

MACRO OAI211HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1274 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1274 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.63945 LAYER M1 ;
  END Z
END OAI211HDMX

MACRO OAI21B2HD1X
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
  END C
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.717 LAYER M1 ;
  END Z
END OAI21B2HD1X

MACRO OAI21B2HD2X
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1261 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.5044 LAYER M1 ;
  END C
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1261 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.17 LAYER M1 ;
  END Z
END OAI21B2HD2X

MACRO OAI21B2HDLX
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END C
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2439 LAYER M1 ;
  END Z
END OAI21B2HDLX

MACRO OAI21B2HDMX
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1508 LAYER M1 ;
  END C
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4067 LAYER M1 ;
  END Z
END OAI21B2HDMX

MACRO OAI21HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2015 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8028 LAYER M1 ;
  END Z
END OAI21HD1X

MACRO OAI21HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1261 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1261 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OAI21HD2X

MACRO OAI21HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1261 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1261 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.36165 LAYER M1 ;
  END Z
END OAI21HDLX

MACRO OAI21HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2171 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2171 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1508 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6234 LAYER M1 ;
  END Z
END OAI21HDMX

MACRO OAI21HDUX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3588 LAYER M1 ;
  END Z
END OAI21HDUX

MACRO OAI221HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1976 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.041 LAYER M1 ;
  END Z
END OAI221HD1X

MACRO OAI221HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.0897 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OAI221HD2X

MACRO OAI221HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.0897 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.45255 LAYER M1 ;
  END Z
END OAI221HDLX

MACRO OAI221HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1274 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6423 LAYER M1 ;
  END Z
END OAI221HDMX

MACRO OAI222HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.2795 LAYER M1 ;
  END Z
END OAI222HD1X

MACRO OAI222HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OAI222HD2X

MACRO OAI222HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.54855 LAYER M1 ;
  END Z
END OAI222HDLX

MACRO OAI222HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.74135 LAYER M1 ;
  END Z
END OAI222HDMX

MACRO OAI22B2HD1X
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.7947 LAYER M1 ;
  END Z
END OAI22B2HD1X

MACRO OAI22B2HD2X
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.5084 LAYER M1 ;
  END Z
END OAI22B2HD2X

MACRO OAI22B2HDLX
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3819 LAYER M1 ;
  END Z
END OAI22B2HDLX

MACRO OAI22B2HDMX
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1937 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1937 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5196 LAYER M1 ;
  END Z
END OAI22B2HDMX

MACRO OAI22HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.91515 LAYER M1 ;
  END Z
END OAI22HD1X

MACRO OAI22HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OAI22HD2X

MACRO OAI22HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2925 LAYER M1 ;
  END Z
END OAI22HDLX

MACRO OAI22HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.429 LAYER M1 ;
  END Z
END OAI22HDMX

MACRO OAI22HDUX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2772 LAYER M1 ;
  END Z
END OAI22HDUX

MACRO OAI31HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0806 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END OAI31HD1X

MACRO OAI31HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0806 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OAI31HD2X

MACRO OAI31HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0806 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4587 LAYER M1 ;
  END Z
END OAI31HDLX

MACRO OAI31HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.104 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.58965 LAYER M1 ;
  END Z
END OAI31HDMX

MACRO OAI32HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END OAI32HD1X

MACRO OAI32HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OAI32HD2X

MACRO OAI32HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4932 LAYER M1 ;
  END Z
END OAI32HDLX

MACRO OAI32HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1495 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1495 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.63345 LAYER M1 ;
  END Z
END OAI32HDMX

MACRO OAI33HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END OAI33HD1X

MACRO OAI33HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OAI33HD2X

MACRO OAI33HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6237 LAYER M1 ;
  END Z
END OAI33HDLX

MACRO OAI33HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.80325 LAYER M1 ;
  END Z
END OAI33HDMX

MACRO OR2HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72315 LAYER M1 ;
  END Z
END OR2HD1X

MACRO OR2HD1XSPG
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
    AntennaGateArea  0.1131 LAYER M2 ;
    AntennaGateArea  0.1131 LAYER M3 ;
    AntennaGateArea  0.1131 LAYER M4 ;
    AntennaGateArea  0.1131 LAYER M5 ;
    AntennaGateArea  0.1131 LAYER M6 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
    AntennaGateArea  0.1131 LAYER M2 ;
    AntennaGateArea  0.1131 LAYER M3 ;
    AntennaGateArea  0.1131 LAYER M4 ;
    AntennaGateArea  0.1131 LAYER M5 ;
    AntennaGateArea  0.1131 LAYER M6 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72315 LAYER M1 ;
    AntennaDiffArea  0.72315 LAYER M2 ;
    AntennaDiffArea  0.72315 LAYER M3 ;
    AntennaDiffArea  0.72315 LAYER M4 ;
    AntennaDiffArea  0.72315 LAYER M5 ;
    AntennaDiffArea  0.72315 LAYER M6 ;
  END Z
END OR2HD1XSPG

MACRO OR2HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2262 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2262 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OR2HD2X

MACRO OR2HD2XSPG
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2262 LAYER M1 ;
    AntennaGateArea  0.2262 LAYER M2 ;
    AntennaGateArea  0.2262 LAYER M3 ;
    AntennaGateArea  0.2262 LAYER M4 ;
    AntennaGateArea  0.2262 LAYER M5 ;
    AntennaGateArea  0.2262 LAYER M6 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2262 LAYER M1 ;
    AntennaGateArea  0.2262 LAYER M2 ;
    AntennaGateArea  0.2262 LAYER M3 ;
    AntennaGateArea  0.2262 LAYER M4 ;
    AntennaGateArea  0.2262 LAYER M5 ;
    AntennaGateArea  0.2262 LAYER M6 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
    AntennaDiffArea  0.8229 LAYER M2 ;
    AntennaDiffArea  0.8229 LAYER M3 ;
    AntennaDiffArea  0.8229 LAYER M4 ;
    AntennaDiffArea  0.8229 LAYER M5 ;
    AntennaDiffArea  0.8229 LAYER M6 ;
  END Z
END OR2HD2XSPG

MACRO OR2HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
END OR2HDLX

MACRO OR2HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END OR2HDMX

MACRO OR2HDUX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0754 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0754 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3249 LAYER M1 ;
  END Z
END OR2HDUX

MACRO OR2ODHD
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1508 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1508 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6468 LAYER M1 ;
  END Z
END OR2ODHD

MACRO OR3HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END OR3HD1X

MACRO OR3HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OR3HD2X

MACRO OR3HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
END OR3HDLX

MACRO OR3HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END OR3HDMX

MACRO OR4HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END OR4HD1X

MACRO OR4HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2236 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2236 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2236 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2236 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OR4HD2X

MACRO OR4HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
END OR4HDLX

MACRO OR4HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END OR4HDMX

MACRO PULLDHD
  PIN EN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END EN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.1095 LAYER M1 ;
  END Z
END PULLDHD

MACRO PULLUHD
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.1095 LAYER M1 ;
  END Z
END PULLUHD

MACRO RSLATHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.65545 LAYER M1 ;
  END Q
  PIN R
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END R
  PIN S
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END S
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6213 LAYER M1 ;
  END QN
END RSLATHD1X

MACRO RSLATHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8844 LAYER M1 ;
  END Q
  PIN R
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END R
  PIN S
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END S
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.97665 LAYER M1 ;
  END QN
END RSLATHD2X

MACRO RSLATHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.252 LAYER M1 ;
  END Q
  PIN R
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END R
  PIN S
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END S
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2415 LAYER M1 ;
  END QN
END RSLATHDLX

MACRO RSLATHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.342 LAYER M1 ;
  END Q
  PIN R
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END R
  PIN S
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END S
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3315 LAYER M1 ;
  END QN
END RSLATHDMX

MACRO RSLATNHD1X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5875 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5845 LAYER M1 ;
  END QN
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END RSLATNHD1X

MACRO RSLATNHD2X
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8977 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END RSLATNHD2X

MACRO RSLATNHDLX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2514 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END RSLATNHDLX

MACRO RSLATNHDMX
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3414 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END QN
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END RSLATNHDMX

MACRO TIEHHD
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.132 LAYER M1 ;
  END Z
END TIEHHD

MACRO TIELHD
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.1245 LAYER M1 ;
  END Z
END TIELHD

MACRO XNOR2HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1092 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.77015 LAYER M1 ;
  END Z
END XNOR2HD1X

MACRO XNOR2HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.3016 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END XNOR2HD2X

MACRO XNOR2HD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.3315 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END XNOR2HD3X

MACRO XNOR2HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2628 LAYER M1 ;
  END Z
END XNOR2HDLX

MACRO XNOR2HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3942 LAYER M1 ;
  END Z
END XNOR2HDMX

MACRO XNOR3HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1092 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.74905 LAYER M1 ;
  END Z
END XNOR3HD1X

MACRO XNOR3HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1755 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1027 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END XNOR3HD2X

MACRO XNOR3HD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1755 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1027 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END XNOR3HD3X

MACRO XNOR3HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2556 LAYER M1 ;
  END Z
END XNOR3HDLX

MACRO XNOR3HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3834 LAYER M1 ;
  END Z
END XNOR3HDMX

MACRO XOR2CLKHD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2145 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5865 LAYER M1 ;
  END Z
END XOR2CLKHD1X

MACRO XOR2CLKHD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2145 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.68835 LAYER M1 ;
  END Z
END XOR2CLKHD2X

MACRO XOR2CLKHD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.221 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.29383 LAYER M1 ;
  END Z
END XOR2CLKHD3X

MACRO XOR2CLKHD4X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.325 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2717 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.3884 LAYER M1 ;
  END Z
END XOR2CLKHD4X

MACRO XOR2HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1846 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1092 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END XOR2HD1X

MACRO XOR2HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.26 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END XOR2HD2X

MACRO XOR2HD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.286 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END XOR2HD3X

MACRO XOR2HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
END XOR2HDLX

MACRO XOR2HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END XOR2HDMX

MACRO XOR3HD1X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1092 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.76485 LAYER M1 ;
  END Z
END XOR3HD1X

MACRO XOR3HD2X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8862 LAYER M1 ;
  END Z
END XOR3HD2X

MACRO XOR3HD3X
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END XOR3HD3X

MACRO XOR3HDLX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
END XOR3HDLX

MACRO XOR3HDMX
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END XOR3HDMX

END LIBRARY
