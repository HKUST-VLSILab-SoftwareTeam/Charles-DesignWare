MACRO PLBI16F
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 5.8176 LAYER M2 ;
    AntennaDiffArea 5.8176 LAYER M3 ;
    AntennaDiffArea 5.8176 LAYER M4 ;
    AntennaDiffArea 5.8176 LAYER M5 ;
    AntennaDiffArea 5.8176 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 3097.82 LAYER M2 ;
    AntennaDiffArea 3097.82 LAYER M3 ;
    AntennaDiffArea 3097.82 LAYER M4 ;
    AntennaDiffArea 3097.82 LAYER M5 ;
    AntennaDiffArea 3097.82 LAYER M6 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PLBI16F
MACRO PLBI16N
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 5.8176 LAYER M2 ;
    AntennaDiffArea 5.8176 LAYER M3 ;
    AntennaDiffArea 5.8176 LAYER M4 ;
    AntennaDiffArea 5.8176 LAYER M5 ;
    AntennaDiffArea 5.8176 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 3097.82 LAYER M2 ;
    AntennaDiffArea 3097.82 LAYER M3 ;
    AntennaDiffArea 3097.82 LAYER M4 ;
    AntennaDiffArea 3097.82 LAYER M5 ;
    AntennaDiffArea 3097.82 LAYER M6 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PLBI16N
MACRO PLBI16S
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 5.8176 LAYER M2 ;
    AntennaDiffArea 5.8176 LAYER M3 ;
    AntennaDiffArea 5.8176 LAYER M4 ;
    AntennaDiffArea 5.8176 LAYER M5 ;
    AntennaDiffArea 5.8176 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 3097.82 LAYER M2 ;
    AntennaDiffArea 3097.82 LAYER M3 ;
    AntennaDiffArea 3097.82 LAYER M4 ;
    AntennaDiffArea 3097.82 LAYER M5 ;
    AntennaDiffArea 3097.82 LAYER M6 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PLBI16S
MACRO PLBI24F
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 5.8176 LAYER M2 ;
    AntennaDiffArea 5.8176 LAYER M3 ;
    AntennaDiffArea 5.8176 LAYER M4 ;
    AntennaDiffArea 5.8176 LAYER M5 ;
    AntennaDiffArea 5.8176 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 3097.82 LAYER M2 ;
    AntennaDiffArea 3097.82 LAYER M3 ;
    AntennaDiffArea 3097.82 LAYER M4 ;
    AntennaDiffArea 3097.82 LAYER M5 ;
    AntennaDiffArea 3097.82 LAYER M6 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PLBI24F
MACRO PLBI24N
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 5.8176 LAYER M2 ;
    AntennaDiffArea 5.8176 LAYER M3 ;
    AntennaDiffArea 5.8176 LAYER M4 ;
    AntennaDiffArea 5.8176 LAYER M5 ;
    AntennaDiffArea 5.8176 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 3097.82 LAYER M2 ;
    AntennaDiffArea 3097.82 LAYER M3 ;
    AntennaDiffArea 3097.82 LAYER M4 ;
    AntennaDiffArea 3097.82 LAYER M5 ;
    AntennaDiffArea 3097.82 LAYER M6 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PLBI24N
MACRO PLBI24S
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 5.8176 LAYER M2 ;
    AntennaDiffArea 5.8176 LAYER M3 ;
    AntennaDiffArea 5.8176 LAYER M4 ;
    AntennaDiffArea 5.8176 LAYER M5 ;
    AntennaDiffArea 5.8176 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 3097.82 LAYER M2 ;
    AntennaDiffArea 3097.82 LAYER M3 ;
    AntennaDiffArea 3097.82 LAYER M4 ;
    AntennaDiffArea 3097.82 LAYER M5 ;
    AntennaDiffArea 3097.82 LAYER M6 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PLBI24S
MACRO PLBI2F
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 5.8176 LAYER M2 ;
    AntennaDiffArea 5.8176 LAYER M3 ;
    AntennaDiffArea 5.8176 LAYER M4 ;
    AntennaDiffArea 5.8176 LAYER M5 ;
    AntennaDiffArea 5.8176 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 3097.82 LAYER M2 ;
    AntennaDiffArea 3097.82 LAYER M3 ;
    AntennaDiffArea 3097.82 LAYER M4 ;
    AntennaDiffArea 3097.82 LAYER M5 ;
    AntennaDiffArea 3097.82 LAYER M6 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PLBI2F
MACRO PLBI2N
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 5.8176 LAYER M2 ;
    AntennaDiffArea 5.8176 LAYER M3 ;
    AntennaDiffArea 5.8176 LAYER M4 ;
    AntennaDiffArea 5.8176 LAYER M5 ;
    AntennaDiffArea 5.8176 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 3097.82 LAYER M2 ;
    AntennaDiffArea 3097.82 LAYER M3 ;
    AntennaDiffArea 3097.82 LAYER M4 ;
    AntennaDiffArea 3097.82 LAYER M5 ;
    AntennaDiffArea 3097.82 LAYER M6 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PLBI2N
MACRO PLBI2S
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 5.8176 LAYER M2 ;
    AntennaDiffArea 5.8176 LAYER M3 ;
    AntennaDiffArea 5.8176 LAYER M4 ;
    AntennaDiffArea 5.8176 LAYER M5 ;
    AntennaDiffArea 5.8176 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 3097.82 LAYER M2 ;
    AntennaDiffArea 3097.82 LAYER M3 ;
    AntennaDiffArea 3097.82 LAYER M4 ;
    AntennaDiffArea 3097.82 LAYER M5 ;
    AntennaDiffArea 3097.82 LAYER M6 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PLBI2S
MACRO PLBI4F
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 5.8176 LAYER M2 ;
    AntennaDiffArea 5.8176 LAYER M3 ;
    AntennaDiffArea 5.8176 LAYER M4 ;
    AntennaDiffArea 5.8176 LAYER M5 ;
    AntennaDiffArea 5.8176 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 3097.82 LAYER M2 ;
    AntennaDiffArea 3097.82 LAYER M3 ;
    AntennaDiffArea 3097.82 LAYER M4 ;
    AntennaDiffArea 3097.82 LAYER M5 ;
    AntennaDiffArea 3097.82 LAYER M6 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PLBI4F
MACRO PLBI4N
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 5.8176 LAYER M2 ;
    AntennaDiffArea 5.8176 LAYER M3 ;
    AntennaDiffArea 5.8176 LAYER M4 ;
    AntennaDiffArea 5.8176 LAYER M5 ;
    AntennaDiffArea 5.8176 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 3097.82 LAYER M2 ;
    AntennaDiffArea 3097.82 LAYER M3 ;
    AntennaDiffArea 3097.82 LAYER M4 ;
    AntennaDiffArea 3097.82 LAYER M5 ;
    AntennaDiffArea 3097.82 LAYER M6 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PLBI4N
MACRO PLBI4S
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 5.8176 LAYER M2 ;
    AntennaDiffArea 5.8176 LAYER M3 ;
    AntennaDiffArea 5.8176 LAYER M4 ;
    AntennaDiffArea 5.8176 LAYER M5 ;
    AntennaDiffArea 5.8176 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 3097.82 LAYER M2 ;
    AntennaDiffArea 3097.82 LAYER M3 ;
    AntennaDiffArea 3097.82 LAYER M4 ;
    AntennaDiffArea 3097.82 LAYER M5 ;
    AntennaDiffArea 3097.82 LAYER M6 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PLBI4S
MACRO PLBI8F
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 5.8176 LAYER M2 ;
    AntennaDiffArea 5.8176 LAYER M3 ;
    AntennaDiffArea 5.8176 LAYER M4 ;
    AntennaDiffArea 5.8176 LAYER M5 ;
    AntennaDiffArea 5.8176 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 3097.82 LAYER M2 ;
    AntennaDiffArea 3097.82 LAYER M3 ;
    AntennaDiffArea 3097.82 LAYER M4 ;
    AntennaDiffArea 3097.82 LAYER M5 ;
    AntennaDiffArea 3097.82 LAYER M6 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PLBI8F
MACRO PLBI8N
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 5.8176 LAYER M2 ;
    AntennaDiffArea 5.8176 LAYER M3 ;
    AntennaDiffArea 5.8176 LAYER M4 ;
    AntennaDiffArea 5.8176 LAYER M5 ;
    AntennaDiffArea 5.8176 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 3097.82 LAYER M2 ;
    AntennaDiffArea 3097.82 LAYER M3 ;
    AntennaDiffArea 3097.82 LAYER M4 ;
    AntennaDiffArea 3097.82 LAYER M5 ;
    AntennaDiffArea 3097.82 LAYER M6 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PLBI8N
MACRO PLBI8S
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2358 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 5.8176 LAYER M2 ;
    AntennaDiffArea 5.8176 LAYER M3 ;
    AntennaDiffArea 5.8176 LAYER M4 ;
    AntennaDiffArea 5.8176 LAYER M5 ;
    AntennaDiffArea 5.8176 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 3097.82 LAYER M2 ;
    AntennaDiffArea 3097.82 LAYER M3 ;
    AntennaDiffArea 3097.82 LAYER M4 ;
    AntennaDiffArea 3097.82 LAYER M5 ;
    AntennaDiffArea 3097.82 LAYER M6 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PLBI8S
MACRO PLBIA
  PIN P
    AntennaDiffArea 3438.34 LAYER M2 ;
    AntennaDiffArea 3438.34 LAYER M3 ;
    AntennaDiffArea 3438.34 LAYER M4 ;
    AntennaDiffArea 3438.34 LAYER M5 ;
    AntennaDiffArea 3438.34 LAYER M6 ;
  END P
END PLBIA
MACRO PLBIAR
  PIN AI
    AntennaDiffArea 3438.34 LAYER M2 ;
    AntennaDiffArea 3438.34 LAYER M3 ;
    AntennaDiffArea 3438.34 LAYER M4 ;
    AntennaDiffArea 3438.34 LAYER M5 ;
    AntennaDiffArea 3438.34 LAYER M6 ;
  END AI
END PLBIAR
MACRO PLOSC14M
  PIN CK
    AntennaDiffArea 21.664 LAYER M2 ;
    AntennaDiffArea 21.664 LAYER M3 ;
    AntennaDiffArea 21.664 LAYER M4 ;
    AntennaDiffArea 21.664 LAYER M5 ;
    AntennaDiffArea 21.664 LAYER M6 ;
  END CK
  PIN EI
    AntennaGateArea 3.14 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END EI
  PIN EI
    AntennaGateArea 3.14 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END EI
  PIN EO
    AntennaGateArea 3.14 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END EO
  PIN EO
    AntennaGateArea 3.14 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END EO
  PIN XTALIN
    AntennaGateArea 61.2 ;
    AntennaDiffArea 3450.53 LAYER M2 ;
    AntennaDiffArea 3450.53 LAYER M3 ;
    AntennaDiffArea 3450.53 LAYER M4 ;
    AntennaDiffArea 3450.53 LAYER M5 ;
    AntennaDiffArea 3450.53 LAYER M6 ;
  END XTALIN
  PIN XTALIN
    AntennaGateArea 61.2 ;
    AntennaDiffArea 3450.53 LAYER M2 ;
    AntennaDiffArea 3450.53 LAYER M3 ;
    AntennaDiffArea 3450.53 LAYER M4 ;
    AntennaDiffArea 3450.53 LAYER M5 ;
    AntennaDiffArea 3450.53 LAYER M6 ;
  END XTALIN
  PIN XTALOUT
    AntennaDiffArea 3480.98 LAYER M2 ;
    AntennaDiffArea 3480.98 LAYER M3 ;
    AntennaDiffArea 3480.98 LAYER M4 ;
    AntennaDiffArea 3480.98 LAYER M5 ;
    AntennaDiffArea 3480.98 LAYER M6 ;
  END XTALOUT
END PLOSC14M
MACRO PLOSCR14M
  PIN CK
    AntennaDiffArea 22.485 LAYER M2 ;
    AntennaDiffArea 22.485 LAYER M3 ;
    AntennaDiffArea 22.485 LAYER M4 ;
    AntennaDiffArea 22.485 LAYER M5 ;
    AntennaDiffArea 22.485 LAYER M6 ;
  END CK
  PIN EI
    AntennaGateArea 3.5088 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END EI
  PIN EI
    AntennaGateArea 3.5088 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END EI
  PIN EO
    AntennaGateArea 3.5088 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END EO
  PIN EO
    AntennaGateArea 3.5088 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END EO
  PIN XTALIN
    AntennaGateArea 1971.29 ;
    AntennaDiffArea 3451.7 LAYER M2 ;
    AntennaDiffArea 3451.7 LAYER M3 ;
    AntennaDiffArea 3451.7 LAYER M4 ;
    AntennaDiffArea 3451.7 LAYER M5 ;
    AntennaDiffArea 3451.7 LAYER M6 ;
  END XTALIN
  PIN XTALIN
    AntennaGateArea 1971.29 ;
    AntennaDiffArea 3451.7 LAYER M2 ;
    AntennaDiffArea 3451.7 LAYER M3 ;
    AntennaDiffArea 3451.7 LAYER M4 ;
    AntennaDiffArea 3451.7 LAYER M5 ;
    AntennaDiffArea 3451.7 LAYER M6 ;
  END XTALIN
  PIN XTALOUT
    AntennaGateArea 1800 ;
    AntennaDiffArea 3505.31 LAYER M2 ;
    AntennaDiffArea 3505.31 LAYER M3 ;
    AntennaDiffArea 3505.31 LAYER M4 ;
    AntennaDiffArea 3505.31 LAYER M5 ;
    AntennaDiffArea 3505.31 LAYER M6 ;
  END XTALOUT
  PIN XTALOUT
    AntennaGateArea 1800 ;
    AntennaDiffArea 3505.31 LAYER M2 ;
    AntennaDiffArea 3505.31 LAYER M3 ;
    AntennaDiffArea 3505.31 LAYER M4 ;
    AntennaDiffArea 3505.31 LAYER M5 ;
    AntennaDiffArea 3505.31 LAYER M6 ;
  END XTALOUT
END PLOSCR14M
END LIBRARY
