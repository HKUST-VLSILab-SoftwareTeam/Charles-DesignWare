VERSION 5.3.1 ;

LAYER M1
    ANTENNACUMAREARATIO  600 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 600 ) ( 0.249 600 ) ( 0.251 2300.4 ) ( 1 2600 ) ) ;
END M1

LAYER V1
    ANTENNACUMAREARATIO  20 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.249 20 ) ( 0.25 92.59 ) ( 1 160 ) ) ;
END V1

LAYER M2
    ANTENNACUMAREARATIO  600 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 600 ) ( 0.249 600 ) ( 0.25 2300.4 ) ( 1 2600 ) ) ;
END M2

LAYER V2
    ANTENNACUMAREARATIO  20 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.249 20 ) ( 0.25 92.59 ) ( 1 160 ) ) ;
END V2

LAYER M3
    ANTENNACUMAREARATIO  600 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 600 ) ( 0.249 600 ) ( 0.25  2300.4 ) ( 1 2600 ) ) ;
END M3

LAYER V3
    ANTENNACUMAREARATIO  20 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.249 20 ) ( 0.25 92.59 ) ( 1 160 ) ) ;
END V3

LAYER M4
    ANTENNACUMAREARATIO  600 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 600 ) ( 0.249 600 ) ( 0.25  2300.4 ) ( 1 2600 ) ) ;
END M4

LAYER V4
    ANTENNACUMAREARATIO  20 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.249 20 ) ( 0.25 92.59 ) ( 1 160 ) ) ;
END V4

LAYER M5
    ANTENNACUMAREARATIO  600 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 600 ) ( 0.249 600 ) ( 0.25  2300.4 ) ( 1 2600 ) ) ;
END M5

LAYER V5
    ANTENNACUMAREARATIO  20 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.249 20 ) ( 0.25 92.59 ) ( 1 160 ) ) ;
END V5

LAYER M6
    ANTENNACUMAREARATIO  600 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 600 ) ( 0.249 600 ) ( 0.25  2300.4 ) ( 1 2600 ) ) ;
END M6

LAYER V6
    ANTENNACUMAREARATIO  20 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.249 20 ) ( 0.25 92.59 ) ( 1 160 ) ) ;
END V6

LAYER M7
    ANTENNACUMAREARATIO  600 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 600 ) ( 0.249 600 ) ( 0.25  2300.4 ) ( 1 2600 ) ) ;
END M7

MACRO AND2CLKHD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.104 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.104 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5865 LAYER M1 ;
  END Z
END AND2CLKHD1XHT

MACRO AND2CLKHD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1664 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1664 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6747 LAYER M1 ;
  END Z
END AND2CLKHD2XHT

MACRO AND2CLKHD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.27155 LAYER M1 ;
  END Z
END AND2CLKHD3XHT

MACRO AND2CLKHD4XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2548 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2548 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.3494 LAYER M1 ;
  END Z
END AND2CLKHD4XHT

MACRO AND2HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END AND2HD1XHT

MACRO AND2HD1XSPGHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
    AntennaGateArea  0.0858 LAYER M2 ;
    AntennaGateArea  0.0858 LAYER M3 ;
    AntennaGateArea  0.0858 LAYER M4 ;
    AntennaGateArea  0.0858 LAYER M5 ;
    AntennaGateArea  0.0858 LAYER M6 ;
    AntennaGateArea  0.0858 LAYER M7 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
    AntennaGateArea  0.0858 LAYER M2 ;
    AntennaGateArea  0.0858 LAYER M3 ;
    AntennaGateArea  0.0858 LAYER M4 ;
    AntennaGateArea  0.0858 LAYER M5 ;
    AntennaGateArea  0.0858 LAYER M6 ;
    AntennaGateArea  0.0858 LAYER M7 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
    AntennaDiffArea  0.72795 LAYER M2 ;
    AntennaDiffArea  0.72795 LAYER M3 ;
    AntennaDiffArea  0.72795 LAYER M4 ;
    AntennaDiffArea  0.72795 LAYER M5 ;
    AntennaDiffArea  0.72795 LAYER M6 ;
    AntennaDiffArea  0.72795 LAYER M7 ;
  END Z
END AND2HD1XSPGHT

MACRO AND2HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1547 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1547 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END AND2HD2XHT

MACRO AND2HD2XSPGHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1547 LAYER M1 ;
    AntennaGateArea  0.1547 LAYER M2 ;
    AntennaGateArea  0.1547 LAYER M3 ;
    AntennaGateArea  0.1547 LAYER M4 ;
    AntennaGateArea  0.1547 LAYER M5 ;
    AntennaGateArea  0.1547 LAYER M6 ;
    AntennaGateArea  0.1547 LAYER M7 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1547 LAYER M1 ;
    AntennaGateArea  0.1547 LAYER M2 ;
    AntennaGateArea  0.1547 LAYER M3 ;
    AntennaGateArea  0.1547 LAYER M4 ;
    AntennaGateArea  0.1547 LAYER M5 ;
    AntennaGateArea  0.1547 LAYER M6 ;
    AntennaGateArea  0.1547 LAYER M7 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
    AntennaDiffArea  0.8229 LAYER M2 ;
    AntennaDiffArea  0.8229 LAYER M3 ;
    AntennaDiffArea  0.8229 LAYER M4 ;
    AntennaDiffArea  0.8229 LAYER M5 ;
    AntennaDiffArea  0.8229 LAYER M6 ;
    AntennaDiffArea  0.8229 LAYER M7 ;
  END Z
END AND2HD2XSPGHT

MACRO AND2HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
END AND2HDLXHT

MACRO AND2HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END AND2HDMXHT

MACRO AND2HDUXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.216 LAYER M1 ;
  END Z
END AND2HDUXHT

MACRO AND3HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0884 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0884 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0884 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END AND3HD1XHT

MACRO AND3HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8651 LAYER M1 ;
  END Z
END AND3HD2XHT

MACRO AND3HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
END AND3HDLXHT

MACRO AND3HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END AND3HDMXHT

MACRO AND4HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.091 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.091 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.091 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.091 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.74905 LAYER M1 ;
  END Z
END AND4HD1XHT

MACRO AND4HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1859 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1859 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1859 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1859 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8651 LAYER M1 ;
  END Z
END AND4HD2XHT

MACRO AND4HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2556 LAYER M1 ;
  END Z
END AND4HDLXHT

MACRO AND4HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3834 LAYER M1 ;
  END Z
END AND4HDMXHT

MACRO ANTFIXHDHT
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.7744 LAYER M1 ;
  END Z
END ANTFIXHDHT

MACRO AOI211HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END AOI211HD1XHT

MACRO AOI211HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END AOI211HD2XHT

MACRO AOI211HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.66735 LAYER M1 ;
  END Z
END AOI211HDLXHT

MACRO AOI211HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END AOI211HDMXHT

MACRO AOI21B2HD1XHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
  END C
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.67715 LAYER M1 ;
  END Z
END AOI21B2HD1XHT

MACRO AOI21B2HD2XHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1209 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.4862 LAYER M1 ;
  END C
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1209 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.9949 LAYER M1 ;
  END Z
END AOI21B2HD2XHT

MACRO AOI21B2HDLXHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END C
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.31365 LAYER M1 ;
  END Z
END AOI21B2HDLXHT

MACRO AOI21B2HDMXHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1703 LAYER M1 ;
  END C
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4722 LAYER M1 ;
  END Z
END AOI21B2HDMXHT

MACRO AOI21HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8328 LAYER M1 ;
  END Z
END AOI21HD1XHT

MACRO AOI21HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END AOI21HD2XHT

MACRO AOI21HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.34755 LAYER M1 ;
  END Z
END AOI21HDLXHT

MACRO AOI21HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1885 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1885 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1703 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5163 LAYER M1 ;
  END Z
END AOI21HDMXHT

MACRO AOI21HDUXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0754 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2569 LAYER M1 ;
  END Z
END AOI21HDUXHT

MACRO AOI221HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END AOI221HD1XHT

MACRO AOI221HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END AOI221HD2XHT

MACRO AOI221HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8514 LAYER M1 ;
  END Z
END AOI221HDLXHT

MACRO AOI221HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1989 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3861 LAYER M1 ;
  END Z
END AOI221HDMXHT

MACRO AOI222HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END AOI222HD1XHT

MACRO AOI222HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END AOI222HD2XHT

MACRO AOI222HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.693 LAYER M1 ;
  END Z
END AOI222HDLXHT

MACRO AOI222HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.1625 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3915 LAYER M1 ;
  END Z
END AOI222HDMXHT

MACRO AOI22B2HD1XHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.73395 LAYER M1 ;
  END Z
END AOI22B2HD1XHT

MACRO AOI22B2HD2XHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1209 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1209 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.0725 LAYER M1 ;
  END Z
END AOI22B2HD2XHT

MACRO AOI22B2HDLXHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3105 LAYER M1 ;
  END Z
END AOI22B2HDLXHT

MACRO AOI22B2HDMXHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1885 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1885 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.454 LAYER M1 ;
  END Z
END AOI22B2HDMXHT

MACRO AOI22HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.99265 LAYER M1 ;
  END Z
END AOI22HD1XHT

MACRO AOI22HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END AOI22HD2XHT

MACRO AOI22HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.303 LAYER M1 ;
  END Z
END AOI22HDLXHT

MACRO AOI22HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.44475 LAYER M1 ;
  END Z
END AOI22HDMXHT

MACRO AOI22HDUXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2772 LAYER M1 ;
  END Z
END AOI22HDUXHT

MACRO AOI31HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.221 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8412 LAYER M1 ;
  END Z
END AOI31HD1XHT

MACRO AOI31HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1404 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END AOI31HD2XHT

MACRO AOI31HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1404 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.47585 LAYER M1 ;
  END Z
END AOI31HDLXHT

MACRO AOI31HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2119 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2119 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2119 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6502 LAYER M1 ;
  END Z
END AOI31HDMXHT

MACRO AOI32HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2392 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2392 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8187 LAYER M1 ;
  END Z
END AOI32HD1XHT

MACRO AOI32HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1326 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1326 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1326 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END AOI32HD2XHT

MACRO AOI32HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1326 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1326 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1326 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4008 LAYER M1 ;
  END Z
END AOI32HDLXHT

MACRO AOI32HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1807 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1807 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1807 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1599 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1599 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5472 LAYER M1 ;
  END Z
END AOI32HDMXHT

MACRO AOI33HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.26105 LAYER M1 ;
  END Z
END AOI33HD1XHT

MACRO AOI33HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END AOI33HD2XHT

MACRO AOI33HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.44205 LAYER M1 ;
  END Z
END AOI33HDLXHT

MACRO AOI33HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.69825 LAYER M1 ;
  END Z
END AOI33HDMXHT

MACRO BUFCLKHD10XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.689 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.1041 LAYER M1 ;
  END Z
END BUFCLKHD10XHT

MACRO BUFCLKHD12XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.689 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.90525 LAYER M1 ;
  END Z
END BUFCLKHD12XHT

MACRO BUFCLKHD14XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.9217 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.6075 LAYER M1 ;
  END Z
END BUFCLKHD14XHT

MACRO BUFCLKHD16XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.157 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  4.3139 LAYER M1 ;
  END Z
END BUFCLKHD16XHT

MACRO BUFCLKHD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5934 LAYER M1 ;
  END Z
END BUFCLKHD1XHT

MACRO BUFCLKHD20XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.521 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  7.3671 LAYER M1 ;
  END Z
END BUFCLKHD20XHT

MACRO BUFCLKHD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.7045 LAYER M1 ;
  END Z
END BUFCLKHD2XHT

MACRO BUFCLKHD30XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.6796 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  10.7733 LAYER M1 ;
  END Z
END BUFCLKHD30XHT

MACRO BUFCLKHD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.35835 LAYER M1 ;
  END Z
END BUFCLKHD3XHT

MACRO BUFCLKHD40XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  2.236 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  13.962 LAYER M1 ;
  END Z
END BUFCLKHD40XHT

MACRO BUFCLKHD4XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2236 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.43775 LAYER M1 ;
  END Z
END BUFCLKHD4XHT

MACRO BUFCLKHD5XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2236 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.0355 LAYER M1 ;
  END Z
END BUFCLKHD5XHT

MACRO BUFCLKHD6XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.3367 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.78875 LAYER M1 ;
  END Z
END BUFCLKHD6XHT

MACRO BUFCLKHD7XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.3367 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.1996 LAYER M1 ;
  END Z
END BUFCLKHD7XHT

MACRO BUFCLKHD80XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  4.5916 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  27.9403 LAYER M1 ;
  END Z
END BUFCLKHD80XHT

MACRO BUFCLKHD8XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4628 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.0508 LAYER M1 ;
  END Z
END BUFCLKHD8XHT

MACRO BUFCLKHDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.36225 LAYER M1 ;
  END Z
END BUFCLKHDLXHT

MACRO BUFCLKHDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4347 LAYER M1 ;
  END Z
END BUFCLKHDMXHT

MACRO BUFCLKHDUXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.091 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2775 LAYER M1 ;
  END Z
END BUFCLKHDUXHT

MACRO BUFHD12XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.0972 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  4.9374 LAYER M1 ;
  END Z
END BUFHD12XHT

MACRO BUFHD16XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.3715 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  6.5832 LAYER M1 ;
  END Z
END BUFHD16XHT

MACRO BUFHD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END BUFHD1XHT

MACRO BUFHD20XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.6458 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  8.229 LAYER M1 ;
  END Z
END BUFHD20XHT

MACRO BUFHD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1846 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END BUFHD2XHT

MACRO BUFHD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END BUFHD3XHT

MACRO BUFHD4XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.3653 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.6458 LAYER M1 ;
  END Z
END BUFHD4XHT

MACRO BUFHD5XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.3653 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.37375 LAYER M1 ;
  END Z
END BUFHD5XHT

MACRO BUFHD6XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4121 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.4687 LAYER M1 ;
  END Z
END BUFHD6XHT

MACRO BUFHD7XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.19665 LAYER M1 ;
  END Z
END BUFHD7XHT

MACRO BUFHD8XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.7306 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.2916 LAYER M1 ;
  END Z
END BUFHD8XHT

MACRO BUFHD8XSPGHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.7306 LAYER M1 ;
    AntennaGateArea  0.7306 LAYER M2 ;
    AntennaGateArea  0.7306 LAYER M3 ;
    AntennaGateArea  0.7306 LAYER M4 ;
    AntennaGateArea  0.7306 LAYER M5 ;
    AntennaGateArea  0.7306 LAYER M6 ;
    AntennaGateArea  0.7306 LAYER M7 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.2916 LAYER M1 ;
    AntennaDiffArea  3.2916 LAYER M2 ;
    AntennaDiffArea  3.2916 LAYER M3 ;
    AntennaDiffArea  3.2916 LAYER M4 ;
    AntennaDiffArea  3.2916 LAYER M5 ;
    AntennaDiffArea  3.2916 LAYER M6 ;
    AntennaDiffArea  3.2916 LAYER M7 ;
  END Z
END BUFHD8XSPGHT

MACRO BUFHDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
END BUFHDLXHT

MACRO BUFHDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END BUFHDMXHT

MACRO BUFHDUXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0624 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.216 LAYER M1 ;
  END Z
END BUFHDUXHT

MACRO BUFTSHD12XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.8229 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.6578 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  5.5704 LAYER M1 ;
  END Z
END BUFTSHD12XHT

MACRO BUFTSHD16XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.6458 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  1.0335 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  7.2162 LAYER M1 ;
  END Z
END BUFTSHD16XHT

MACRO BUFTSHD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2613 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6694 LAYER M1 ;
  END Z
END BUFTSHD1XHT

MACRO BUFTSHD20XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.9201 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  1.209 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  8.862 LAYER M1 ;
  END Z
END BUFTSHD20XHT

MACRO BUFTSHD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1924 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.034 LAYER M1 ;
  END Z
END BUFTSHD2XHT

MACRO BUFTSHD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.2349 LAYER M1 ;
  END Z
END BUFTSHD3XHT

MACRO BUFTSHD4XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4368 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.299 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.89385 LAYER M1 ;
  END Z
END BUFTSHD4XHT

MACRO BUFTSHD5XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4992 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.3432 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.37375 LAYER M1 ;
  END Z
END BUFTSHD5XHT

MACRO BUFTSHD6XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.3705 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.4687 LAYER M1 ;
  END Z
END BUFTSHD6XHT

MACRO BUFTSHD7XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.7488 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.442 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.19665 LAYER M1 ;
  END Z
END BUFTSHD7XHT

MACRO BUFTSHD8XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.8229 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.4186 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.9246 LAYER M1 ;
  END Z
END BUFTSHD8XHT

MACRO BUFTSHDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1443 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.40365 LAYER M1 ;
  END Z
END BUFTSHDLXHT

MACRO BUFTSHDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1703 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6072 LAYER M1 ;
  END Z
END BUFTSHDMXHT

MACRO BUFTSHDUXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0624 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.0884 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2275 LAYER M1 ;
  END Z
END BUFTSHDUXHT

MACRO DEL1HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.7042 LAYER M1 ;
  END Z
END DEL1HD1XHT

MACRO DEL1HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END DEL1HDMXHT

MACRO DEL1HDMXSPGHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
    AntennaGateArea  0.0936 LAYER M2 ;
    AntennaGateArea  0.0936 LAYER M3 ;
    AntennaGateArea  0.0936 LAYER M4 ;
    AntennaGateArea  0.0936 LAYER M5 ;
    AntennaGateArea  0.0936 LAYER M6 ;
    AntennaGateArea  0.0936 LAYER M7 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.35835 LAYER M1 ;
    AntennaDiffArea  0.35835 LAYER M2 ;
    AntennaDiffArea  0.35835 LAYER M3 ;
    AntennaDiffArea  0.35835 LAYER M4 ;
    AntennaDiffArea  0.35835 LAYER M5 ;
    AntennaDiffArea  0.35835 LAYER M6 ;
    AntennaDiffArea  0.35835 LAYER M7 ;
  END Z
END DEL1HDMXSPGHT

MACRO DEL2HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END DEL2HD1XHT

MACRO DEL2HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END DEL2HDMXHT

MACRO DEL2HDMXSPGHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
    AntennaGateArea  0.0936 LAYER M2 ;
    AntennaGateArea  0.0936 LAYER M3 ;
    AntennaGateArea  0.0936 LAYER M4 ;
    AntennaGateArea  0.0936 LAYER M5 ;
    AntennaGateArea  0.0936 LAYER M6 ;
    AntennaGateArea  0.0936 LAYER M7 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
    AntennaDiffArea  0.327 LAYER M2 ;
    AntennaDiffArea  0.327 LAYER M3 ;
    AntennaDiffArea  0.327 LAYER M4 ;
    AntennaDiffArea  0.327 LAYER M5 ;
    AntennaDiffArea  0.327 LAYER M6 ;
    AntennaDiffArea  0.327 LAYER M7 ;
  END Z
END DEL2HDMXSPGHT

MACRO DEL3HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END DEL3HD1XHT

MACRO DEL3HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END DEL3HDMXHT

MACRO DEL4HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END DEL4HD1XHT

MACRO DEL4HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END DEL4HDMXHT

MACRO DEL4HDMXSPGHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
    AntennaGateArea  0.0936 LAYER M2 ;
    AntennaGateArea  0.0936 LAYER M3 ;
    AntennaGateArea  0.0936 LAYER M4 ;
    AntennaGateArea  0.0936 LAYER M5 ;
    AntennaGateArea  0.0936 LAYER M6 ;
    AntennaGateArea  0.0936 LAYER M7 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
    AntennaDiffArea  0.327 LAYER M2 ;
    AntennaDiffArea  0.327 LAYER M3 ;
    AntennaDiffArea  0.327 LAYER M4 ;
    AntennaDiffArea  0.327 LAYER M5 ;
    AntennaDiffArea  0.327 LAYER M6 ;
    AntennaDiffArea  0.327 LAYER M7 ;
  END Z
END DEL4HDMXSPGHT

MACRO FAHD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4368 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.3211 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END S
  PIN CI
    #DIRECTION INPUT ;
    AntennaGateArea  0.2886 LAYER M1 ;
  END CI
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5845 LAYER M1 ;
  END CO
END FAHD1XHT

MACRO FAHD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.4823 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END S
  PIN CI
    #DIRECTION INPUT ;
    AntennaGateArea  0.3939 LAYER M1 ;
  END CI
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END CO
END FAHD2XHT

MACRO FAHDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.3744 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.3211 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END S
  PIN CI
    #DIRECTION INPUT ;
    AntennaGateArea  0.2626 LAYER M1 ;
  END CI
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.261 LAYER M1 ;
  END CO
END FAHDLXHT

MACRO FAHDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.3744 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.3211 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.36225 LAYER M1 ;
  END S
  PIN CI
    #DIRECTION INPUT ;
    AntennaGateArea  0.2626 LAYER M1 ;
  END CI
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.38115 LAYER M1 ;
  END CO
END FAHDMXHT

MACRO FAHDUXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.216 LAYER M1 ;
  END S
  PIN CI
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END CI
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.216 LAYER M1 ;
  END CO
END FAHDUXHT

MACRO FAHHD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END S
  PIN CI
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END CI
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.73985 LAYER M1 ;
  END CO
END FAHHD1XHT

MACRO FAHHD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1651 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.3029 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END S
  PIN CI
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END CI
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END CO
END FAHHD2XHT

MACRO FAHHDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2499 LAYER M1 ;
  END S
  PIN CI
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END CI
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.255 LAYER M1 ;
  END CO
END FAHHDLXHT

MACRO FAHHDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3741 LAYER M1 ;
  END S
  PIN CI
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END CI
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3855 LAYER M1 ;
  END CO
END FAHHDMXHT

MACRO FFDCRHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
END FFDCRHD1XHT

MACRO FFDCRHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1144 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1144 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
END FFDCRHD2XHT

MACRO FFDCRHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.24 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.052 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.052 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
END FFDCRHDLXHT

MACRO FFDCRHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.33 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0637 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0637 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
END FFDCRHDMXHT

MACRO FFDHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
END FFDHD1XHT

MACRO FFDHD1XSPGHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
    AntennaDiffArea  0.72795 LAYER M2 ;
    AntennaDiffArea  0.72795 LAYER M3 ;
    AntennaDiffArea  0.72795 LAYER M4 ;
    AntennaDiffArea  0.72795 LAYER M5 ;
    AntennaDiffArea  0.72795 LAYER M6 ;
    AntennaDiffArea  0.72795 LAYER M7 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
    AntennaDiffArea  0.72795 LAYER M2 ;
    AntennaDiffArea  0.72795 LAYER M3 ;
    AntennaDiffArea  0.72795 LAYER M4 ;
    AntennaDiffArea  0.72795 LAYER M5 ;
    AntennaDiffArea  0.72795 LAYER M6 ;
    AntennaDiffArea  0.72795 LAYER M7 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
    AntennaGateArea  0.117 LAYER M2 ;
    AntennaGateArea  0.117 LAYER M3 ;
    AntennaGateArea  0.117 LAYER M4 ;
    AntennaGateArea  0.117 LAYER M5 ;
    AntennaGateArea  0.117 LAYER M6 ;
    AntennaGateArea  0.117 LAYER M7 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
    AntennaGateArea  0.078 LAYER M2 ;
    AntennaGateArea  0.078 LAYER M3 ;
    AntennaGateArea  0.078 LAYER M4 ;
    AntennaGateArea  0.078 LAYER M5 ;
    AntennaGateArea  0.078 LAYER M6 ;
    AntennaGateArea  0.078 LAYER M7 ;
  END CK
END FFDHD1XSPGHT

MACRO FFDHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
END FFDHD2XHT

MACRO FFDHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
END FFDHDLXHT

MACRO FFDHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
END FFDHDMXHT

MACRO FFDHQHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
END FFDHQHD1XHT

MACRO FFDHQHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
END FFDHQHD2XHT

MACRO FFDHQHD3XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
END FFDHQHD3XHT

MACRO FFDHQHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
END FFDHQHDMXHT

MACRO FFDNHD1XHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
END FFDNHD1XHT

MACRO FFDNHD2XHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
END FFDNHD2XHT

MACRO FFDNHDLXHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.065 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
END FFDNHDLXHT

MACRO FFDNHDMXHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
END FFDNHDMXHT

MACRO FFDNRHD1XHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
END FFDNRHD1XHT

MACRO FFDNRHD2XHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
END FFDNRHD2XHT

MACRO FFDNRHDLXHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.065 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
END FFDNRHDLXHT

MACRO FFDNRHDMXHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
END FFDNRHDMXHT

MACRO FFDNSHD1XHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFDNSHD1XHT

MACRO FFDNSHD2XHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3094 LAYER M1 ;
  END SN
END FFDNSHD2XHT

MACRO FFDNSHDLXHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.065 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFDNSHDLXHT

MACRO FFDNSHDMXHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFDNSHDMXHT

MACRO FFDNSRHD1XHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6814 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6168 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFDNSRHD1XHT

MACRO FFDNSRHD2XHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.338 LAYER M1 ;
  END SN
END FFDNSRHD2XHT

MACRO FFDNSRHDLXHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.065 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFDNSRHDLXHT

MACRO FFDNSRHDMXHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFDNSRHDMXHT

MACRO FFDQHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
END FFDQHD1XHT

MACRO FFDQHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
END FFDQHD2XHT

MACRO FFDQHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.27255 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
END FFDQHDLXHT

MACRO FFDQHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
END FFDQHDMXHT

MACRO FFDQRHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
END FFDQRHD1XHT

MACRO FFDQRHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
END FFDQRHD2XHT

MACRO FFDQRHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
END FFDQRHDLXHT

MACRO FFDQRHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
END FFDQRHDMXHT

MACRO FFDQSHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1859 LAYER M1 ;
  END SN
END FFDQSHD1XHT

MACRO FFDQSHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2405 LAYER M1 ;
  END SN
END FFDQSHD2XHT

MACRO FFDQSHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFDQSHDLXHT

MACRO FFDQSHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFDQSHDMXHT

MACRO FFDQSRHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1859 LAYER M1 ;
  END SN
END FFDQSRHD1XHT

MACRO FFDQSRHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2405 LAYER M1 ;
  END SN
END FFDQSRHD2XHT

MACRO FFDQSRHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFDQSRHDLXHT

MACRO FFDQSRHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFDQSRHDMXHT

MACRO FFDRHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
END FFDRHD1XHT

MACRO FFDRHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
END FFDRHD2XHT

MACRO FFDRHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
END FFDRHDLXHT

MACRO FFDRHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
END FFDRHDMXHT

MACRO FFDRHQHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
END FFDRHQHD1XHT

MACRO FFDRHQHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1755 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1404 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
END FFDRHQHD2XHT

MACRO FFDRHQHD3XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.5043 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2145 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
END FFDRHQHD3XHT

MACRO FFDRHQHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
END FFDRHQHDMXHT

MACRO FFDSHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFDSHD1XHT

MACRO FFDSHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3094 LAYER M1 ;
  END SN
END FFDSHD2XHT

MACRO FFDSHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFDSHDLXHT

MACRO FFDSHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFDSHDMXHT

MACRO FFDSHQHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2574 LAYER M1 ;
  END SN
END FFDSHQHD1XHT

MACRO FFDSHQHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.4559 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1755 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3198 LAYER M1 ;
  END SN
END FFDSHQHD2XHT

MACRO FFDSHQHD3XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2145 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3783 LAYER M1 ;
  END SN
END FFDSHQHD3XHT

MACRO FFDSHQHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFDSHQHDMXHT

MACRO FFDSRHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.70515 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.70515 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFDSRHD1XHT

MACRO FFDSRHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.338 LAYER M1 ;
  END SN
END FFDSRHD2XHT

MACRO FFDSRHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFDSRHDLXHT

MACRO FFDSRHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.35835 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.35835 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFDSRHDMXHT

MACRO FFDSRHQHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
  END SN
END FFDSRHQHD1XHT

MACRO FFDSRHQHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1755 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1404 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3198 LAYER M1 ;
  END SN
END FFDSRHQHD2XHT

MACRO FFDSRHQHD3XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2145 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3783 LAYER M1 ;
  END SN
END FFDSRHQHD3XHT

MACRO FFDSRHQHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3945 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.208 LAYER M1 ;
  END SN
END FFDSRHQHDMXHT

MACRO FFEDCRHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
END FFEDCRHD1XHT

MACRO FFEDCRHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
END FFEDCRHD2XHT

MACRO FFEDCRHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END E
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
END FFEDCRHDLXHT

MACRO FFEDCRHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3945 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1794 LAYER M1 ;
  END E
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
END FFEDCRHDMXHT

MACRO FFEDHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.7042 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
END FFEDHD1XHT

MACRO FFEDHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.2659 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
END FFEDHD2XHT

MACRO FFEDHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1794 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
END FFEDHDLXHT

MACRO FFEDHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
END FFEDHDMXHT

MACRO FFEDHQHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
END FFEDHQHD1XHT

MACRO FFEDHQHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.234 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.3276 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
END FFEDHQHD2XHT

MACRO FFEDHQHD3XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2756 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.3692 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
END FFEDHQHD3XHT

MACRO FFEDHQHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.52095 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
END FFEDHQHDMXHT

MACRO FFEDQHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
END FFEDQHD1XHT

MACRO FFEDQHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
END FFEDQHD2XHT

MACRO FFEDQHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
END FFEDQHDLXHT

MACRO FFEDQHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1794 LAYER M1 ;
  END E
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
END FFEDQHDMXHT

MACRO FFSDCRHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSDCRHD1XHT

MACRO FFSDCRHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSDCRHD2XHT

MACRO FFSDCRHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.169 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0689 LAYER M1 ;
  END TI
END FFSDCRHDLXHT

MACRO FFSDCRHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1144 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1144 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1846 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0689 LAYER M1 ;
  END TI
END FFSDCRHDMXHT

MACRO FFSDHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDHD1XHT

MACRO FFSDHD1XSPGHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
    AntennaDiffArea  0.72795 LAYER M2 ;
    AntennaDiffArea  0.72795 LAYER M3 ;
    AntennaDiffArea  0.72795 LAYER M4 ;
    AntennaDiffArea  0.72795 LAYER M5 ;
    AntennaDiffArea  0.72795 LAYER M6 ;
    AntennaDiffArea  0.72795 LAYER M7 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
    AntennaDiffArea  0.72795 LAYER M2 ;
    AntennaDiffArea  0.72795 LAYER M3 ;
    AntennaDiffArea  0.72795 LAYER M4 ;
    AntennaDiffArea  0.72795 LAYER M5 ;
    AntennaDiffArea  0.72795 LAYER M6 ;
    AntennaDiffArea  0.72795 LAYER M7 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
    AntennaGateArea  0.156 LAYER M2 ;
    AntennaGateArea  0.156 LAYER M3 ;
    AntennaGateArea  0.156 LAYER M4 ;
    AntennaGateArea  0.156 LAYER M5 ;
    AntennaGateArea  0.156 LAYER M6 ;
    AntennaGateArea  0.156 LAYER M7 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
    AntennaGateArea  0.2366 LAYER M2 ;
    AntennaGateArea  0.2366 LAYER M3 ;
    AntennaGateArea  0.2366 LAYER M4 ;
    AntennaGateArea  0.2366 LAYER M5 ;
    AntennaGateArea  0.2366 LAYER M6 ;
    AntennaGateArea  0.2366 LAYER M7 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
    AntennaGateArea  0.078 LAYER M2 ;
    AntennaGateArea  0.078 LAYER M3 ;
    AntennaGateArea  0.078 LAYER M4 ;
    AntennaGateArea  0.078 LAYER M5 ;
    AntennaGateArea  0.078 LAYER M6 ;
    AntennaGateArea  0.078 LAYER M7 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
    AntennaGateArea  0.117 LAYER M2 ;
    AntennaGateArea  0.117 LAYER M3 ;
    AntennaGateArea  0.117 LAYER M4 ;
    AntennaGateArea  0.117 LAYER M5 ;
    AntennaGateArea  0.117 LAYER M6 ;
    AntennaGateArea  0.117 LAYER M7 ;
  END TI
END FFSDHD1XSPGHT

MACRO FFSDHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDHD2XHT

MACRO FFSDHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
END FFSDHDLXHT

MACRO FFSDHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
END FFSDHDMXHT

MACRO FFSDHQHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDHQHD1XHT

MACRO FFSDHQHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.234 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2886 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDHQHD2XHT

MACRO FFSDHQHD3XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2925 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDHQHD3XHT

MACRO FFSDHQHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4752 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDHQHDMXHT

MACRO FFSDNHD1XHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDNHD1XHT

MACRO FFSDNHD2XHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDNHD2XHT

MACRO FFSDNHDLXHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.065 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
END FFSDNHDLXHT

MACRO FFSDNHDMXHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
END FFSDNHDMXHT

MACRO FFSDNRHD1XHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.70515 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDNRHD1XHT

MACRO FFSDNRHD2XHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDNRHD2XHT

MACRO FFSDNRHDLXHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.065 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
END FFSDNRHDLXHT

MACRO FFSDNRHDMXHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
END FFSDNRHDMXHT

MACRO FFSDNSHD1XHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFSDNSHD1XHT

MACRO FFSDNSHD2XHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3094 LAYER M1 ;
  END SN
END FFSDNSHD2XHT

MACRO FFSDNSHDLXHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.065 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFSDNSHDLXHT

MACRO FFSDNSHDMXHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFSDNSHDMXHT

MACRO FFSDNSRHD1XHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6814 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6168 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFSDNSRHD1XHT

MACRO FFSDNSRHD2XHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.338 LAYER M1 ;
  END SN
END FFSDNSRHD2XHT

MACRO FFSDNSRHDLXHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.065 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFSDNSRHDLXHT

MACRO FFSDNSRHDMXHT
  PIN CKN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END CKN
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFSDNSRHDMXHT

MACRO FFSDQHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDQHD1XHT

MACRO FFSDQHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDQHD2XHT

MACRO FFSDQHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
END FFSDQHDLXHT

MACRO FFSDQHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
END FFSDQHDMXHT

MACRO FFSDQRHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDQRHD1XHT

MACRO FFSDQRHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDQRHD2XHT

MACRO FFSDQRHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
END FFSDQRHDLXHT

MACRO FFSDQRHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
END FFSDQRHDMXHT

MACRO FFSDQSHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1859 LAYER M1 ;
  END SN
END FFSDQSHD1XHT

MACRO FFSDQSHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2405 LAYER M1 ;
  END SN
END FFSDQSHD2XHT

MACRO FFSDQSHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2709 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFSDQSHDLXHT

MACRO FFSDQSHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFSDQSHDMXHT

MACRO FFSDQSRHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1859 LAYER M1 ;
  END SN
END FFSDQSRHD1XHT

MACRO FFSDQSRHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2405 LAYER M1 ;
  END SN
END FFSDQSRHD2XHT

MACRO FFSDQSRHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFSDQSRHDLXHT

MACRO FFSDQSRHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFSDQSRHDMXHT

MACRO FFSDRHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDRHD1XHT

MACRO FFSDRHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDRHD2XHT

MACRO FFSDRHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
END FFSDRHDLXHT

MACRO FFSDRHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
END FFSDRHDMXHT

MACRO FFSDRHQHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDRHQHD1XHT

MACRO FFSDRHQHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.234 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1404 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2886 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDRHQHD2XHT

MACRO FFSDRHQHD3XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2925 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDRHQHD3XHT

MACRO FFSDRHQHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSDRHQHDMXHT

MACRO FFSDSHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFSDSHD1XHT

MACRO FFSDSHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3094 LAYER M1 ;
  END SN
END FFSDSHD2XHT

MACRO FFSDSHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFSDSHDLXHT

MACRO FFSDSHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFSDSHDMXHT

MACRO FFSDSHQHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2574 LAYER M1 ;
  END SN
END FFSDSHQHD1XHT

MACRO FFSDSHQHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.234 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2886 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3198 LAYER M1 ;
  END SN
END FFSDSHQHD2XHT

MACRO FFSDSHQHD3XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2925 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3783 LAYER M1 ;
  END SN
END FFSDSHQHD3XHT

MACRO FFSDSHQHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFSDSHQHDMXHT

MACRO FFSDSRHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.70515 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.70515 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END SN
END FFSDSRHD1XHT

MACRO FFSDSRHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.338 LAYER M1 ;
  END SN
END FFSDSRHD2XHT

MACRO FFSDSRHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END SN
END FFSDSRHDLXHT

MACRO FFSDSRHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END SN
END FFSDSRHDMXHT

MACRO FFSDSRHQHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
  END SN
END FFSDSRHQHD1XHT

MACRO FFSDSRHQHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.234 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1404 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2886 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3198 LAYER M1 ;
  END SN
END FFSDSRHQHD2XHT

MACRO FFSDSRHQHD3XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.49955 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2925 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3783 LAYER M1 ;
  END SN
END FFSDSRHQHD3XHT

MACRO FFSDSRHQHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.208 LAYER M1 ;
  END SN
END FFSDSRHQHDMXHT

MACRO FFSEDCRHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSEDCRHD1XHT

MACRO FFSEDCRHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END TI
END FFSEDCRHD2XHT

MACRO FFSEDCRHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END E
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END TI
END FFSEDCRHDLXHT

MACRO FFSEDCRHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1794 LAYER M1 ;
  END E
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END TI
END FFSEDCRHDMXHT

MACRO FFSEDHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDHD1XHT

MACRO FFSEDHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDHD2XHT

MACRO FFSEDHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDHDLXHT

MACRO FFSEDHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.35835 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.35835 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1794 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDHDMXHT

MACRO FFSEDHQHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDHQHD1XHT

MACRO FFSEDHQHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDHQHD2XHT

MACRO FFSEDHQHD3XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.39 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDHQHD3XHT

MACRO FFSEDHQHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.52095 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.195 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDHQHDMXHT

MACRO FFSEDQHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDQHD1XHT

MACRO FFSEDQHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDQHD2XHT

MACRO FFSEDQHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.1742 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0468 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDQHDLXHT

MACRO FFSEDQHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1794 LAYER M1 ;
  END E
  PIN TE
    #DIRECTION INPUT ;
    AntennaGateArea  0.2002 LAYER M1 ;
  END TE
  PIN CK
    #DIRECTION INPUT ;
    AntennaGateArea  0.0572 LAYER M1 ;
  END CK
  PIN TI
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END TI
END FFSEDQHDMXHT

MACRO FILLER16HDHT
END FILLER16HDHT

MACRO FILLER1HDHT
END FILLER1HDHT

MACRO FILLER2HDHT
END FILLER2HDHT

MACRO FILLER32HDHT
END FILLER32HDHT

MACRO FILLER3HDHT
END FILLER3HDHT

MACRO FILLER4HDHT
END FILLER4HDHT

MACRO FILLER64HDHT
END FILLER64HDHT

MACRO FILLER6HDHT
END FILLER6HDHT

MACRO FILLER8HDHT
END FILLER8HDHT

MACRO FILLERC16HDHT
END FILLERC16HDHT

MACRO FILLERC1HDHT
END FILLERC1HDHT

MACRO FILLERC2HDHT
END FILLERC2HDHT

MACRO FILLERC32HDHT
END FILLERC32HDHT

MACRO FILLERC3HDHT
END FILLERC3HDHT

MACRO FILLERC4HDHT
END FILLERC4HDHT

MACRO FILLERC64HDHT
END FILLERC64HDHT

MACRO FILLERC6HDHT
END FILLERC6HDHT

MACRO FILLERC8HDHT
END FILLERC8HDHT

MACRO HAHD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1885 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END S
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END CO
END HAHD1XHT

MACRO HAHD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.3276 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.4108 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END S
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END CO
END HAHD2XHT

MACRO HAHDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1794 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2574 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END S
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END CO
END HAHDLXHT

MACRO HAHDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1794 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2574 LAYER M1 ;
  END B
  PIN S
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END S
  PIN CO
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END CO
END HAHDMXHT

MACRO HOLDHDHT
  PIN Z
    #DIRECTION INOUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
    AntennaDiffArea  0.32445 LAYER M1 ;
  END Z
END HOLDHDHT

MACRO INVCLKHD10XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.911 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.09885 LAYER M1 ;
  END Z
END INVCLKHD10XHT

MACRO INVCLKHD12XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  2.262 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.393 LAYER M1 ;
  END Z
END INVCLKHD12XHT

MACRO INVCLKHD14XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  2.7807 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  4.3834 LAYER M1 ;
  END Z
END INVCLKHD14XHT

MACRO INVCLKHD16XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  3.484 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  5.2326 LAYER M1 ;
  END Z
END INVCLKHD16XHT

MACRO INVCLKHD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2236 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5934 LAYER M1 ;
  END Z
END INVCLKHD1XHT

MACRO INVCLKHD20XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  4.537 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  6.8066 LAYER M1 ;
  END Z
END INVCLKHD20XHT

MACRO INVCLKHD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4498 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6747 LAYER M1 ;
  END Z
END INVCLKHD2XHT

MACRO INVCLKHD30XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.455 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  10.3545 LAYER M1 ;
  END Z
END INVCLKHD30XHT

MACRO INVCLKHD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.6838 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.2897 LAYER M1 ;
  END Z
END INVCLKHD3XHT

MACRO INVCLKHD40XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5642 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  14.0082 LAYER M1 ;
  END Z
END INVCLKHD40XHT

MACRO INVCLKHD4XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.9087 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.3636 LAYER M1 ;
  END Z
END INVCLKHD4XHT

MACRO INVCLKHD5XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.053 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.8225 LAYER M1 ;
  END Z
END INVCLKHD5XHT

MACRO INVCLKHD6XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.2324 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.8486 LAYER M1 ;
  END Z
END INVCLKHD6XHT

MACRO INVCLKHD7XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.417 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.2324 LAYER M1 ;
  END Z
END INVCLKHD7XHT

MACRO INVCLKHD80XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.1193 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  28.0111 LAYER M1 ;
  END Z
END INVCLKHD80XHT

MACRO INVCLKHD8XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.638 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.4659 LAYER M1 ;
  END Z
END INVCLKHD8XHT

MACRO INVCLKHDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.36225 LAYER M1 ;
  END Z
END INVCLKHDLXHT

MACRO INVCLKHDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4347 LAYER M1 ;
  END Z
END INVCLKHDMXHT

MACRO INVCLKHDUXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.091 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2775 LAYER M1 ;
  END Z
END INVCLKHDUXHT

MACRO INVHD12XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  4.9374 LAYER M1 ;
  END Z
END INVHD12XHT

MACRO INVHD16XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4875 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  6.5832 LAYER M1 ;
  END Z
END INVHD16XHT

MACRO INVHD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END INVHD1XHT

MACRO INVHD1XSPGHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
    AntennaGateArea  0.2743 LAYER M2 ;
    AntennaGateArea  0.2743 LAYER M3 ;
    AntennaGateArea  0.2743 LAYER M4 ;
    AntennaGateArea  0.2743 LAYER M5 ;
    AntennaGateArea  0.2743 LAYER M6 ;
    AntennaGateArea  0.2743 LAYER M7 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
    AntennaDiffArea  0.72795 LAYER M2 ;
    AntennaDiffArea  0.72795 LAYER M3 ;
    AntennaDiffArea  0.72795 LAYER M4 ;
    AntennaDiffArea  0.72795 LAYER M5 ;
    AntennaDiffArea  0.72795 LAYER M6 ;
    AntennaDiffArea  0.72795 LAYER M7 ;
  END Z
END INVHD1XSPGHT

MACRO INVHD20XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  8.862 LAYER M1 ;
  END Z
END INVHD20XHT

MACRO INVHD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END INVHD2XHT

MACRO INVHD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.8229 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END INVHD3XHT

MACRO INVHD4XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.0972 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.6458 LAYER M1 ;
  END Z
END INVHD4XHT

MACRO INVHD5XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.3715 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.37375 LAYER M1 ;
  END Z
END INVHD5XHT

MACRO INVHD6XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.6458 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.4687 LAYER M1 ;
  END Z
END INVHD6XHT

MACRO INVHD7XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  1.9201 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.19665 LAYER M1 ;
  END Z
END INVHD7XHT

MACRO INVHD8XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  2.1944 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.2916 LAYER M1 ;
  END Z
END INVHD8XHT

MACRO INVHDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
END INVHDLXHT

MACRO INVHDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1404 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END INVHDMXHT

MACRO INVHDPXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.247 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6555 LAYER M1 ;
  END Z
END INVHDPXHT

MACRO INVHDUXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0624 LAYER M1 ;
  END A
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2246 LAYER M1 ;
  END Z
END INVHDUXHT

MACRO INVODHD8XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN Z0
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z0
  PIN Z1
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z1
  PIN Z2
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z2
  PIN Z3
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z3
  PIN Z4
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z4
  PIN Z5
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z5
  PIN Z6
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z6
  PIN Z7
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z7
END INVODHD8XHT

MACRO INVTSHD12XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.6578 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  5.5704 LAYER M1 ;
  END Z
END INVTSHD12XHT

MACRO INVTSHD16XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  1.0335 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  7.2162 LAYER M1 ;
  END Z
END INVTSHD16XHT

MACRO INVTSHD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4459 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2587 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6694 LAYER M1 ;
  END Z
END INVTSHD1XHT

MACRO INVTSHD20XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  1.209 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  8.862 LAYER M1 ;
  END Z
END INVTSHD20XHT

MACRO INVTSHD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.8918 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.5174 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.3388 LAYER M1 ;
  END Z
END INVTSHD2XHT

MACRO INVTSHD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.2349 LAYER M1 ;
  END Z
END INVTSHD3XHT

MACRO INVTSHD4XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1495 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.299 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.89385 LAYER M1 ;
  END Z
END INVTSHD4XHT

MACRO INVTSHD5XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1677 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.3432 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.06505 LAYER M1 ;
  END Z
END INVTSHD5XHT

MACRO INVTSHD6XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1833 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.3705 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.74215 LAYER M1 ;
  END Z
END INVTSHD6XHT

MACRO INVTSHD7XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.442 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.88195 LAYER M1 ;
  END Z
END INVTSHD7XHT

MACRO INVTSHD8XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.4186 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  3.9246 LAYER M1 ;
  END Z
END INVTSHD8XHT

MACRO INVTSHDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1534 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1456 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4071 LAYER M1 ;
  END Z
END INVTSHDLXHT

MACRO INVTSHDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2288 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1703 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6072 LAYER M1 ;
  END Z
END INVTSHDMXHT

MACRO INVTSHDUXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1014 LAYER M1 ;
  END A
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.0962 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2889 LAYER M1 ;
  END Z
END INVTSHDUXHT

MACRO LATHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
END LATHD1XHT

MACRO LATHD1XSPGHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
    AntennaDiffArea  0.72795 LAYER M2 ;
    AntennaDiffArea  0.72795 LAYER M3 ;
    AntennaDiffArea  0.72795 LAYER M4 ;
    AntennaDiffArea  0.72795 LAYER M5 ;
    AntennaDiffArea  0.72795 LAYER M6 ;
    AntennaDiffArea  0.72795 LAYER M7 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
    AntennaDiffArea  0.72795 LAYER M2 ;
    AntennaDiffArea  0.72795 LAYER M3 ;
    AntennaDiffArea  0.72795 LAYER M4 ;
    AntennaDiffArea  0.72795 LAYER M5 ;
    AntennaDiffArea  0.72795 LAYER M6 ;
    AntennaDiffArea  0.72795 LAYER M7 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
    AntennaGateArea  0.156 LAYER M2 ;
    AntennaGateArea  0.156 LAYER M3 ;
    AntennaGateArea  0.156 LAYER M4 ;
    AntennaGateArea  0.156 LAYER M5 ;
    AntennaGateArea  0.156 LAYER M6 ;
    AntennaGateArea  0.156 LAYER M7 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
    AntennaGateArea  0.117 LAYER M2 ;
    AntennaGateArea  0.117 LAYER M3 ;
    AntennaGateArea  0.117 LAYER M4 ;
    AntennaGateArea  0.117 LAYER M5 ;
    AntennaGateArea  0.117 LAYER M6 ;
    AntennaGateArea  0.117 LAYER M7 ;
  END G
END LATHD1XSPGHT

MACRO LATHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2405 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
END LATHD2XHT

MACRO LATHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2442 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2589 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END G
END LATHDLXHT

MACRO LATHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END G
END LATHDMXHT

MACRO LATNHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
END LATNHD1XHT

MACRO LATNHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2405 LAYER M1 ;
  END D
END LATNHD2XHT

MACRO LATNHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
END LATNHDLXHT

MACRO LATNHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
END LATNHDMXHT

MACRO LATNRHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6396 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2288 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END RN
END LATNRHD1XHT

MACRO LATNRHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3523 LAYER M1 ;
  END RN
END LATNRHD2XHT

MACRO LATNRHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2376 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1508 LAYER M1 ;
  END RN
END LATNRHDLXHT

MACRO LATNRHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.34125 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2132 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2145 LAYER M1 ;
  END RN
END LATNRHDMXHT

MACRO LATNSHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.67285 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
  END D
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END LATNSHD1XHT

MACRO LATNSHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1261 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
  END D
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END SN
END LATNSHD2XHT

MACRO LATNSHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1885 LAYER M1 ;
  END D
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END LATNSHDLXHT

MACRO LATNSHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.35835 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2262 LAYER M1 ;
  END D
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END LATNSHDMXHT

MACRO LATNSRHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6168 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6814 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2652 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END SN
END LATNSRHD1XHT

MACRO LATNSRHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3523 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END SN
END LATNSRHD2XHT

MACRO LATNSRHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.221 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END LATNSRHDLXHT

MACRO LATNSRHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END Q
  PIN GN
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END GN
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END D
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2652 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END SN
END LATNSRHDMXHT

MACRO LATRHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6396 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2288 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END RN
END LATRHD1XHT

MACRO LATRHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3523 LAYER M1 ;
  END RN
END LATRHD2XHT

MACRO LATRHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END G
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1508 LAYER M1 ;
  END RN
END LATRHDLXHT

MACRO LATRHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.34125 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2132 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2145 LAYER M1 ;
  END RN
END LATRHDMXHT

MACRO LATSHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.67285 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END LATSHD1XHT

MACRO LATSHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END SN
END LATSHD2XHT

MACRO LATSHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1885 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END G
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END LATSHDLXHT

MACRO LATSHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.35835 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2262 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END LATSHDMXHT

MACRO LATSRHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6168 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6814 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2652 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END SN
END LATSRHD1XHT

MACRO LATSRHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.3523 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END SN
END LATSRHD2XHT

MACRO LATSRHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.237 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END G
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.221 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END LATSRHDLXHT

MACRO LATSRHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END QN
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END D
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.2652 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1378 LAYER M1 ;
  END SN
END LATSRHDMXHT

MACRO LATTSHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.3938 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.312 LAYER M1 ;
  END E
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
END LATTSHD1XHT

MACRO LATTSHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END E
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
END LATTSHD2XHT

MACRO LATTSHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.32515 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1456 LAYER M1 ;
  END E
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END G
END LATTSHDLXHT

MACRO LATTSHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4968 LAYER M1 ;
  END Q
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END E
  PIN G
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END G
END LATTSHDMXHT

MACRO MUX2CLKHD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5865 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END S0
END MUX2CLKHD1XHT

MACRO MUX2CLKHD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.69615 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2366 LAYER M1 ;
  END S0
END MUX2CLKHD2XHT

MACRO MUX2CLKHD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2197 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2197 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.30605 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.3133 LAYER M1 ;
  END S0
END MUX2CLKHD3XHT

MACRO MUX2CLKHD4XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.312 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.312 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.3701 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.4056 LAYER M1 ;
  END S0
END MUX2CLKHD4XHT

MACRO MUX2HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2184 LAYER M1 ;
  END S0
END MUX2HD1XHT

MACRO MUX2HD1XSPGHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
    AntennaGateArea  0.1248 LAYER M2 ;
    AntennaGateArea  0.1248 LAYER M3 ;
    AntennaGateArea  0.1248 LAYER M4 ;
    AntennaGateArea  0.1248 LAYER M5 ;
    AntennaGateArea  0.1248 LAYER M6 ;
    AntennaGateArea  0.1248 LAYER M7 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
    AntennaGateArea  0.1248 LAYER M2 ;
    AntennaGateArea  0.1248 LAYER M3 ;
    AntennaGateArea  0.1248 LAYER M4 ;
    AntennaGateArea  0.1248 LAYER M5 ;
    AntennaGateArea  0.1248 LAYER M6 ;
    AntennaGateArea  0.1248 LAYER M7 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
    AntennaDiffArea  0.72795 LAYER M2 ;
    AntennaDiffArea  0.72795 LAYER M3 ;
    AntennaDiffArea  0.72795 LAYER M4 ;
    AntennaDiffArea  0.72795 LAYER M5 ;
    AntennaDiffArea  0.72795 LAYER M6 ;
    AntennaDiffArea  0.72795 LAYER M7 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2184 LAYER M1 ;
    AntennaGateArea  0.2184 LAYER M2 ;
    AntennaGateArea  0.2184 LAYER M3 ;
    AntennaGateArea  0.2184 LAYER M4 ;
    AntennaGateArea  0.2184 LAYER M5 ;
    AntennaGateArea  0.2184 LAYER M6 ;
    AntennaGateArea  0.2184 LAYER M7 ;
  END S0
END MUX2HD1XSPGHT

MACRO MUX2HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.89675 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.3432 LAYER M1 ;
  END S0
END MUX2HD2XHT

MACRO MUX2HD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.3679 LAYER M1 ;
  END S0
END MUX2HD3XHT

MACRO MUX2HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S0
END MUX2HDLXHT

MACRO MUX2HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S0
END MUX2HDMXHT

MACRO MUX2HDUXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0624 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0624 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.461 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END S0
END MUX2HDUXHT

MACRO MUX4HD1XHT
  PIN S1
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S1
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6814 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END S0
END MUX4HD1XHT

MACRO MUX4HD2XHT
  PIN S1
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S1
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END S0
END MUX4HD2XHT

MACRO MUX4HDLXHT
  PIN S1
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S1
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END S0
END MUX4HDLXHT

MACRO MUX4HDMXHT
  PIN S1
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S1
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END S0
END MUX4HDMXHT

MACRO MUXI2HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S0
END MUXI2HD1XHT

MACRO MUXI2HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S0
END MUXI2HD2XHT

MACRO MUXI2HD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S0
END MUXI2HD3XHT

MACRO MUXI2HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S0
END MUXI2HDLXHT

MACRO MUXI2HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S0
END MUXI2HDMXHT

MACRO MUXI4HD1XHT
  PIN S1
    #DIRECTION INPUT ;
    AntennaGateArea  0.2184 LAYER M1 ;
  END S1
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END S0
END MUXI4HD1XHT

MACRO MUXI4HD2XHT
  PIN S1
    #DIRECTION INPUT ;
    AntennaGateArea  0.3432 LAYER M1 ;
  END S1
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.3198 LAYER M1 ;
  END S0
END MUXI4HD2XHT

MACRO MUXI4HDLXHT
  PIN S1
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S1
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END S0
END MUXI4HDLXHT

MACRO MUXI4HDMXHT
  PIN S1
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END S1
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
  PIN S0
    #DIRECTION INPUT ;
    AntennaGateArea  0.2808 LAYER M1 ;
  END S0
END MUXI4HDMXHT

MACRO NAND2B1HD1XHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.717 LAYER M1 ;
  END Z
END NAND2B1HD1XHT

MACRO NAND2B1HD2XHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.5044 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1404 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.17 LAYER M1 ;
  END Z
END NAND2B1HD2XHT

MACRO NAND2B1HDLXHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2439 LAYER M1 ;
  END Z
END NAND2B1HDLXHT

MACRO NAND2B1HDMXHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1508 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4067 LAYER M1 ;
  END Z
END NAND2B1HDMXHT

MACRO NAND2B1HDUXHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0624 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.318 LAYER M1 ;
  END Z
END NAND2B1HDUXHT

MACRO NAND2HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.0438 LAYER M1 ;
  END Z
END NAND2HD1XHT

MACRO NAND2HD1XSPGHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
    AntennaGateArea  0.2522 LAYER M2 ;
    AntennaGateArea  0.2522 LAYER M3 ;
    AntennaGateArea  0.2522 LAYER M4 ;
    AntennaGateArea  0.2522 LAYER M5 ;
    AntennaGateArea  0.2522 LAYER M6 ;
    AntennaGateArea  0.2522 LAYER M7 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
    AntennaGateArea  0.2522 LAYER M2 ;
    AntennaGateArea  0.2522 LAYER M3 ;
    AntennaGateArea  0.2522 LAYER M4 ;
    AntennaGateArea  0.2522 LAYER M5 ;
    AntennaGateArea  0.2522 LAYER M6 ;
    AntennaGateArea  0.2522 LAYER M7 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.0186 LAYER M1 ;
    AntennaDiffArea  1.0186 LAYER M2 ;
    AntennaDiffArea  1.0186 LAYER M3 ;
    AntennaDiffArea  1.0186 LAYER M4 ;
    AntennaDiffArea  1.0186 LAYER M5 ;
    AntennaDiffArea  1.0186 LAYER M6 ;
    AntennaDiffArea  1.0186 LAYER M7 ;
  END Z
END NAND2HD1XSPGHT

MACRO NAND2HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5044 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.5044 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.17 LAYER M1 ;
  END Z
END NAND2HD2XHT

MACRO NAND2HD2XSPGHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.5044 LAYER M1 ;
    AntennaGateArea  0.5044 LAYER M2 ;
    AntennaGateArea  0.5044 LAYER M3 ;
    AntennaGateArea  0.5044 LAYER M4 ;
    AntennaGateArea  0.5044 LAYER M5 ;
    AntennaGateArea  0.5044 LAYER M6 ;
    AntennaGateArea  0.5044 LAYER M7 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.5044 LAYER M1 ;
    AntennaGateArea  0.5044 LAYER M2 ;
    AntennaGateArea  0.5044 LAYER M3 ;
    AntennaGateArea  0.5044 LAYER M4 ;
    AntennaGateArea  0.5044 LAYER M5 ;
    AntennaGateArea  0.5044 LAYER M6 ;
    AntennaGateArea  0.5044 LAYER M7 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.17 LAYER M1 ;
    AntennaDiffArea  1.17 LAYER M2 ;
    AntennaDiffArea  1.17 LAYER M3 ;
    AntennaDiffArea  1.17 LAYER M4 ;
    AntennaDiffArea  1.17 LAYER M5 ;
    AntennaDiffArea  1.17 LAYER M6 ;
    AntennaDiffArea  1.17 LAYER M7 ;
  END Z
END NAND2HD2XSPGHT

MACRO NAND2HD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.7566 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.7566 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  2.205 LAYER M1 ;
  END Z
END NAND2HD3XHT

MACRO NAND2HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2439 LAYER M1 ;
  END Z
END NAND2HDLXHT

MACRO NAND2HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1508 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1508 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.42855 LAYER M1 ;
  END Z
END NAND2HDMXHT

MACRO NAND2HDUXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0676 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0676 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.321 LAYER M1 ;
  END Z
END NAND2HDUXHT

MACRO NAND2ODHDHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z
END NAND2ODHDHT

MACRO NAND3B1HD1XHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2288 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2288 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.9548 LAYER M1 ;
  END Z
END NAND3B1HD1XHT

MACRO NAND3B1HD2XHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NAND3B1HD2XHT

MACRO NAND3B1HDLXHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4705 LAYER M1 ;
  END Z
END NAND3B1HDLXHT

MACRO NAND3B1HDMXHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.78895 LAYER M1 ;
  END Z
END NAND3B1HDMXHT

MACRO NAND3HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2288 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2288 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2288 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.9352 LAYER M1 ;
  END Z
END NAND3HD1XHT

MACRO NAND3HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NAND3HD2XHT

MACRO NAND3HD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END NAND3HD3XHT

MACRO NAND3HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3285 LAYER M1 ;
  END Z
END NAND3HDLXHT

MACRO NAND3HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.68985 LAYER M1 ;
  END Z
END NAND3HDMXHT

MACRO NAND3ODHDHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.078 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3036 LAYER M1 ;
  END Z
END NAND3ODHDHT

MACRO NAND4B1HD1XHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END NAND4B1HD1XHT

MACRO NAND4B1HD2XHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NAND4B1HD2XHT

MACRO NAND4B1HDLXHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.471 LAYER M1 ;
  END Z
END NAND4B1HDLXHT

MACRO NAND4B1HDMXHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.7329 LAYER M1 ;
  END Z
END NAND4B1HDMXHT

MACRO NAND4B2HD1XHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END NAND4B2HD1XHT

MACRO NAND4B2HD2XHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NAND4B2HD2XHT

MACRO NAND4B2HDLXHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.345 LAYER M1 ;
  END Z
END NAND4B2HDLXHT

MACRO NAND4B2HDMXHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.7272 LAYER M1 ;
  END Z
END NAND4B2HDMXHT

MACRO NAND4HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END NAND4HD1XHT

MACRO NAND4HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NAND4HD2XHT

MACRO NAND4HD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END NAND4HD3XHT

MACRO NAND4HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0819 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.34785 LAYER M1 ;
  END Z
END NAND4HDLXHT

MACRO NAND4HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6949 LAYER M1 ;
  END Z
END NAND4HDMXHT

MACRO NOR2B1HD1XHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.67395 LAYER M1 ;
  END Z
END NOR2B1HD1XHT

MACRO NOR2B1HD2XHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.4862 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1404 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.9789 LAYER M1 ;
  END Z
END NOR2B1HD2XHT

MACRO NOR2B1HDLXHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3165 LAYER M1 ;
  END Z
END NOR2B1HDLXHT

MACRO NOR2B1HDMXHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1703 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4765 LAYER M1 ;
  END Z
END NOR2B1HDMXHT

MACRO NOR2B1HDUXHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0754 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0624 LAYER M1 ;
  END AN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2511 LAYER M1 ;
  END Z
END NOR2B1HDUXHT

MACRO NOR2HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6801 LAYER M1 ;
  END Z
END NOR2HD1XHT

MACRO NOR2HD1XSPGHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
    AntennaGateArea  0.2431 LAYER M2 ;
    AntennaGateArea  0.2431 LAYER M3 ;
    AntennaGateArea  0.2431 LAYER M4 ;
    AntennaGateArea  0.2431 LAYER M5 ;
    AntennaGateArea  0.2431 LAYER M6 ;
    AntennaGateArea  0.2431 LAYER M7 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2431 LAYER M1 ;
    AntennaGateArea  0.2431 LAYER M2 ;
    AntennaGateArea  0.2431 LAYER M3 ;
    AntennaGateArea  0.2431 LAYER M4 ;
    AntennaGateArea  0.2431 LAYER M5 ;
    AntennaGateArea  0.2431 LAYER M6 ;
    AntennaGateArea  0.2431 LAYER M7 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6801 LAYER M1 ;
    AntennaDiffArea  0.6801 LAYER M2 ;
    AntennaDiffArea  0.6801 LAYER M3 ;
    AntennaDiffArea  0.6801 LAYER M4 ;
    AntennaDiffArea  0.6801 LAYER M5 ;
    AntennaDiffArea  0.6801 LAYER M6 ;
    AntennaDiffArea  0.6801 LAYER M7 ;
  END Z
END NOR2HD1XSPGHT

MACRO NOR2HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4862 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.4862 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.0286 LAYER M1 ;
  END Z
END NOR2HD2XHT

MACRO NOR2HD2XSPGHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.4862 LAYER M1 ;
    AntennaGateArea  0.4862 LAYER M2 ;
    AntennaGateArea  0.4862 LAYER M3 ;
    AntennaGateArea  0.4862 LAYER M4 ;
    AntennaGateArea  0.4862 LAYER M5 ;
    AntennaGateArea  0.4862 LAYER M6 ;
    AntennaGateArea  0.4862 LAYER M7 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.4862 LAYER M1 ;
    AntennaGateArea  0.4862 LAYER M2 ;
    AntennaGateArea  0.4862 LAYER M3 ;
    AntennaGateArea  0.4862 LAYER M4 ;
    AntennaGateArea  0.4862 LAYER M5 ;
    AntennaGateArea  0.4862 LAYER M6 ;
    AntennaGateArea  0.4862 LAYER M7 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.0286 LAYER M1 ;
    AntennaDiffArea  1.0286 LAYER M2 ;
    AntennaDiffArea  1.0286 LAYER M3 ;
    AntennaDiffArea  1.0286 LAYER M4 ;
    AntennaDiffArea  1.0286 LAYER M5 ;
    AntennaDiffArea  1.0286 LAYER M6 ;
    AntennaDiffArea  1.0286 LAYER M7 ;
  END Z
END NOR2HD2XSPGHT

MACRO NOR2HD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.7332 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.7332 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.87255 LAYER M1 ;
  END Z
END NOR2HD3XHT

MACRO NOR2HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.31365 LAYER M1 ;
  END Z
END NOR2HDLXHT

MACRO NOR2HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1703 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1703 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4722 LAYER M1 ;
  END Z
END NOR2HDMXHT

MACRO NOR2HDUXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0754 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0754 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4029 LAYER M1 ;
  END Z
END NOR2HDUXHT

MACRO NOR3B1HD1XHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.83595 LAYER M1 ;
  END Z
END NOR3B1HD1XHT

MACRO NOR3B1HD2XHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NOR3B1HD2XHT

MACRO NOR3B1HDLXHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5943 LAYER M1 ;
  END Z
END NOR3B1HDLXHT

MACRO NOR3B1HDMXHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.65805 LAYER M1 ;
  END Z
END NOR3B1HDMXHT

MACRO NOR3HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.83595 LAYER M1 ;
  END Z
END NOR3HD1XHT

MACRO NOR3HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NOR3HD2XHT

MACRO NOR3HD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END NOR3HD3XHT

MACRO NOR3HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4463 LAYER M1 ;
  END Z
END NOR3HDLXHT

MACRO NOR3HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6723 LAYER M1 ;
  END Z
END NOR3HDMXHT

MACRO NOR4B1HD1XHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END NOR4B1HD1XHT

MACRO NOR4B1HD2XHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NOR4B1HD2XHT

MACRO NOR4B1HDLXHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.62025 LAYER M1 ;
  END Z
END NOR4B1HDLXHT

MACRO NOR4B1HDMXHT
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END B
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.93295 LAYER M1 ;
  END Z
END NOR4B1HDMXHT

MACRO NOR4B2HD1XHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.7042 LAYER M1 ;
  END Z
END NOR4B2HD1XHT

MACRO NOR4B2HD2XHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NOR4B2HD2XHT

MACRO NOR4B2HDLXHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.49275 LAYER M1 ;
  END Z
END NOR4B2HDLXHT

MACRO NOR4B2HDMXHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.74085 LAYER M1 ;
  END Z
END NOR4B2HDMXHT

MACRO NOR4HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END NOR4HD1XHT

MACRO NOR4HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END NOR4HD2XHT

MACRO NOR4HD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END NOR4HD3XHT

MACRO NOR4HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.53025 LAYER M1 ;
  END Z
END NOR4HDLXHT

MACRO NOR4HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.79715 LAYER M1 ;
  END Z
END NOR4HDMXHT

MACRO OAI211HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1976 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1976 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.999 LAYER M1 ;
  END Z
END OAI211HD1XHT

MACRO OAI211HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0897 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0897 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OAI211HD2XHT

MACRO OAI211HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0897 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0897 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4503 LAYER M1 ;
  END Z
END OAI211HDLXHT

MACRO OAI211HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1274 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1274 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.63945 LAYER M1 ;
  END Z
END OAI211HDMXHT

MACRO OAI21B2HD1XHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2522 LAYER M1 ;
  END C
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.717 LAYER M1 ;
  END Z
END OAI21B2HD1XHT

MACRO OAI21B2HD2XHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1261 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.5044 LAYER M1 ;
  END C
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.1261 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.17 LAYER M1 ;
  END Z
END OAI21B2HD2XHT

MACRO OAI21B2HDLXHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END C
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2439 LAYER M1 ;
  END Z
END OAI21B2HDLXHT

MACRO OAI21B2HDMXHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1508 LAYER M1 ;
  END C
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4067 LAYER M1 ;
  END Z
END OAI21B2HDMXHT

MACRO OAI21HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2015 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8028 LAYER M1 ;
  END Z
END OAI21HD1XHT

MACRO OAI21HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1261 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1261 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OAI21HD2XHT

MACRO OAI21HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1261 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1261 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.36165 LAYER M1 ;
  END Z
END OAI21HDLXHT

MACRO OAI21HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2171 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2171 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1508 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6234 LAYER M1 ;
  END Z
END OAI21HDMXHT

MACRO OAI21HDUXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0702 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3588 LAYER M1 ;
  END Z
END OAI21HDUXHT

MACRO OAI221HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1976 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.041 LAYER M1 ;
  END Z
END OAI221HD1XHT

MACRO OAI221HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.0897 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OAI221HD2XHT

MACRO OAI221HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1222 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.0897 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.45255 LAYER M1 ;
  END Z
END OAI221HDLXHT

MACRO OAI221HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1729 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1274 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6423 LAYER M1 ;
  END Z
END OAI221HDMXHT

MACRO OAI222HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.2704 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.2795 LAYER M1 ;
  END Z
END OAI222HD1XHT

MACRO OAI222HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OAI222HD2XHT

MACRO OAI222HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.0949 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.54855 LAYER M1 ;
  END Z
END OAI222HDLXHT

MACRO OAI222HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.156 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.74135 LAYER M1 ;
  END Z
END OAI222HDMXHT

MACRO OAI22B2HD1XHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.7947 LAYER M1 ;
  END Z
END OAI22B2HD1XHT

MACRO OAI22B2HD2XHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.5486 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.5084 LAYER M1 ;
  END Z
END OAI22B2HD2XHT

MACRO OAI22B2HDLXHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3819 LAYER M1 ;
  END Z
END OAI22B2HDLXHT

MACRO OAI22B2HDMXHT
  PIN AN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END AN
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1937 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1937 LAYER M1 ;
  END D
  PIN BN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0858 LAYER M1 ;
  END BN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5196 LAYER M1 ;
  END Z
END OAI22B2HDMXHT

MACRO OAI22HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.91515 LAYER M1 ;
  END Z
END OAI22HD1XHT

MACRO OAI22HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OAI22HD2XHT

MACRO OAI22HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0975 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2925 LAYER M1 ;
  END Z
END OAI22HDLXHT

MACRO OAI22HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.143 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.429 LAYER M1 ;
  END Z
END OAI22HDMXHT

MACRO OAI22HDUXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0832 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2772 LAYER M1 ;
  END Z
END OAI22HDUXHT

MACRO OAI31HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0806 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END OAI31HD1XHT

MACRO OAI31HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0806 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OAI31HD2XHT

MACRO OAI31HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.0806 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4587 LAYER M1 ;
  END Z
END OAI31HDLXHT

MACRO OAI31HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.104 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.58965 LAYER M1 ;
  END Z
END OAI31HDMXHT

MACRO OAI32HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END OAI32HD1XHT

MACRO OAI32HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OAI32HD2XHT

MACRO OAI32HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.117 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.4932 LAYER M1 ;
  END Z
END OAI32HDLXHT

MACRO OAI32HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1495 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1495 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.63345 LAYER M1 ;
  END Z
END OAI32HDMXHT

MACRO OAI33HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END OAI33HD1XHT

MACRO OAI33HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OAI33HD2XHT

MACRO OAI33HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.1638 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6237 LAYER M1 ;
  END Z
END OAI33HDLXHT

MACRO OAI33HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END D
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END E
  PIN F
    #DIRECTION INPUT ;
    AntennaGateArea  0.2106 LAYER M1 ;
  END F
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.80325 LAYER M1 ;
  END Z
END OAI33HDMXHT

MACRO OR2HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72315 LAYER M1 ;
  END Z
END OR2HD1XHT

MACRO OR2HD1XSPGHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
    AntennaGateArea  0.1131 LAYER M2 ;
    AntennaGateArea  0.1131 LAYER M3 ;
    AntennaGateArea  0.1131 LAYER M4 ;
    AntennaGateArea  0.1131 LAYER M5 ;
    AntennaGateArea  0.1131 LAYER M6 ;
    AntennaGateArea  0.1131 LAYER M7 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
    AntennaGateArea  0.1131 LAYER M2 ;
    AntennaGateArea  0.1131 LAYER M3 ;
    AntennaGateArea  0.1131 LAYER M4 ;
    AntennaGateArea  0.1131 LAYER M5 ;
    AntennaGateArea  0.1131 LAYER M6 ;
    AntennaGateArea  0.1131 LAYER M7 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72315 LAYER M1 ;
    AntennaDiffArea  0.72315 LAYER M2 ;
    AntennaDiffArea  0.72315 LAYER M3 ;
    AntennaDiffArea  0.72315 LAYER M4 ;
    AntennaDiffArea  0.72315 LAYER M5 ;
    AntennaDiffArea  0.72315 LAYER M6 ;
    AntennaDiffArea  0.72315 LAYER M7 ;
  END Z
END OR2HD1XSPGHT

MACRO OR2HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2262 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2262 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OR2HD2XHT

MACRO OR2HD2XSPGHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2262 LAYER M1 ;
    AntennaGateArea  0.2262 LAYER M2 ;
    AntennaGateArea  0.2262 LAYER M3 ;
    AntennaGateArea  0.2262 LAYER M4 ;
    AntennaGateArea  0.2262 LAYER M5 ;
    AntennaGateArea  0.2262 LAYER M6 ;
    AntennaGateArea  0.2262 LAYER M7 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2262 LAYER M1 ;
    AntennaGateArea  0.2262 LAYER M2 ;
    AntennaGateArea  0.2262 LAYER M3 ;
    AntennaGateArea  0.2262 LAYER M4 ;
    AntennaGateArea  0.2262 LAYER M5 ;
    AntennaGateArea  0.2262 LAYER M6 ;
    AntennaGateArea  0.2262 LAYER M7 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
    AntennaDiffArea  0.8229 LAYER M2 ;
    AntennaDiffArea  0.8229 LAYER M3 ;
    AntennaDiffArea  0.8229 LAYER M4 ;
    AntennaDiffArea  0.8229 LAYER M5 ;
    AntennaDiffArea  0.8229 LAYER M6 ;
    AntennaDiffArea  0.8229 LAYER M7 ;
  END Z
END OR2HD2XSPGHT

MACRO OR2HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
END OR2HDLXHT

MACRO OR2HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1131 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END OR2HDMXHT

MACRO OR2HDUXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.0754 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0754 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3249 LAYER M1 ;
  END Z
END OR2HDUXHT

MACRO OR2ODHDHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1508 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1508 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6468 LAYER M1 ;
  END Z
END OR2ODHDHT

MACRO OR3HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END OR3HD1XHT

MACRO OR3HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2327 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OR3HD2XHT

MACRO OR3HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
END OR3HDLXHT

MACRO OR3HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END OR3HDMXHT

MACRO OR4HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END OR4HD1XHT

MACRO OR4HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2236 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2236 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2236 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.2236 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END OR4HD2XHT

MACRO OR4HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
END OR4HDLXHT

MACRO OR4HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END C
  PIN D
    #DIRECTION INPUT ;
    AntennaGateArea  0.1248 LAYER M1 ;
  END D
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END OR4HDMXHT

MACRO PULLDHDHT
  PIN EN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END EN
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.1095 LAYER M1 ;
  END Z
END PULLDHDHT

MACRO PULLUHDHT
  PIN E
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END E
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.1095 LAYER M1 ;
  END Z
END PULLUHDHT

MACRO RSLATHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.65545 LAYER M1 ;
  END Q
  PIN R
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END R
  PIN S
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END S
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.6213 LAYER M1 ;
  END QN
END RSLATHD1XHT

MACRO RSLATHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8844 LAYER M1 ;
  END Q
  PIN R
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END R
  PIN S
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END S
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.97665 LAYER M1 ;
  END QN
END RSLATHD2XHT

MACRO RSLATHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.252 LAYER M1 ;
  END Q
  PIN R
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END R
  PIN S
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END S
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2415 LAYER M1 ;
  END QN
END RSLATHDLXHT

MACRO RSLATHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.342 LAYER M1 ;
  END Q
  PIN R
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END R
  PIN S
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END S
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3315 LAYER M1 ;
  END QN
END RSLATHDMXHT

MACRO RSLATNHD1XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5875 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5845 LAYER M1 ;
  END QN
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END RSLATNHD1XHT

MACRO RSLATNHD2XHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8977 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END QN
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END RSLATNHD2XHT

MACRO RSLATNHDLXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2514 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END QN
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END RSLATNHDLXHT

MACRO RSLATNHDMXHT
  PIN Q
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3414 LAYER M1 ;
  END Q
  PIN QN
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.327 LAYER M1 ;
  END QN
  PIN RN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END RN
  PIN SN
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END SN
END RSLATNHDMXHT

MACRO TIEHHDHT
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.132 LAYER M1 ;
  END Z
END TIEHHDHT

MACRO TIELHDHT
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.1245 LAYER M1 ;
  END Z
END TIELHDHT

MACRO XNOR2HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2054 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1092 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.77015 LAYER M1 ;
  END Z
END XNOR2HD1XHT

MACRO XNOR2HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.3016 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END XNOR2HD2XHT

MACRO XNOR2HD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.3315 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END XNOR2HD3XHT

MACRO XNOR2HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2628 LAYER M1 ;
  END Z
END XNOR2HDLXHT

MACRO XNOR2HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3942 LAYER M1 ;
  END Z
END XNOR2HDMXHT

MACRO XNOR3HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1092 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.74905 LAYER M1 ;
  END Z
END XNOR3HD1XHT

MACRO XNOR3HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1755 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1027 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END XNOR3HD2XHT

MACRO XNOR3HD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1755 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1027 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END XNOR3HD3XHT

MACRO XNOR3HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2556 LAYER M1 ;
  END Z
END XNOR3HDLXHT

MACRO XNOR3HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3834 LAYER M1 ;
  END Z
END XNOR3HDMXHT

MACRO XOR2CLKHD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2145 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.5865 LAYER M1 ;
  END Z
END XOR2CLKHD1XHT

MACRO XOR2CLKHD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2145 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1365 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.68835 LAYER M1 ;
  END Z
END XOR2CLKHD2XHT

MACRO XOR2CLKHD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.2743 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.221 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.29383 LAYER M1 ;
  END Z
END XOR2CLKHD3XHT

MACRO XOR2CLKHD4XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.325 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2717 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.3884 LAYER M1 ;
  END Z
END XOR2CLKHD4XHT

MACRO XOR2HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1846 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1092 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.72795 LAYER M1 ;
  END Z
END XOR2HD1XHT

MACRO XOR2HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.26 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8229 LAYER M1 ;
  END Z
END XOR2HD2XHT

MACRO XOR2HD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.286 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END XOR2HD3XHT

MACRO XOR2HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
END XOR2HDLXHT

MACRO XOR2HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1716 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END XOR2HDMXHT

MACRO XOR3HD1XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1092 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.76485 LAYER M1 ;
  END Z
END XOR3HD1XHT

MACRO XOR3HD2XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.8862 LAYER M1 ;
  END Z
END XOR3HD2XHT

MACRO XOR3HD3XHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.2496 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  1.55085 LAYER M1 ;
  END Z
END XOR3HD3XHT

MACRO XOR3HDLXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.2484 LAYER M1 ;
  END Z
END XOR3HDLXHT

MACRO XOR3HDMXHT
  PIN A
    #DIRECTION INPUT ;
    AntennaGateArea  0.1872 LAYER M1 ;
  END A
  PIN B
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END B
  PIN C
    #DIRECTION INPUT ;
    AntennaGateArea  0.0936 LAYER M1 ;
  END C
  PIN Z
    #DIRECTION OUTPUT ;
    AntennaDiffArea  0.3726 LAYER M1 ;
  END Z
END XOR3HDMXHT

END LIBRARY
