
SITE  IOSite
    CLASS       PAD ;
    SYMMETRY    Y ;
    SIZE        0.005 BY 189.000 ;
END  IOSite

SITE  CornerSite
    CLASS	PAD ;
    SYMMETRY	R90 Y ;
    SIZE	189.000 BY 189.000 ;
END  CornerSite

MACRO PSESDCLAMP
  CLASS  PAD ;
  FOREIGN PSESDCLAMP 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 72.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 0.445 71.440 0.700 78.100 ;
        RECT 0.445 63.270 0.700 68.270 ;
        RECT 0.445 51.630 0.700 59.770 ;
        RECT 0.445 39.130 0.700 48.130 ;
        RECT 0.445 26.270 0.700 35.270 ;
        RECT 0.445 14.630 0.700 22.770 ;
        RECT 0.445 3.610 0.700 11.130 ;
        RECT 0.445 0.040 1.275 0.700 ;
        RECT 0.445 0.040 0.700 2.960 ;
        RECT 4.835 0.090 4.845 0.700 ;
        RECT 4.845 0.100 4.855 0.700 ;
        RECT 4.855 0.110 4.865 0.700 ;
        RECT 4.865 0.120 4.875 0.700 ;
        RECT 4.875 0.130 4.885 0.700 ;
        RECT 4.885 0.140 4.895 0.700 ;
        RECT 4.895 0.150 4.905 0.700 ;
        RECT 4.905 0.160 4.915 0.700 ;
        RECT 4.915 0.170 4.925 0.700 ;
        RECT 4.925 0.180 4.935 0.700 ;
        RECT 4.935 0.190 4.945 0.700 ;
        RECT 4.945 0.200 4.955 0.700 ;
        RECT 4.955 0.210 4.965 0.700 ;
        RECT 4.965 0.220 4.975 0.700 ;
        RECT 4.975 0.230 4.985 0.700 ;
        RECT 4.985 0.240 4.995 0.700 ;
        RECT 4.995 0.250 5.005 0.700 ;
        RECT 5.005 0.260 5.015 0.700 ;
        RECT 5.015 0.270 5.025 0.700 ;
        RECT 5.025 0.280 5.035 0.700 ;
        RECT 5.035 0.290 5.045 0.700 ;
        RECT 5.045 0.300 5.055 0.700 ;
        RECT 5.055 0.310 5.065 0.700 ;
        RECT 5.065 0.320 5.075 0.700 ;
        RECT 5.075 0.330 5.085 0.700 ;
        RECT 5.085 0.340 5.095 0.700 ;
        RECT 5.095 0.350 5.105 0.700 ;
        RECT 5.105 0.360 5.115 0.700 ;
        RECT 5.115 0.370 5.125 0.700 ;
        RECT 5.125 0.380 5.135 0.700 ;
        RECT 5.135 0.390 5.145 0.700 ;
        RECT 5.145 0.400 5.155 0.700 ;
        RECT 5.155 0.410 5.165 0.700 ;
        RECT 5.165 0.420 5.175 0.700 ;
        RECT 5.175 0.430 5.185 0.700 ;
        RECT 5.185 0.440 5.195 0.700 ;
        RECT 5.195 0.450 5.205 0.700 ;
        RECT 5.205 0.460 5.215 0.700 ;
        RECT 5.215 0.470 5.225 0.700 ;
        RECT 5.225 0.480 5.235 0.700 ;
        RECT 5.235 0.490 5.245 0.700 ;
        RECT 5.245 0.500 5.255 0.700 ;
        RECT 5.255 0.510 5.265 0.700 ;
        RECT 5.265 0.520 5.275 0.700 ;
        RECT 5.275 0.530 5.285 0.700 ;
        RECT 5.285 0.540 5.295 0.700 ;
        RECT 5.295 0.550 5.305 0.700 ;
        RECT 5.305 0.560 5.315 0.700 ;
        RECT 5.315 0.570 5.325 0.700 ;
        RECT 2.475 0.570 2.485 0.700 ;
        RECT 2.485 0.560 2.495 0.700 ;
        RECT 2.495 0.550 2.505 0.700 ;
        RECT 2.505 0.540 2.515 0.700 ;
        RECT 2.515 0.530 2.525 0.700 ;
        RECT 2.525 0.520 2.535 0.700 ;
        RECT 2.535 0.510 2.545 0.700 ;
        RECT 2.545 0.500 2.555 0.700 ;
        RECT 2.555 0.490 2.565 0.700 ;
        RECT 2.565 0.480 2.575 0.700 ;
        RECT 2.575 0.470 2.585 0.700 ;
        RECT 2.585 0.460 2.595 0.700 ;
        RECT 2.595 0.450 2.605 0.700 ;
        RECT 2.605 0.440 2.615 0.700 ;
        RECT 2.615 0.430 2.625 0.700 ;
        RECT 2.625 0.420 2.635 0.700 ;
        RECT 2.635 0.410 2.645 0.700 ;
        RECT 2.645 0.400 2.655 0.700 ;
        RECT 2.655 0.390 2.665 0.700 ;
        RECT 2.665 0.380 2.675 0.700 ;
        RECT 2.675 0.370 2.685 0.700 ;
        RECT 2.685 0.360 2.695 0.700 ;
        RECT 2.695 0.350 2.705 0.700 ;
        RECT 2.705 0.340 2.715 0.700 ;
        RECT 2.715 0.330 2.725 0.700 ;
        RECT 2.725 0.320 2.735 0.700 ;
        RECT 2.735 0.310 2.745 0.700 ;
        RECT 2.745 0.300 2.755 0.700 ;
        RECT 2.755 0.290 2.765 0.700 ;
        RECT 2.765 0.280 2.775 0.700 ;
        RECT 2.775 0.270 2.785 0.700 ;
        RECT 2.785 0.260 2.795 0.700 ;
        RECT 2.795 0.250 2.805 0.700 ;
        RECT 2.805 0.240 2.815 0.700 ;
        RECT 2.815 0.230 2.825 0.700 ;
        RECT 2.825 0.220 2.835 0.700 ;
        RECT 2.835 0.210 2.845 0.700 ;
        RECT 2.845 0.200 2.855 0.700 ;
        RECT 2.855 0.190 2.865 0.700 ;
        RECT 2.865 0.180 2.875 0.700 ;
        RECT 2.875 0.170 2.885 0.700 ;
        RECT 2.885 0.160 2.895 0.700 ;
        RECT 2.895 0.150 2.905 0.700 ;
        RECT 2.905 0.140 2.915 0.700 ;
        RECT 2.915 0.130 2.925 0.700 ;
        RECT 2.925 0.120 2.935 0.700 ;
        RECT 2.935 0.110 2.945 0.700 ;
        RECT 2.945 0.100 2.955 0.700 ;
        RECT 2.955 0.090 2.965 0.700 ;
        RECT 2.965 0.080 4.835 0.700 ;
        RECT 11.255 0.090 11.265 0.700 ;
        RECT 11.265 0.100 11.275 0.700 ;
        RECT 11.275 0.110 11.285 0.700 ;
        RECT 11.285 0.120 11.295 0.700 ;
        RECT 11.295 0.130 11.305 0.700 ;
        RECT 11.305 0.140 11.315 0.700 ;
        RECT 11.315 0.150 11.325 0.700 ;
        RECT 11.325 0.160 11.335 0.700 ;
        RECT 11.335 0.170 11.345 0.700 ;
        RECT 11.345 0.180 11.355 0.700 ;
        RECT 11.355 0.190 11.365 0.700 ;
        RECT 11.365 0.200 11.375 0.700 ;
        RECT 11.375 0.210 11.385 0.700 ;
        RECT 11.385 0.220 11.395 0.700 ;
        RECT 11.395 0.230 11.405 0.700 ;
        RECT 11.405 0.240 11.415 0.700 ;
        RECT 11.415 0.250 11.425 0.700 ;
        RECT 11.425 0.260 11.435 0.700 ;
        RECT 11.435 0.270 11.445 0.700 ;
        RECT 11.445 0.280 11.455 0.700 ;
        RECT 11.455 0.290 11.465 0.700 ;
        RECT 11.465 0.300 11.475 0.700 ;
        RECT 11.475 0.310 11.485 0.700 ;
        RECT 11.485 0.320 11.495 0.700 ;
        RECT 11.495 0.330 11.505 0.700 ;
        RECT 11.505 0.340 11.515 0.700 ;
        RECT 11.515 0.350 11.525 0.700 ;
        RECT 11.525 0.360 11.535 0.700 ;
        RECT 11.535 0.370 11.545 0.700 ;
        RECT 11.545 0.380 11.555 0.700 ;
        RECT 11.555 0.390 11.565 0.700 ;
        RECT 11.565 0.400 11.575 0.700 ;
        RECT 11.575 0.410 11.585 0.700 ;
        RECT 11.585 0.420 11.595 0.700 ;
        RECT 11.595 0.430 11.605 0.700 ;
        RECT 11.605 0.440 11.615 0.700 ;
        RECT 11.615 0.450 11.625 0.700 ;
        RECT 11.625 0.460 11.635 0.700 ;
        RECT 11.635 0.470 11.645 0.700 ;
        RECT 11.645 0.480 11.655 0.700 ;
        RECT 11.655 0.490 11.665 0.700 ;
        RECT 11.665 0.500 11.675 0.700 ;
        RECT 11.675 0.510 11.685 0.700 ;
        RECT 11.685 0.520 11.695 0.700 ;
        RECT 11.695 0.530 11.705 0.700 ;
        RECT 11.705 0.540 11.715 0.700 ;
        RECT 11.715 0.550 11.725 0.700 ;
        RECT 11.725 0.560 11.735 0.700 ;
        RECT 11.735 0.570 11.745 0.700 ;
        RECT 8.895 0.570 8.905 0.700 ;
        RECT 8.905 0.560 8.915 0.700 ;
        RECT 8.915 0.550 8.925 0.700 ;
        RECT 8.925 0.540 8.935 0.700 ;
        RECT 8.935 0.530 8.945 0.700 ;
        RECT 8.945 0.520 8.955 0.700 ;
        RECT 8.955 0.510 8.965 0.700 ;
        RECT 8.965 0.500 8.975 0.700 ;
        RECT 8.975 0.490 8.985 0.700 ;
        RECT 8.985 0.480 8.995 0.700 ;
        RECT 8.995 0.470 9.005 0.700 ;
        RECT 9.005 0.460 9.015 0.700 ;
        RECT 9.015 0.450 9.025 0.700 ;
        RECT 9.025 0.440 9.035 0.700 ;
        RECT 9.035 0.430 9.045 0.700 ;
        RECT 9.045 0.420 9.055 0.700 ;
        RECT 9.055 0.410 9.065 0.700 ;
        RECT 9.065 0.400 9.075 0.700 ;
        RECT 9.075 0.390 9.085 0.700 ;
        RECT 9.085 0.380 9.095 0.700 ;
        RECT 9.095 0.370 9.105 0.700 ;
        RECT 9.105 0.360 9.115 0.700 ;
        RECT 9.115 0.350 9.125 0.700 ;
        RECT 9.125 0.340 9.135 0.700 ;
        RECT 9.135 0.330 9.145 0.700 ;
        RECT 9.145 0.320 9.155 0.700 ;
        RECT 9.155 0.310 9.165 0.700 ;
        RECT 9.165 0.300 9.175 0.700 ;
        RECT 9.175 0.290 9.185 0.700 ;
        RECT 9.185 0.280 9.195 0.700 ;
        RECT 9.195 0.270 9.205 0.700 ;
        RECT 9.205 0.260 9.215 0.700 ;
        RECT 9.215 0.250 9.225 0.700 ;
        RECT 9.225 0.240 9.235 0.700 ;
        RECT 9.235 0.230 9.245 0.700 ;
        RECT 9.245 0.220 9.255 0.700 ;
        RECT 9.255 0.210 9.265 0.700 ;
        RECT 9.265 0.200 9.275 0.700 ;
        RECT 9.275 0.190 9.285 0.700 ;
        RECT 9.285 0.180 9.295 0.700 ;
        RECT 9.295 0.170 9.305 0.700 ;
        RECT 9.305 0.160 9.315 0.700 ;
        RECT 9.315 0.150 9.325 0.700 ;
        RECT 9.325 0.140 9.335 0.700 ;
        RECT 9.335 0.130 9.345 0.700 ;
        RECT 9.345 0.120 9.355 0.700 ;
        RECT 9.355 0.110 9.365 0.700 ;
        RECT 9.365 0.100 9.375 0.700 ;
        RECT 9.375 0.090 9.385 0.700 ;
        RECT 9.385 0.080 11.255 0.700 ;
        RECT 17.675 0.090 17.685 0.700 ;
        RECT 17.685 0.100 17.695 0.700 ;
        RECT 17.695 0.110 17.705 0.700 ;
        RECT 17.705 0.120 17.715 0.700 ;
        RECT 17.715 0.130 17.725 0.700 ;
        RECT 17.725 0.140 17.735 0.700 ;
        RECT 17.735 0.150 17.745 0.700 ;
        RECT 17.745 0.160 17.755 0.700 ;
        RECT 17.755 0.170 17.765 0.700 ;
        RECT 17.765 0.180 17.775 0.700 ;
        RECT 17.775 0.190 17.785 0.700 ;
        RECT 17.785 0.200 17.795 0.700 ;
        RECT 17.795 0.210 17.805 0.700 ;
        RECT 17.805 0.220 17.815 0.700 ;
        RECT 17.815 0.230 17.825 0.700 ;
        RECT 17.825 0.240 17.835 0.700 ;
        RECT 17.835 0.250 17.845 0.700 ;
        RECT 17.845 0.260 17.855 0.700 ;
        RECT 17.855 0.270 17.865 0.700 ;
        RECT 17.865 0.280 17.875 0.700 ;
        RECT 17.875 0.290 17.885 0.700 ;
        RECT 17.885 0.300 17.895 0.700 ;
        RECT 17.895 0.310 17.905 0.700 ;
        RECT 17.905 0.320 17.915 0.700 ;
        RECT 17.915 0.330 17.925 0.700 ;
        RECT 17.925 0.340 17.935 0.700 ;
        RECT 17.935 0.350 17.945 0.700 ;
        RECT 17.945 0.360 17.955 0.700 ;
        RECT 17.955 0.370 17.965 0.700 ;
        RECT 17.965 0.380 17.975 0.700 ;
        RECT 17.975 0.390 17.985 0.700 ;
        RECT 17.985 0.400 17.995 0.700 ;
        RECT 17.995 0.410 18.005 0.700 ;
        RECT 18.005 0.420 18.015 0.700 ;
        RECT 18.015 0.430 18.025 0.700 ;
        RECT 18.025 0.440 18.035 0.700 ;
        RECT 18.035 0.450 18.045 0.700 ;
        RECT 18.045 0.460 18.055 0.700 ;
        RECT 18.055 0.470 18.065 0.700 ;
        RECT 18.065 0.480 18.075 0.700 ;
        RECT 18.075 0.490 18.085 0.700 ;
        RECT 18.085 0.500 18.095 0.700 ;
        RECT 18.095 0.510 18.105 0.700 ;
        RECT 18.105 0.520 18.115 0.700 ;
        RECT 18.115 0.530 18.125 0.700 ;
        RECT 18.125 0.540 18.135 0.700 ;
        RECT 18.135 0.550 18.145 0.700 ;
        RECT 18.145 0.560 18.155 0.700 ;
        RECT 18.155 0.570 18.165 0.700 ;
        RECT 15.315 0.570 15.325 0.700 ;
        RECT 15.325 0.560 15.335 0.700 ;
        RECT 15.335 0.550 15.345 0.700 ;
        RECT 15.345 0.540 15.355 0.700 ;
        RECT 15.355 0.530 15.365 0.700 ;
        RECT 15.365 0.520 15.375 0.700 ;
        RECT 15.375 0.510 15.385 0.700 ;
        RECT 15.385 0.500 15.395 0.700 ;
        RECT 15.395 0.490 15.405 0.700 ;
        RECT 15.405 0.480 15.415 0.700 ;
        RECT 15.415 0.470 15.425 0.700 ;
        RECT 15.425 0.460 15.435 0.700 ;
        RECT 15.435 0.450 15.445 0.700 ;
        RECT 15.445 0.440 15.455 0.700 ;
        RECT 15.455 0.430 15.465 0.700 ;
        RECT 15.465 0.420 15.475 0.700 ;
        RECT 15.475 0.410 15.485 0.700 ;
        RECT 15.485 0.400 15.495 0.700 ;
        RECT 15.495 0.390 15.505 0.700 ;
        RECT 15.505 0.380 15.515 0.700 ;
        RECT 15.515 0.370 15.525 0.700 ;
        RECT 15.525 0.360 15.535 0.700 ;
        RECT 15.535 0.350 15.545 0.700 ;
        RECT 15.545 0.340 15.555 0.700 ;
        RECT 15.555 0.330 15.565 0.700 ;
        RECT 15.565 0.320 15.575 0.700 ;
        RECT 15.575 0.310 15.585 0.700 ;
        RECT 15.585 0.300 15.595 0.700 ;
        RECT 15.595 0.290 15.605 0.700 ;
        RECT 15.605 0.280 15.615 0.700 ;
        RECT 15.615 0.270 15.625 0.700 ;
        RECT 15.625 0.260 15.635 0.700 ;
        RECT 15.635 0.250 15.645 0.700 ;
        RECT 15.645 0.240 15.655 0.700 ;
        RECT 15.655 0.230 15.665 0.700 ;
        RECT 15.665 0.220 15.675 0.700 ;
        RECT 15.675 0.210 15.685 0.700 ;
        RECT 15.685 0.200 15.695 0.700 ;
        RECT 15.695 0.190 15.705 0.700 ;
        RECT 15.705 0.180 15.715 0.700 ;
        RECT 15.715 0.170 15.725 0.700 ;
        RECT 15.725 0.160 15.735 0.700 ;
        RECT 15.735 0.150 15.745 0.700 ;
        RECT 15.745 0.140 15.755 0.700 ;
        RECT 15.755 0.130 15.765 0.700 ;
        RECT 15.765 0.120 15.775 0.700 ;
        RECT 15.775 0.110 15.785 0.700 ;
        RECT 15.785 0.100 15.795 0.700 ;
        RECT 15.795 0.090 15.805 0.700 ;
        RECT 15.805 0.080 17.675 0.700 ;
        RECT 24.095 0.090 24.105 0.700 ;
        RECT 24.105 0.100 24.115 0.700 ;
        RECT 24.115 0.110 24.125 0.700 ;
        RECT 24.125 0.120 24.135 0.700 ;
        RECT 24.135 0.130 24.145 0.700 ;
        RECT 24.145 0.140 24.155 0.700 ;
        RECT 24.155 0.150 24.165 0.700 ;
        RECT 24.165 0.160 24.175 0.700 ;
        RECT 24.175 0.170 24.185 0.700 ;
        RECT 24.185 0.180 24.195 0.700 ;
        RECT 24.195 0.190 24.205 0.700 ;
        RECT 24.205 0.200 24.215 0.700 ;
        RECT 24.215 0.210 24.225 0.700 ;
        RECT 24.225 0.220 24.235 0.700 ;
        RECT 24.235 0.230 24.245 0.700 ;
        RECT 24.245 0.240 24.255 0.700 ;
        RECT 24.255 0.250 24.265 0.700 ;
        RECT 24.265 0.260 24.275 0.700 ;
        RECT 24.275 0.270 24.285 0.700 ;
        RECT 24.285 0.280 24.295 0.700 ;
        RECT 24.295 0.290 24.305 0.700 ;
        RECT 24.305 0.300 24.315 0.700 ;
        RECT 24.315 0.310 24.325 0.700 ;
        RECT 24.325 0.320 24.335 0.700 ;
        RECT 24.335 0.330 24.345 0.700 ;
        RECT 24.345 0.340 24.355 0.700 ;
        RECT 24.355 0.350 24.365 0.700 ;
        RECT 24.365 0.360 24.375 0.700 ;
        RECT 24.375 0.370 24.385 0.700 ;
        RECT 24.385 0.380 24.395 0.700 ;
        RECT 24.395 0.390 24.405 0.700 ;
        RECT 24.405 0.400 24.415 0.700 ;
        RECT 24.415 0.410 24.425 0.700 ;
        RECT 24.425 0.420 24.435 0.700 ;
        RECT 24.435 0.430 24.445 0.700 ;
        RECT 24.445 0.440 24.455 0.700 ;
        RECT 24.455 0.450 24.465 0.700 ;
        RECT 24.465 0.460 24.475 0.700 ;
        RECT 24.475 0.470 24.485 0.700 ;
        RECT 24.485 0.480 24.495 0.700 ;
        RECT 24.495 0.490 24.505 0.700 ;
        RECT 24.505 0.500 24.515 0.700 ;
        RECT 24.515 0.510 24.525 0.700 ;
        RECT 24.525 0.520 24.535 0.700 ;
        RECT 24.535 0.530 24.545 0.700 ;
        RECT 24.545 0.540 24.555 0.700 ;
        RECT 24.555 0.550 24.565 0.700 ;
        RECT 24.565 0.560 24.575 0.700 ;
        RECT 24.575 0.570 24.585 0.700 ;
        RECT 21.735 0.570 21.745 0.700 ;
        RECT 21.745 0.560 21.755 0.700 ;
        RECT 21.755 0.550 21.765 0.700 ;
        RECT 21.765 0.540 21.775 0.700 ;
        RECT 21.775 0.530 21.785 0.700 ;
        RECT 21.785 0.520 21.795 0.700 ;
        RECT 21.795 0.510 21.805 0.700 ;
        RECT 21.805 0.500 21.815 0.700 ;
        RECT 21.815 0.490 21.825 0.700 ;
        RECT 21.825 0.480 21.835 0.700 ;
        RECT 21.835 0.470 21.845 0.700 ;
        RECT 21.845 0.460 21.855 0.700 ;
        RECT 21.855 0.450 21.865 0.700 ;
        RECT 21.865 0.440 21.875 0.700 ;
        RECT 21.875 0.430 21.885 0.700 ;
        RECT 21.885 0.420 21.895 0.700 ;
        RECT 21.895 0.410 21.905 0.700 ;
        RECT 21.905 0.400 21.915 0.700 ;
        RECT 21.915 0.390 21.925 0.700 ;
        RECT 21.925 0.380 21.935 0.700 ;
        RECT 21.935 0.370 21.945 0.700 ;
        RECT 21.945 0.360 21.955 0.700 ;
        RECT 21.955 0.350 21.965 0.700 ;
        RECT 21.965 0.340 21.975 0.700 ;
        RECT 21.975 0.330 21.985 0.700 ;
        RECT 21.985 0.320 21.995 0.700 ;
        RECT 21.995 0.310 22.005 0.700 ;
        RECT 22.005 0.300 22.015 0.700 ;
        RECT 22.015 0.290 22.025 0.700 ;
        RECT 22.025 0.280 22.035 0.700 ;
        RECT 22.035 0.270 22.045 0.700 ;
        RECT 22.045 0.260 22.055 0.700 ;
        RECT 22.055 0.250 22.065 0.700 ;
        RECT 22.065 0.240 22.075 0.700 ;
        RECT 22.075 0.230 22.085 0.700 ;
        RECT 22.085 0.220 22.095 0.700 ;
        RECT 22.095 0.210 22.105 0.700 ;
        RECT 22.105 0.200 22.115 0.700 ;
        RECT 22.115 0.190 22.125 0.700 ;
        RECT 22.125 0.180 22.135 0.700 ;
        RECT 22.135 0.170 22.145 0.700 ;
        RECT 22.145 0.160 22.155 0.700 ;
        RECT 22.155 0.150 22.165 0.700 ;
        RECT 22.165 0.140 22.175 0.700 ;
        RECT 22.175 0.130 22.185 0.700 ;
        RECT 22.185 0.120 22.195 0.700 ;
        RECT 22.195 0.110 22.205 0.700 ;
        RECT 22.205 0.100 22.215 0.700 ;
        RECT 22.215 0.090 22.225 0.700 ;
        RECT 22.225 0.080 24.095 0.700 ;
        RECT 30.515 0.090 30.525 0.700 ;
        RECT 30.525 0.100 30.535 0.700 ;
        RECT 30.535 0.110 30.545 0.700 ;
        RECT 30.545 0.120 30.555 0.700 ;
        RECT 30.555 0.130 30.565 0.700 ;
        RECT 30.565 0.140 30.575 0.700 ;
        RECT 30.575 0.150 30.585 0.700 ;
        RECT 30.585 0.160 30.595 0.700 ;
        RECT 30.595 0.170 30.605 0.700 ;
        RECT 30.605 0.180 30.615 0.700 ;
        RECT 30.615 0.190 30.625 0.700 ;
        RECT 30.625 0.200 30.635 0.700 ;
        RECT 30.635 0.210 30.645 0.700 ;
        RECT 30.645 0.220 30.655 0.700 ;
        RECT 30.655 0.230 30.665 0.700 ;
        RECT 30.665 0.240 30.675 0.700 ;
        RECT 30.675 0.250 30.685 0.700 ;
        RECT 30.685 0.260 30.695 0.700 ;
        RECT 30.695 0.270 30.705 0.700 ;
        RECT 30.705 0.280 30.715 0.700 ;
        RECT 30.715 0.290 30.725 0.700 ;
        RECT 30.725 0.300 30.735 0.700 ;
        RECT 30.735 0.310 30.745 0.700 ;
        RECT 30.745 0.320 30.755 0.700 ;
        RECT 30.755 0.330 30.765 0.700 ;
        RECT 30.765 0.340 30.775 0.700 ;
        RECT 30.775 0.350 30.785 0.700 ;
        RECT 30.785 0.360 30.795 0.700 ;
        RECT 30.795 0.370 30.805 0.700 ;
        RECT 30.805 0.380 30.815 0.700 ;
        RECT 30.815 0.390 30.825 0.700 ;
        RECT 30.825 0.400 30.835 0.700 ;
        RECT 30.835 0.410 30.845 0.700 ;
        RECT 30.845 0.420 30.855 0.700 ;
        RECT 30.855 0.430 30.865 0.700 ;
        RECT 30.865 0.440 30.875 0.700 ;
        RECT 30.875 0.450 30.885 0.700 ;
        RECT 30.885 0.460 30.895 0.700 ;
        RECT 30.895 0.470 30.905 0.700 ;
        RECT 30.905 0.480 30.915 0.700 ;
        RECT 30.915 0.490 30.925 0.700 ;
        RECT 30.925 0.500 30.935 0.700 ;
        RECT 30.935 0.510 30.945 0.700 ;
        RECT 30.945 0.520 30.955 0.700 ;
        RECT 30.955 0.530 30.965 0.700 ;
        RECT 30.965 0.540 30.975 0.700 ;
        RECT 30.975 0.550 30.985 0.700 ;
        RECT 30.985 0.560 30.995 0.700 ;
        RECT 30.995 0.570 31.005 0.700 ;
        RECT 28.155 0.570 28.165 0.700 ;
        RECT 28.165 0.560 28.175 0.700 ;
        RECT 28.175 0.550 28.185 0.700 ;
        RECT 28.185 0.540 28.195 0.700 ;
        RECT 28.195 0.530 28.205 0.700 ;
        RECT 28.205 0.520 28.215 0.700 ;
        RECT 28.215 0.510 28.225 0.700 ;
        RECT 28.225 0.500 28.235 0.700 ;
        RECT 28.235 0.490 28.245 0.700 ;
        RECT 28.245 0.480 28.255 0.700 ;
        RECT 28.255 0.470 28.265 0.700 ;
        RECT 28.265 0.460 28.275 0.700 ;
        RECT 28.275 0.450 28.285 0.700 ;
        RECT 28.285 0.440 28.295 0.700 ;
        RECT 28.295 0.430 28.305 0.700 ;
        RECT 28.305 0.420 28.315 0.700 ;
        RECT 28.315 0.410 28.325 0.700 ;
        RECT 28.325 0.400 28.335 0.700 ;
        RECT 28.335 0.390 28.345 0.700 ;
        RECT 28.345 0.380 28.355 0.700 ;
        RECT 28.355 0.370 28.365 0.700 ;
        RECT 28.365 0.360 28.375 0.700 ;
        RECT 28.375 0.350 28.385 0.700 ;
        RECT 28.385 0.340 28.395 0.700 ;
        RECT 28.395 0.330 28.405 0.700 ;
        RECT 28.405 0.320 28.415 0.700 ;
        RECT 28.415 0.310 28.425 0.700 ;
        RECT 28.425 0.300 28.435 0.700 ;
        RECT 28.435 0.290 28.445 0.700 ;
        RECT 28.445 0.280 28.455 0.700 ;
        RECT 28.455 0.270 28.465 0.700 ;
        RECT 28.465 0.260 28.475 0.700 ;
        RECT 28.475 0.250 28.485 0.700 ;
        RECT 28.485 0.240 28.495 0.700 ;
        RECT 28.495 0.230 28.505 0.700 ;
        RECT 28.505 0.220 28.515 0.700 ;
        RECT 28.515 0.210 28.525 0.700 ;
        RECT 28.525 0.200 28.535 0.700 ;
        RECT 28.535 0.190 28.545 0.700 ;
        RECT 28.545 0.180 28.555 0.700 ;
        RECT 28.555 0.170 28.565 0.700 ;
        RECT 28.565 0.160 28.575 0.700 ;
        RECT 28.575 0.150 28.585 0.700 ;
        RECT 28.585 0.140 28.595 0.700 ;
        RECT 28.595 0.130 28.605 0.700 ;
        RECT 28.605 0.120 28.615 0.700 ;
        RECT 28.615 0.110 28.625 0.700 ;
        RECT 28.625 0.100 28.635 0.700 ;
        RECT 28.635 0.090 28.645 0.700 ;
        RECT 28.645 0.080 30.515 0.700 ;
        RECT 36.935 0.090 36.945 0.700 ;
        RECT 36.945 0.100 36.955 0.700 ;
        RECT 36.955 0.110 36.965 0.700 ;
        RECT 36.965 0.120 36.975 0.700 ;
        RECT 36.975 0.130 36.985 0.700 ;
        RECT 36.985 0.140 36.995 0.700 ;
        RECT 36.995 0.150 37.005 0.700 ;
        RECT 37.005 0.160 37.015 0.700 ;
        RECT 37.015 0.170 37.025 0.700 ;
        RECT 37.025 0.180 37.035 0.700 ;
        RECT 37.035 0.190 37.045 0.700 ;
        RECT 37.045 0.200 37.055 0.700 ;
        RECT 37.055 0.210 37.065 0.700 ;
        RECT 37.065 0.220 37.075 0.700 ;
        RECT 37.075 0.230 37.085 0.700 ;
        RECT 37.085 0.240 37.095 0.700 ;
        RECT 37.095 0.250 37.105 0.700 ;
        RECT 37.105 0.260 37.115 0.700 ;
        RECT 37.115 0.270 37.125 0.700 ;
        RECT 37.125 0.280 37.135 0.700 ;
        RECT 37.135 0.290 37.145 0.700 ;
        RECT 37.145 0.300 37.155 0.700 ;
        RECT 37.155 0.310 37.165 0.700 ;
        RECT 37.165 0.320 37.175 0.700 ;
        RECT 37.175 0.330 37.185 0.700 ;
        RECT 37.185 0.340 37.195 0.700 ;
        RECT 37.195 0.350 37.205 0.700 ;
        RECT 37.205 0.360 37.215 0.700 ;
        RECT 37.215 0.370 37.225 0.700 ;
        RECT 37.225 0.380 37.235 0.700 ;
        RECT 37.235 0.390 37.245 0.700 ;
        RECT 37.245 0.400 37.255 0.700 ;
        RECT 37.255 0.410 37.265 0.700 ;
        RECT 37.265 0.420 37.275 0.700 ;
        RECT 37.275 0.430 37.285 0.700 ;
        RECT 37.285 0.440 37.295 0.700 ;
        RECT 37.295 0.450 37.305 0.700 ;
        RECT 37.305 0.460 37.315 0.700 ;
        RECT 37.315 0.470 37.325 0.700 ;
        RECT 37.325 0.480 37.335 0.700 ;
        RECT 37.335 0.490 37.345 0.700 ;
        RECT 37.345 0.500 37.355 0.700 ;
        RECT 37.355 0.510 37.365 0.700 ;
        RECT 37.365 0.520 37.375 0.700 ;
        RECT 37.375 0.530 37.385 0.700 ;
        RECT 37.385 0.540 37.395 0.700 ;
        RECT 37.395 0.550 37.405 0.700 ;
        RECT 37.405 0.560 37.415 0.700 ;
        RECT 37.415 0.570 37.425 0.700 ;
        RECT 34.575 0.570 34.585 0.700 ;
        RECT 34.585 0.560 34.595 0.700 ;
        RECT 34.595 0.550 34.605 0.700 ;
        RECT 34.605 0.540 34.615 0.700 ;
        RECT 34.615 0.530 34.625 0.700 ;
        RECT 34.625 0.520 34.635 0.700 ;
        RECT 34.635 0.510 34.645 0.700 ;
        RECT 34.645 0.500 34.655 0.700 ;
        RECT 34.655 0.490 34.665 0.700 ;
        RECT 34.665 0.480 34.675 0.700 ;
        RECT 34.675 0.470 34.685 0.700 ;
        RECT 34.685 0.460 34.695 0.700 ;
        RECT 34.695 0.450 34.705 0.700 ;
        RECT 34.705 0.440 34.715 0.700 ;
        RECT 34.715 0.430 34.725 0.700 ;
        RECT 34.725 0.420 34.735 0.700 ;
        RECT 34.735 0.410 34.745 0.700 ;
        RECT 34.745 0.400 34.755 0.700 ;
        RECT 34.755 0.390 34.765 0.700 ;
        RECT 34.765 0.380 34.775 0.700 ;
        RECT 34.775 0.370 34.785 0.700 ;
        RECT 34.785 0.360 34.795 0.700 ;
        RECT 34.795 0.350 34.805 0.700 ;
        RECT 34.805 0.340 34.815 0.700 ;
        RECT 34.815 0.330 34.825 0.700 ;
        RECT 34.825 0.320 34.835 0.700 ;
        RECT 34.835 0.310 34.845 0.700 ;
        RECT 34.845 0.300 34.855 0.700 ;
        RECT 34.855 0.290 34.865 0.700 ;
        RECT 34.865 0.280 34.875 0.700 ;
        RECT 34.875 0.270 34.885 0.700 ;
        RECT 34.885 0.260 34.895 0.700 ;
        RECT 34.895 0.250 34.905 0.700 ;
        RECT 34.905 0.240 34.915 0.700 ;
        RECT 34.915 0.230 34.925 0.700 ;
        RECT 34.925 0.220 34.935 0.700 ;
        RECT 34.935 0.210 34.945 0.700 ;
        RECT 34.945 0.200 34.955 0.700 ;
        RECT 34.955 0.190 34.965 0.700 ;
        RECT 34.965 0.180 34.975 0.700 ;
        RECT 34.975 0.170 34.985 0.700 ;
        RECT 34.985 0.160 34.995 0.700 ;
        RECT 34.995 0.150 35.005 0.700 ;
        RECT 35.005 0.140 35.015 0.700 ;
        RECT 35.015 0.130 35.025 0.700 ;
        RECT 35.025 0.120 35.035 0.700 ;
        RECT 35.035 0.110 35.045 0.700 ;
        RECT 35.045 0.100 35.055 0.700 ;
        RECT 35.055 0.090 35.065 0.700 ;
        RECT 35.065 0.080 36.935 0.700 ;
        RECT 43.355 0.090 43.365 0.700 ;
        RECT 43.365 0.100 43.375 0.700 ;
        RECT 43.375 0.110 43.385 0.700 ;
        RECT 43.385 0.120 43.395 0.700 ;
        RECT 43.395 0.130 43.405 0.700 ;
        RECT 43.405 0.140 43.415 0.700 ;
        RECT 43.415 0.150 43.425 0.700 ;
        RECT 43.425 0.160 43.435 0.700 ;
        RECT 43.435 0.170 43.445 0.700 ;
        RECT 43.445 0.180 43.455 0.700 ;
        RECT 43.455 0.190 43.465 0.700 ;
        RECT 43.465 0.200 43.475 0.700 ;
        RECT 43.475 0.210 43.485 0.700 ;
        RECT 43.485 0.220 43.495 0.700 ;
        RECT 43.495 0.230 43.505 0.700 ;
        RECT 43.505 0.240 43.515 0.700 ;
        RECT 43.515 0.250 43.525 0.700 ;
        RECT 43.525 0.260 43.535 0.700 ;
        RECT 43.535 0.270 43.545 0.700 ;
        RECT 43.545 0.280 43.555 0.700 ;
        RECT 43.555 0.290 43.565 0.700 ;
        RECT 43.565 0.300 43.575 0.700 ;
        RECT 43.575 0.310 43.585 0.700 ;
        RECT 43.585 0.320 43.595 0.700 ;
        RECT 43.595 0.330 43.605 0.700 ;
        RECT 43.605 0.340 43.615 0.700 ;
        RECT 43.615 0.350 43.625 0.700 ;
        RECT 43.625 0.360 43.635 0.700 ;
        RECT 43.635 0.370 43.645 0.700 ;
        RECT 43.645 0.380 43.655 0.700 ;
        RECT 43.655 0.390 43.665 0.700 ;
        RECT 43.665 0.400 43.675 0.700 ;
        RECT 43.675 0.410 43.685 0.700 ;
        RECT 43.685 0.420 43.695 0.700 ;
        RECT 43.695 0.430 43.705 0.700 ;
        RECT 43.705 0.440 43.715 0.700 ;
        RECT 43.715 0.450 43.725 0.700 ;
        RECT 43.725 0.460 43.735 0.700 ;
        RECT 43.735 0.470 43.745 0.700 ;
        RECT 43.745 0.480 43.755 0.700 ;
        RECT 43.755 0.490 43.765 0.700 ;
        RECT 43.765 0.500 43.775 0.700 ;
        RECT 43.775 0.510 43.785 0.700 ;
        RECT 43.785 0.520 43.795 0.700 ;
        RECT 43.795 0.530 43.805 0.700 ;
        RECT 43.805 0.540 43.815 0.700 ;
        RECT 43.815 0.550 43.825 0.700 ;
        RECT 43.825 0.560 43.835 0.700 ;
        RECT 43.835 0.570 43.845 0.700 ;
        RECT 40.995 0.570 41.005 0.700 ;
        RECT 41.005 0.560 41.015 0.700 ;
        RECT 41.015 0.550 41.025 0.700 ;
        RECT 41.025 0.540 41.035 0.700 ;
        RECT 41.035 0.530 41.045 0.700 ;
        RECT 41.045 0.520 41.055 0.700 ;
        RECT 41.055 0.510 41.065 0.700 ;
        RECT 41.065 0.500 41.075 0.700 ;
        RECT 41.075 0.490 41.085 0.700 ;
        RECT 41.085 0.480 41.095 0.700 ;
        RECT 41.095 0.470 41.105 0.700 ;
        RECT 41.105 0.460 41.115 0.700 ;
        RECT 41.115 0.450 41.125 0.700 ;
        RECT 41.125 0.440 41.135 0.700 ;
        RECT 41.135 0.430 41.145 0.700 ;
        RECT 41.145 0.420 41.155 0.700 ;
        RECT 41.155 0.410 41.165 0.700 ;
        RECT 41.165 0.400 41.175 0.700 ;
        RECT 41.175 0.390 41.185 0.700 ;
        RECT 41.185 0.380 41.195 0.700 ;
        RECT 41.195 0.370 41.205 0.700 ;
        RECT 41.205 0.360 41.215 0.700 ;
        RECT 41.215 0.350 41.225 0.700 ;
        RECT 41.225 0.340 41.235 0.700 ;
        RECT 41.235 0.330 41.245 0.700 ;
        RECT 41.245 0.320 41.255 0.700 ;
        RECT 41.255 0.310 41.265 0.700 ;
        RECT 41.265 0.300 41.275 0.700 ;
        RECT 41.275 0.290 41.285 0.700 ;
        RECT 41.285 0.280 41.295 0.700 ;
        RECT 41.295 0.270 41.305 0.700 ;
        RECT 41.305 0.260 41.315 0.700 ;
        RECT 41.315 0.250 41.325 0.700 ;
        RECT 41.325 0.240 41.335 0.700 ;
        RECT 41.335 0.230 41.345 0.700 ;
        RECT 41.345 0.220 41.355 0.700 ;
        RECT 41.355 0.210 41.365 0.700 ;
        RECT 41.365 0.200 41.375 0.700 ;
        RECT 41.375 0.190 41.385 0.700 ;
        RECT 41.385 0.180 41.395 0.700 ;
        RECT 41.395 0.170 41.405 0.700 ;
        RECT 41.405 0.160 41.415 0.700 ;
        RECT 41.415 0.150 41.425 0.700 ;
        RECT 41.425 0.140 41.435 0.700 ;
        RECT 41.435 0.130 41.445 0.700 ;
        RECT 41.445 0.120 41.455 0.700 ;
        RECT 41.455 0.110 41.465 0.700 ;
        RECT 41.465 0.100 41.475 0.700 ;
        RECT 41.475 0.090 41.485 0.700 ;
        RECT 41.485 0.080 43.355 0.700 ;
        RECT 49.775 0.090 49.785 0.700 ;
        RECT 49.785 0.100 49.795 0.700 ;
        RECT 49.795 0.110 49.805 0.700 ;
        RECT 49.805 0.120 49.815 0.700 ;
        RECT 49.815 0.130 49.825 0.700 ;
        RECT 49.825 0.140 49.835 0.700 ;
        RECT 49.835 0.150 49.845 0.700 ;
        RECT 49.845 0.160 49.855 0.700 ;
        RECT 49.855 0.170 49.865 0.700 ;
        RECT 49.865 0.180 49.875 0.700 ;
        RECT 49.875 0.190 49.885 0.700 ;
        RECT 49.885 0.200 49.895 0.700 ;
        RECT 49.895 0.210 49.905 0.700 ;
        RECT 49.905 0.220 49.915 0.700 ;
        RECT 49.915 0.230 49.925 0.700 ;
        RECT 49.925 0.240 49.935 0.700 ;
        RECT 49.935 0.250 49.945 0.700 ;
        RECT 49.945 0.260 49.955 0.700 ;
        RECT 49.955 0.270 49.965 0.700 ;
        RECT 49.965 0.280 49.975 0.700 ;
        RECT 49.975 0.290 49.985 0.700 ;
        RECT 49.985 0.300 49.995 0.700 ;
        RECT 49.995 0.310 50.005 0.700 ;
        RECT 50.005 0.320 50.015 0.700 ;
        RECT 50.015 0.330 50.025 0.700 ;
        RECT 50.025 0.340 50.035 0.700 ;
        RECT 50.035 0.350 50.045 0.700 ;
        RECT 50.045 0.360 50.055 0.700 ;
        RECT 50.055 0.370 50.065 0.700 ;
        RECT 50.065 0.380 50.075 0.700 ;
        RECT 50.075 0.390 50.085 0.700 ;
        RECT 50.085 0.400 50.095 0.700 ;
        RECT 50.095 0.410 50.105 0.700 ;
        RECT 50.105 0.420 50.115 0.700 ;
        RECT 50.115 0.430 50.125 0.700 ;
        RECT 50.125 0.440 50.135 0.700 ;
        RECT 50.135 0.450 50.145 0.700 ;
        RECT 50.145 0.460 50.155 0.700 ;
        RECT 50.155 0.470 50.165 0.700 ;
        RECT 50.165 0.480 50.175 0.700 ;
        RECT 50.175 0.490 50.185 0.700 ;
        RECT 50.185 0.500 50.195 0.700 ;
        RECT 50.195 0.510 50.205 0.700 ;
        RECT 50.205 0.520 50.215 0.700 ;
        RECT 50.215 0.530 50.225 0.700 ;
        RECT 50.225 0.540 50.235 0.700 ;
        RECT 50.235 0.550 50.245 0.700 ;
        RECT 50.245 0.560 50.255 0.700 ;
        RECT 50.255 0.570 50.265 0.700 ;
        RECT 47.415 0.570 47.425 0.700 ;
        RECT 47.425 0.560 47.435 0.700 ;
        RECT 47.435 0.550 47.445 0.700 ;
        RECT 47.445 0.540 47.455 0.700 ;
        RECT 47.455 0.530 47.465 0.700 ;
        RECT 47.465 0.520 47.475 0.700 ;
        RECT 47.475 0.510 47.485 0.700 ;
        RECT 47.485 0.500 47.495 0.700 ;
        RECT 47.495 0.490 47.505 0.700 ;
        RECT 47.505 0.480 47.515 0.700 ;
        RECT 47.515 0.470 47.525 0.700 ;
        RECT 47.525 0.460 47.535 0.700 ;
        RECT 47.535 0.450 47.545 0.700 ;
        RECT 47.545 0.440 47.555 0.700 ;
        RECT 47.555 0.430 47.565 0.700 ;
        RECT 47.565 0.420 47.575 0.700 ;
        RECT 47.575 0.410 47.585 0.700 ;
        RECT 47.585 0.400 47.595 0.700 ;
        RECT 47.595 0.390 47.605 0.700 ;
        RECT 47.605 0.380 47.615 0.700 ;
        RECT 47.615 0.370 47.625 0.700 ;
        RECT 47.625 0.360 47.635 0.700 ;
        RECT 47.635 0.350 47.645 0.700 ;
        RECT 47.645 0.340 47.655 0.700 ;
        RECT 47.655 0.330 47.665 0.700 ;
        RECT 47.665 0.320 47.675 0.700 ;
        RECT 47.675 0.310 47.685 0.700 ;
        RECT 47.685 0.300 47.695 0.700 ;
        RECT 47.695 0.290 47.705 0.700 ;
        RECT 47.705 0.280 47.715 0.700 ;
        RECT 47.715 0.270 47.725 0.700 ;
        RECT 47.725 0.260 47.735 0.700 ;
        RECT 47.735 0.250 47.745 0.700 ;
        RECT 47.745 0.240 47.755 0.700 ;
        RECT 47.755 0.230 47.765 0.700 ;
        RECT 47.765 0.220 47.775 0.700 ;
        RECT 47.775 0.210 47.785 0.700 ;
        RECT 47.785 0.200 47.795 0.700 ;
        RECT 47.795 0.190 47.805 0.700 ;
        RECT 47.805 0.180 47.815 0.700 ;
        RECT 47.815 0.170 47.825 0.700 ;
        RECT 47.825 0.160 47.835 0.700 ;
        RECT 47.835 0.150 47.845 0.700 ;
        RECT 47.845 0.140 47.855 0.700 ;
        RECT 47.855 0.130 47.865 0.700 ;
        RECT 47.865 0.120 47.875 0.700 ;
        RECT 47.875 0.110 47.885 0.700 ;
        RECT 47.885 0.100 47.895 0.700 ;
        RECT 47.895 0.090 47.905 0.700 ;
        RECT 47.905 0.080 49.775 0.700 ;
        RECT 56.195 0.090 56.205 0.700 ;
        RECT 56.205 0.100 56.215 0.700 ;
        RECT 56.215 0.110 56.225 0.700 ;
        RECT 56.225 0.120 56.235 0.700 ;
        RECT 56.235 0.130 56.245 0.700 ;
        RECT 56.245 0.140 56.255 0.700 ;
        RECT 56.255 0.150 56.265 0.700 ;
        RECT 56.265 0.160 56.275 0.700 ;
        RECT 56.275 0.170 56.285 0.700 ;
        RECT 56.285 0.180 56.295 0.700 ;
        RECT 56.295 0.190 56.305 0.700 ;
        RECT 56.305 0.200 56.315 0.700 ;
        RECT 56.315 0.210 56.325 0.700 ;
        RECT 56.325 0.220 56.335 0.700 ;
        RECT 56.335 0.230 56.345 0.700 ;
        RECT 56.345 0.240 56.355 0.700 ;
        RECT 56.355 0.250 56.365 0.700 ;
        RECT 56.365 0.260 56.375 0.700 ;
        RECT 56.375 0.270 56.385 0.700 ;
        RECT 56.385 0.280 56.395 0.700 ;
        RECT 56.395 0.290 56.405 0.700 ;
        RECT 56.405 0.300 56.415 0.700 ;
        RECT 56.415 0.310 56.425 0.700 ;
        RECT 56.425 0.320 56.435 0.700 ;
        RECT 56.435 0.330 56.445 0.700 ;
        RECT 56.445 0.340 56.455 0.700 ;
        RECT 56.455 0.350 56.465 0.700 ;
        RECT 56.465 0.360 56.475 0.700 ;
        RECT 56.475 0.370 56.485 0.700 ;
        RECT 56.485 0.380 56.495 0.700 ;
        RECT 56.495 0.390 56.505 0.700 ;
        RECT 56.505 0.400 56.515 0.700 ;
        RECT 56.515 0.410 56.525 0.700 ;
        RECT 56.525 0.420 56.535 0.700 ;
        RECT 56.535 0.430 56.545 0.700 ;
        RECT 56.545 0.440 56.555 0.700 ;
        RECT 56.555 0.450 56.565 0.700 ;
        RECT 56.565 0.460 56.575 0.700 ;
        RECT 56.575 0.470 56.585 0.700 ;
        RECT 56.585 0.480 56.595 0.700 ;
        RECT 56.595 0.490 56.605 0.700 ;
        RECT 56.605 0.500 56.615 0.700 ;
        RECT 56.615 0.510 56.625 0.700 ;
        RECT 56.625 0.520 56.635 0.700 ;
        RECT 56.635 0.530 56.645 0.700 ;
        RECT 56.645 0.540 56.655 0.700 ;
        RECT 56.655 0.550 56.665 0.700 ;
        RECT 56.665 0.560 56.675 0.700 ;
        RECT 56.675 0.570 56.685 0.700 ;
        RECT 53.835 0.570 53.845 0.700 ;
        RECT 53.845 0.560 53.855 0.700 ;
        RECT 53.855 0.550 53.865 0.700 ;
        RECT 53.865 0.540 53.875 0.700 ;
        RECT 53.875 0.530 53.885 0.700 ;
        RECT 53.885 0.520 53.895 0.700 ;
        RECT 53.895 0.510 53.905 0.700 ;
        RECT 53.905 0.500 53.915 0.700 ;
        RECT 53.915 0.490 53.925 0.700 ;
        RECT 53.925 0.480 53.935 0.700 ;
        RECT 53.935 0.470 53.945 0.700 ;
        RECT 53.945 0.460 53.955 0.700 ;
        RECT 53.955 0.450 53.965 0.700 ;
        RECT 53.965 0.440 53.975 0.700 ;
        RECT 53.975 0.430 53.985 0.700 ;
        RECT 53.985 0.420 53.995 0.700 ;
        RECT 53.995 0.410 54.005 0.700 ;
        RECT 54.005 0.400 54.015 0.700 ;
        RECT 54.015 0.390 54.025 0.700 ;
        RECT 54.025 0.380 54.035 0.700 ;
        RECT 54.035 0.370 54.045 0.700 ;
        RECT 54.045 0.360 54.055 0.700 ;
        RECT 54.055 0.350 54.065 0.700 ;
        RECT 54.065 0.340 54.075 0.700 ;
        RECT 54.075 0.330 54.085 0.700 ;
        RECT 54.085 0.320 54.095 0.700 ;
        RECT 54.095 0.310 54.105 0.700 ;
        RECT 54.105 0.300 54.115 0.700 ;
        RECT 54.115 0.290 54.125 0.700 ;
        RECT 54.125 0.280 54.135 0.700 ;
        RECT 54.135 0.270 54.145 0.700 ;
        RECT 54.145 0.260 54.155 0.700 ;
        RECT 54.155 0.250 54.165 0.700 ;
        RECT 54.165 0.240 54.175 0.700 ;
        RECT 54.175 0.230 54.185 0.700 ;
        RECT 54.185 0.220 54.195 0.700 ;
        RECT 54.195 0.210 54.205 0.700 ;
        RECT 54.205 0.200 54.215 0.700 ;
        RECT 54.215 0.190 54.225 0.700 ;
        RECT 54.225 0.180 54.235 0.700 ;
        RECT 54.235 0.170 54.245 0.700 ;
        RECT 54.245 0.160 54.255 0.700 ;
        RECT 54.255 0.150 54.265 0.700 ;
        RECT 54.265 0.140 54.275 0.700 ;
        RECT 54.275 0.130 54.285 0.700 ;
        RECT 54.285 0.120 54.295 0.700 ;
        RECT 54.295 0.110 54.305 0.700 ;
        RECT 54.305 0.100 54.315 0.700 ;
        RECT 54.315 0.090 54.325 0.700 ;
        RECT 54.325 0.080 56.195 0.700 ;
        RECT 62.615 0.090 62.625 0.700 ;
        RECT 62.625 0.100 62.635 0.700 ;
        RECT 62.635 0.110 62.645 0.700 ;
        RECT 62.645 0.120 62.655 0.700 ;
        RECT 62.655 0.130 62.665 0.700 ;
        RECT 62.665 0.140 62.675 0.700 ;
        RECT 62.675 0.150 62.685 0.700 ;
        RECT 62.685 0.160 62.695 0.700 ;
        RECT 62.695 0.170 62.705 0.700 ;
        RECT 62.705 0.180 62.715 0.700 ;
        RECT 62.715 0.190 62.725 0.700 ;
        RECT 62.725 0.200 62.735 0.700 ;
        RECT 62.735 0.210 62.745 0.700 ;
        RECT 62.745 0.220 62.755 0.700 ;
        RECT 62.755 0.230 62.765 0.700 ;
        RECT 62.765 0.240 62.775 0.700 ;
        RECT 62.775 0.250 62.785 0.700 ;
        RECT 62.785 0.260 62.795 0.700 ;
        RECT 62.795 0.270 62.805 0.700 ;
        RECT 62.805 0.280 62.815 0.700 ;
        RECT 62.815 0.290 62.825 0.700 ;
        RECT 62.825 0.300 62.835 0.700 ;
        RECT 62.835 0.310 62.845 0.700 ;
        RECT 62.845 0.320 62.855 0.700 ;
        RECT 62.855 0.330 62.865 0.700 ;
        RECT 62.865 0.340 62.875 0.700 ;
        RECT 62.875 0.350 62.885 0.700 ;
        RECT 62.885 0.360 62.895 0.700 ;
        RECT 62.895 0.370 62.905 0.700 ;
        RECT 62.905 0.380 62.915 0.700 ;
        RECT 62.915 0.390 62.925 0.700 ;
        RECT 62.925 0.400 62.935 0.700 ;
        RECT 62.935 0.410 62.945 0.700 ;
        RECT 62.945 0.420 62.955 0.700 ;
        RECT 62.955 0.430 62.965 0.700 ;
        RECT 62.965 0.440 62.975 0.700 ;
        RECT 62.975 0.450 62.985 0.700 ;
        RECT 62.985 0.460 62.995 0.700 ;
        RECT 62.995 0.470 63.005 0.700 ;
        RECT 63.005 0.480 63.015 0.700 ;
        RECT 63.015 0.490 63.025 0.700 ;
        RECT 63.025 0.500 63.035 0.700 ;
        RECT 63.035 0.510 63.045 0.700 ;
        RECT 63.045 0.520 63.055 0.700 ;
        RECT 63.055 0.530 63.065 0.700 ;
        RECT 63.065 0.540 63.075 0.700 ;
        RECT 63.075 0.550 63.085 0.700 ;
        RECT 63.085 0.560 63.095 0.700 ;
        RECT 63.095 0.570 63.105 0.700 ;
        RECT 60.255 0.570 60.265 0.700 ;
        RECT 60.265 0.560 60.275 0.700 ;
        RECT 60.275 0.550 60.285 0.700 ;
        RECT 60.285 0.540 60.295 0.700 ;
        RECT 60.295 0.530 60.305 0.700 ;
        RECT 60.305 0.520 60.315 0.700 ;
        RECT 60.315 0.510 60.325 0.700 ;
        RECT 60.325 0.500 60.335 0.700 ;
        RECT 60.335 0.490 60.345 0.700 ;
        RECT 60.345 0.480 60.355 0.700 ;
        RECT 60.355 0.470 60.365 0.700 ;
        RECT 60.365 0.460 60.375 0.700 ;
        RECT 60.375 0.450 60.385 0.700 ;
        RECT 60.385 0.440 60.395 0.700 ;
        RECT 60.395 0.430 60.405 0.700 ;
        RECT 60.405 0.420 60.415 0.700 ;
        RECT 60.415 0.410 60.425 0.700 ;
        RECT 60.425 0.400 60.435 0.700 ;
        RECT 60.435 0.390 60.445 0.700 ;
        RECT 60.445 0.380 60.455 0.700 ;
        RECT 60.455 0.370 60.465 0.700 ;
        RECT 60.465 0.360 60.475 0.700 ;
        RECT 60.475 0.350 60.485 0.700 ;
        RECT 60.485 0.340 60.495 0.700 ;
        RECT 60.495 0.330 60.505 0.700 ;
        RECT 60.505 0.320 60.515 0.700 ;
        RECT 60.515 0.310 60.525 0.700 ;
        RECT 60.525 0.300 60.535 0.700 ;
        RECT 60.535 0.290 60.545 0.700 ;
        RECT 60.545 0.280 60.555 0.700 ;
        RECT 60.555 0.270 60.565 0.700 ;
        RECT 60.565 0.260 60.575 0.700 ;
        RECT 60.575 0.250 60.585 0.700 ;
        RECT 60.585 0.240 60.595 0.700 ;
        RECT 60.595 0.230 60.605 0.700 ;
        RECT 60.605 0.220 60.615 0.700 ;
        RECT 60.615 0.210 60.625 0.700 ;
        RECT 60.625 0.200 60.635 0.700 ;
        RECT 60.635 0.190 60.645 0.700 ;
        RECT 60.645 0.180 60.655 0.700 ;
        RECT 60.655 0.170 60.665 0.700 ;
        RECT 60.665 0.160 60.675 0.700 ;
        RECT 60.675 0.150 60.685 0.700 ;
        RECT 60.685 0.140 60.695 0.700 ;
        RECT 60.695 0.130 60.705 0.700 ;
        RECT 60.705 0.120 60.715 0.700 ;
        RECT 60.715 0.110 60.725 0.700 ;
        RECT 60.725 0.100 60.735 0.700 ;
        RECT 60.735 0.090 60.745 0.700 ;
        RECT 60.745 0.080 62.615 0.700 ;
        RECT 69.035 0.090 69.045 0.700 ;
        RECT 69.045 0.100 69.055 0.700 ;
        RECT 69.055 0.110 69.065 0.700 ;
        RECT 69.065 0.120 69.075 0.700 ;
        RECT 69.075 0.130 69.085 0.700 ;
        RECT 69.085 0.140 69.095 0.700 ;
        RECT 69.095 0.150 69.105 0.700 ;
        RECT 69.105 0.160 69.115 0.700 ;
        RECT 69.115 0.170 69.125 0.700 ;
        RECT 69.125 0.180 69.135 0.700 ;
        RECT 69.135 0.190 69.145 0.700 ;
        RECT 69.145 0.200 69.155 0.700 ;
        RECT 69.155 0.210 69.165 0.700 ;
        RECT 69.165 0.220 69.175 0.700 ;
        RECT 69.175 0.230 69.185 0.700 ;
        RECT 69.185 0.240 69.195 0.700 ;
        RECT 69.195 0.250 69.205 0.700 ;
        RECT 69.205 0.260 69.215 0.700 ;
        RECT 69.215 0.270 69.225 0.700 ;
        RECT 69.225 0.280 69.235 0.700 ;
        RECT 69.235 0.290 69.245 0.700 ;
        RECT 69.245 0.300 69.255 0.700 ;
        RECT 69.255 0.310 69.265 0.700 ;
        RECT 69.265 0.320 69.275 0.700 ;
        RECT 69.275 0.330 69.285 0.700 ;
        RECT 69.285 0.340 69.295 0.700 ;
        RECT 69.295 0.350 69.305 0.700 ;
        RECT 69.305 0.360 69.315 0.700 ;
        RECT 69.315 0.370 69.325 0.700 ;
        RECT 69.325 0.380 69.335 0.700 ;
        RECT 69.335 0.390 69.345 0.700 ;
        RECT 69.345 0.400 69.355 0.700 ;
        RECT 69.355 0.410 69.365 0.700 ;
        RECT 69.365 0.420 69.375 0.700 ;
        RECT 69.375 0.430 69.385 0.700 ;
        RECT 69.385 0.440 69.395 0.700 ;
        RECT 69.395 0.450 69.405 0.700 ;
        RECT 69.405 0.460 69.415 0.700 ;
        RECT 69.415 0.470 69.425 0.700 ;
        RECT 69.425 0.480 69.435 0.700 ;
        RECT 69.435 0.490 69.445 0.700 ;
        RECT 69.445 0.500 69.455 0.700 ;
        RECT 69.455 0.510 69.465 0.700 ;
        RECT 69.465 0.520 69.475 0.700 ;
        RECT 69.475 0.530 69.485 0.700 ;
        RECT 69.485 0.540 69.495 0.700 ;
        RECT 69.495 0.550 69.505 0.700 ;
        RECT 69.505 0.560 69.515 0.700 ;
        RECT 69.515 0.570 69.525 0.700 ;
        RECT 66.675 0.570 66.685 0.700 ;
        RECT 66.685 0.560 66.695 0.700 ;
        RECT 66.695 0.550 66.705 0.700 ;
        RECT 66.705 0.540 66.715 0.700 ;
        RECT 66.715 0.530 66.725 0.700 ;
        RECT 66.725 0.520 66.735 0.700 ;
        RECT 66.735 0.510 66.745 0.700 ;
        RECT 66.745 0.500 66.755 0.700 ;
        RECT 66.755 0.490 66.765 0.700 ;
        RECT 66.765 0.480 66.775 0.700 ;
        RECT 66.775 0.470 66.785 0.700 ;
        RECT 66.785 0.460 66.795 0.700 ;
        RECT 66.795 0.450 66.805 0.700 ;
        RECT 66.805 0.440 66.815 0.700 ;
        RECT 66.815 0.430 66.825 0.700 ;
        RECT 66.825 0.420 66.835 0.700 ;
        RECT 66.835 0.410 66.845 0.700 ;
        RECT 66.845 0.400 66.855 0.700 ;
        RECT 66.855 0.390 66.865 0.700 ;
        RECT 66.865 0.380 66.875 0.700 ;
        RECT 66.875 0.370 66.885 0.700 ;
        RECT 66.885 0.360 66.895 0.700 ;
        RECT 66.895 0.350 66.905 0.700 ;
        RECT 66.905 0.340 66.915 0.700 ;
        RECT 66.915 0.330 66.925 0.700 ;
        RECT 66.925 0.320 66.935 0.700 ;
        RECT 66.935 0.310 66.945 0.700 ;
        RECT 66.945 0.300 66.955 0.700 ;
        RECT 66.955 0.290 66.965 0.700 ;
        RECT 66.965 0.280 66.975 0.700 ;
        RECT 66.975 0.270 66.985 0.700 ;
        RECT 66.985 0.260 66.995 0.700 ;
        RECT 66.995 0.250 67.005 0.700 ;
        RECT 67.005 0.240 67.015 0.700 ;
        RECT 67.015 0.230 67.025 0.700 ;
        RECT 67.025 0.220 67.035 0.700 ;
        RECT 67.035 0.210 67.045 0.700 ;
        RECT 67.045 0.200 67.055 0.700 ;
        RECT 67.055 0.190 67.065 0.700 ;
        RECT 67.065 0.180 67.075 0.700 ;
        RECT 67.075 0.170 67.085 0.700 ;
        RECT 67.085 0.160 67.095 0.700 ;
        RECT 67.095 0.150 67.105 0.700 ;
        RECT 67.105 0.140 67.115 0.700 ;
        RECT 67.115 0.130 67.125 0.700 ;
        RECT 67.125 0.120 67.135 0.700 ;
        RECT 67.135 0.110 67.145 0.700 ;
        RECT 67.145 0.100 67.155 0.700 ;
        RECT 67.155 0.090 67.165 0.700 ;
        RECT 67.165 0.080 69.035 0.700 ;
        RECT 1.100 1.100 70.900 187.900 ;
        RECT 71.300 71.440 71.555 78.100 ;
        RECT 71.300 63.270 71.555 68.270 ;
        RECT 71.300 51.630 71.555 59.770 ;
        RECT 71.300 39.130 71.555 48.130 ;
        RECT 71.300 26.270 71.555 35.270 ;
        RECT 71.300 14.630 71.555 22.770 ;
        RECT 71.300 3.610 71.555 11.130 ;
        RECT 70.725 0.040 71.555 0.700 ;
        RECT 71.300 0.040 71.555 2.960 ;
      LAYER M1 ;
        RECT 1.100 1.100 70.900 187.900 ;
        RECT 0.000 0.000 72.000 0.400 ;
        RECT 0.000 0.000 1.800 0.700 ;
        RECT 70.200 0.000 72.000 0.700 ;
        RECT 0.000 0.000 0.700 78.100 ;
        RECT 71.300 0.000 72.000 78.100 ;
      LAYER M3 ;
        RECT 0.560 0.120 1.275 0.700 ;
        RECT 0.560 0.120 0.700 78.100 ;
        RECT 1.100 1.100 70.900 187.900 ;
        RECT 70.725 0.120 71.455 0.700 ;
        RECT 71.300 0.120 71.455 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 70.900 187.900 ;
        RECT 71.300 185.015 72.000 187.775 ;
        RECT 71.300 177.615 72.000 184.415 ;
        RECT 71.300 170.640 72.000 176.940 ;
        RECT 71.300 162.140 72.000 170.040 ;
        RECT 71.300 154.840 72.000 161.540 ;
        RECT 71.300 139.530 72.000 150.030 ;
        RECT 71.300 127.890 72.000 136.030 ;
        RECT 71.300 116.930 72.000 124.390 ;
        RECT 71.300 105.930 72.000 113.930 ;
        RECT 71.300 94.290 72.000 102.430 ;
        RECT 71.300 90.340 72.000 92.340 ;
        RECT 71.300 85.080 72.000 87.960 ;
        RECT 71.300 79.590 72.000 84.480 ;
        RECT 71.300 71.440 72.000 79.110 ;
        RECT 71.300 57.770 72.000 68.270 ;
        RECT 71.300 45.630 72.000 54.270 ;
        RECT 71.300 32.770 72.000 42.130 ;
        RECT 71.300 20.470 72.000 28.910 ;
        RECT 71.300 9.130 72.000 16.970 ;
        RECT 71.300 3.610 72.000 5.630 ;
        RECT 0.000 0.000 72.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 71.300 0.000 72.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 70.900 187.900 ;
        RECT 71.300 185.400 72.000 187.775 ;
        RECT 71.300 177.615 72.000 184.955 ;
        RECT 71.300 170.640 72.000 176.940 ;
        RECT 71.300 162.140 72.000 170.040 ;
        RECT 71.300 154.840 72.000 161.540 ;
        RECT 71.300 145.030 72.000 150.030 ;
        RECT 71.300 133.390 72.000 141.530 ;
        RECT 71.300 122.170 72.000 129.890 ;
        RECT 71.300 111.430 72.000 119.170 ;
        RECT 71.300 99.790 72.000 107.930 ;
        RECT 71.300 90.340 72.000 96.290 ;
        RECT 71.300 85.080 72.000 87.960 ;
        RECT 71.300 79.590 72.000 84.780 ;
        RECT 71.300 71.440 72.000 79.110 ;
        RECT 71.300 63.270 72.000 68.270 ;
        RECT 71.300 51.630 72.000 59.770 ;
        RECT 71.300 39.130 72.000 48.130 ;
        RECT 71.300 26.270 72.000 35.270 ;
        RECT 71.300 14.630 72.000 22.770 ;
        RECT 71.300 3.610 72.000 11.130 ;
        RECT 0.000 0.000 72.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 71.300 0.000 72.000 2.960 ;
      LAYER M2 ;
        RECT 0.000 0.000 0.925 0.700 ;
        RECT 0.000 0.000 0.700 78.100 ;
        RECT 1.100 1.100 70.900 187.900 ;
        RECT 71.040 0.000 72.000 0.700 ;
        RECT 71.300 0.000 72.000 78.100 ;
  END 
END PSESDCLAMP

MACRO PSSPLIT_OSC
  CLASS  PAD ;
  FOREIGN PSSPLIT_OSC 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 1.320 0.000 6.540 0.700 ;
        RECT 33.460 0.000 38.680 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
      LAYER M1 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 162.140 40.000 170.040 ;
      LAYER M3 ;
        RECT 1.320 0.000 6.540 0.700 ;
        RECT 33.460 0.000 38.680 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 170.640 0.700 184.415 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 0.000 5.995 0.700 ;
        RECT 0.000 0.000 0.700 79.110 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 170.640 40.000 184.415 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 34.005 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 79.110 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 170.635 0.700 184.955 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 0.000 5.995 0.700 ;
        RECT 0.000 0.000 0.700 79.110 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 170.635 40.000 184.955 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 34.005 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 79.110 ;
      LAYER M2 ;
        RECT 1.100 1.100 38.900 187.900 ;
  END 
END PSSPLIT_OSC

MACRO PSCORNER
  CLASS  ENDCAP BOTTOMLEFT ;
  FOREIGN PSCORNER 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 189.000 BY 189.000 ;
  SYMMETRY Y R90  ;
  SITE CornerSite ;
  OBS 
      LAYER M4 ;
        RECT 108.345 0.000 188.400 188.895 ;
        RECT 0.000 108.420 188.895 188.400 ;
        RECT 0.105 0.105 188.895 188.895 ;
      LAYER M1 ;
        RECT 108.345 0.000 188.400 188.915 ;
        RECT 0.000 108.420 188.915 188.400 ;
        RECT 0.085 0.085 188.915 188.915 ;
      LAYER M3 ;
        RECT 108.345 0.000 188.400 188.895 ;
        RECT 0.000 108.420 188.895 188.400 ;
        RECT 0.105 0.105 188.895 188.895 ;
      LAYER M6 ;
        RECT 108.345 0.000 189.000 2.960 ;
        RECT 0.230 0.230 189.000 2.960 ;
        RECT 0.230 3.610 189.000 5.630 ;
        RECT 0.230 9.130 189.000 16.970 ;
        RECT 0.230 20.470 189.000 28.910 ;
        RECT 0.230 32.770 189.000 42.130 ;
        RECT 0.230 45.630 189.000 54.270 ;
        RECT 0.230 57.770 189.000 68.270 ;
        RECT 0.230 71.440 189.000 79.110 ;
        RECT 0.230 79.590 189.000 84.480 ;
        RECT 0.230 85.080 189.000 87.960 ;
        RECT 0.230 90.340 189.000 92.340 ;
        RECT 0.230 94.290 189.000 102.430 ;
        RECT 0.230 0.230 188.770 188.770 ;
        RECT 0.230 105.930 189.000 113.930 ;
        RECT 0.000 108.420 189.000 113.930 ;
        RECT 0.000 116.930 189.000 124.390 ;
        RECT 0.000 127.890 189.000 136.030 ;
        RECT 0.000 139.530 189.000 150.030 ;
        RECT 0.000 154.840 189.000 161.540 ;
        RECT 0.000 162.140 189.000 170.040 ;
        RECT 0.000 170.640 189.000 176.940 ;
        RECT 0.000 177.615 189.000 184.415 ;
        RECT 0.000 185.015 189.000 187.775 ;
        RECT 108.345 0.000 188.770 188.770 ;
        RECT 0.000 108.420 188.770 188.770 ;
        RECT 0.230 0.230 2.960 189.000 ;
        RECT 0.000 108.420 2.960 189.000 ;
        RECT 3.610 0.230 5.630 189.000 ;
        RECT 9.130 0.230 16.970 189.000 ;
        RECT 20.470 0.230 28.910 189.000 ;
        RECT 32.770 0.230 42.130 189.000 ;
        RECT 45.630 0.230 54.270 189.000 ;
        RECT 57.770 0.230 68.270 189.000 ;
        RECT 71.440 0.230 79.110 189.000 ;
        RECT 79.590 0.230 84.480 189.000 ;
        RECT 85.080 0.230 87.960 189.000 ;
        RECT 90.340 0.230 92.340 189.000 ;
        RECT 94.290 0.230 102.430 189.000 ;
        RECT 108.345 0.000 113.930 189.000 ;
        RECT 105.930 0.230 113.930 189.000 ;
        RECT 116.930 0.000 124.390 189.000 ;
        RECT 127.890 0.000 136.030 189.000 ;
        RECT 139.530 0.000 150.030 189.000 ;
        RECT 154.840 0.000 161.540 189.000 ;
        RECT 162.140 0.000 170.040 189.000 ;
        RECT 170.640 0.000 176.940 189.000 ;
        RECT 177.615 0.000 184.415 189.000 ;
        RECT 185.015 0.000 187.775 189.000 ;
      LAYER M5 ;
        RECT 108.345 0.000 189.000 2.960 ;
        RECT 0.105 0.105 189.000 2.960 ;
        RECT 0.105 3.610 189.000 11.130 ;
        RECT 0.105 14.630 189.000 22.770 ;
        RECT 0.105 26.270 189.000 35.270 ;
        RECT 0.105 39.130 189.000 48.130 ;
        RECT 0.105 51.630 189.000 59.770 ;
        RECT 0.105 63.270 189.000 68.270 ;
        RECT 0.105 71.440 189.000 79.110 ;
        RECT 0.105 79.590 189.000 84.780 ;
        RECT 0.105 85.080 189.000 87.960 ;
        RECT 0.105 90.340 189.000 96.290 ;
        RECT 0.105 99.790 189.000 107.930 ;
        RECT 0.105 0.105 188.895 188.895 ;
        RECT 0.000 111.430 189.000 119.170 ;
        RECT 0.000 122.170 189.000 129.890 ;
        RECT 0.000 133.390 189.000 141.530 ;
        RECT 0.000 145.030 189.000 150.030 ;
        RECT 0.000 154.840 189.000 161.540 ;
        RECT 0.000 162.140 189.000 170.040 ;
        RECT 0.000 170.640 189.000 176.940 ;
        RECT 0.000 177.615 189.000 184.955 ;
        RECT 0.000 185.400 189.000 187.775 ;
        RECT 108.345 0.000 188.895 188.895 ;
        RECT 0.000 108.420 188.895 188.895 ;
        RECT 0.105 0.105 2.960 189.000 ;
        RECT 0.000 108.420 2.960 189.000 ;
        RECT 3.610 0.105 11.130 189.000 ;
        RECT 14.630 0.105 22.770 189.000 ;
        RECT 26.270 0.105 35.270 189.000 ;
        RECT 39.130 0.105 48.130 189.000 ;
        RECT 51.630 0.105 59.770 189.000 ;
        RECT 63.270 0.105 68.270 189.000 ;
        RECT 71.440 0.105 79.110 189.000 ;
        RECT 79.590 0.105 84.780 189.000 ;
        RECT 85.080 0.105 87.960 189.000 ;
        RECT 90.340 0.105 96.290 189.000 ;
        RECT 99.790 0.105 107.930 189.000 ;
        RECT 111.430 0.000 119.170 189.000 ;
        RECT 122.170 0.000 129.890 189.000 ;
        RECT 133.390 0.000 141.530 189.000 ;
        RECT 145.030 0.000 150.030 189.000 ;
        RECT 154.840 0.000 161.540 189.000 ;
        RECT 162.140 0.000 170.040 189.000 ;
        RECT 170.640 0.000 176.940 189.000 ;
        RECT 177.615 0.000 184.955 189.000 ;
        RECT 185.400 0.000 187.775 189.000 ;
      LAYER M2 ;
        RECT 108.345 0.000 188.400 188.950 ;
        RECT 0.050 86.045 189.000 89.040 ;
        RECT 0.000 108.420 188.950 188.400 ;
        RECT 0.050 0.050 188.950 188.950 ;
  END 
END PSCORNER

MACRO PSVSSO
  CLASS  PAD ;
  FOREIGN PSVSSO 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN VSSO
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 4.210 188.300 35.790 189.000 ;
      LAYER V3 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M3 ;
        RECT 4.210 188.300 35.790 189.000 ;
      LAYER V2 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M2 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V1 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M1 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER M6 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V5 ;
        RECT 4.555 188.510 4.915 188.870 ;
        RECT 5.265 188.510 5.625 188.870 ;
        RECT 5.975 188.510 6.335 188.870 ;
        RECT 6.685 188.510 7.045 188.870 ;
        RECT 7.395 188.510 7.755 188.870 ;
        RECT 8.105 188.510 8.465 188.870 ;
        RECT 8.815 188.510 9.175 188.870 ;
        RECT 9.525 188.510 9.885 188.870 ;
        RECT 10.235 188.510 10.595 188.870 ;
        RECT 10.945 188.510 11.305 188.870 ;
        RECT 11.655 188.510 12.015 188.870 ;
        RECT 12.365 188.510 12.725 188.870 ;
        RECT 13.075 188.510 13.435 188.870 ;
        RECT 13.785 188.510 14.145 188.870 ;
        RECT 14.495 188.510 14.855 188.870 ;
        RECT 15.205 188.510 15.565 188.870 ;
        RECT 15.915 188.510 16.275 188.870 ;
        RECT 16.625 188.510 16.985 188.870 ;
        RECT 17.335 188.510 17.695 188.870 ;
        RECT 18.045 188.510 18.405 188.870 ;
        RECT 18.755 188.510 19.115 188.870 ;
        RECT 19.465 188.510 19.825 188.870 ;
        RECT 20.175 188.510 20.535 188.870 ;
        RECT 20.885 188.510 21.245 188.870 ;
        RECT 21.595 188.510 21.955 188.870 ;
        RECT 22.305 188.510 22.665 188.870 ;
        RECT 23.015 188.510 23.375 188.870 ;
        RECT 23.725 188.510 24.085 188.870 ;
        RECT 24.435 188.510 24.795 188.870 ;
        RECT 25.145 188.510 25.505 188.870 ;
        RECT 25.855 188.510 26.215 188.870 ;
        RECT 26.565 188.510 26.925 188.870 ;
        RECT 27.275 188.510 27.635 188.870 ;
        RECT 27.985 188.510 28.345 188.870 ;
        RECT 28.695 188.510 29.055 188.870 ;
        RECT 29.405 188.510 29.765 188.870 ;
        RECT 30.115 188.510 30.475 188.870 ;
        RECT 30.825 188.510 31.185 188.870 ;
        RECT 31.535 188.510 31.895 188.870 ;
        RECT 32.245 188.510 32.605 188.870 ;
        RECT 32.955 188.510 33.315 188.870 ;
        RECT 33.665 188.510 34.025 188.870 ;
        RECT 34.375 188.510 34.735 188.870 ;
        RECT 35.085 188.510 35.445 188.870 ;
      LAYER M5 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V4 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
    END
  END VSSO
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.700 187.720 ;
        RECT 0.130 177.560 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.885 ;
        RECT 0.130 162.085 0.700 170.040 ;
        RECT 0.130 154.785 0.700 160.610 ;
        RECT 0.130 86.045 0.700 87.905 ;
        RECT 0.130 79.535 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 74.280 ;
        RECT 0.000 0.000 0.345 78.095 ;
        RECT 0.000 77.765 0.700 78.095 ;
        RECT 4.680 0.000 10.595 0.700 ;
        RECT 12.895 0.000 18.815 0.700 ;
        RECT 21.150 0.000 27.070 0.700 ;
        RECT 29.405 0.000 35.325 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.720 ;
        RECT 39.300 177.560 39.870 184.900 ;
        RECT 39.300 171.540 39.870 176.885 ;
        RECT 39.300 162.140 39.870 169.985 ;
        RECT 39.300 154.840 39.870 160.555 ;
        RECT 39.300 86.045 39.870 87.905 ;
        RECT 39.300 79.535 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 74.280 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.700 187.775 ;
        RECT 0.000 177.565 0.700 184.480 ;
        RECT 0.000 171.540 0.700 176.885 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 40.000 187.775 ;
        RECT 39.300 177.565 40.000 184.480 ;
        RECT 39.300 171.540 40.000 176.885 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 85.980 40.000 160.610 ;
        RECT 39.300 79.600 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 74.280 ;
        RECT 0.000 0.000 0.700 76.370 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 39.625 0.000 40.000 78.100 ;
        RECT 39.300 77.770 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.700 187.720 ;
        RECT 0.130 177.560 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.885 ;
        RECT 0.130 162.085 0.700 170.040 ;
        RECT 0.130 154.785 0.700 160.610 ;
        RECT 0.130 86.045 0.700 87.905 ;
        RECT 0.130 79.535 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 74.280 ;
        RECT 0.000 0.000 0.345 78.095 ;
        RECT 0.000 77.765 0.700 78.095 ;
        RECT 4.680 0.000 10.595 0.700 ;
        RECT 12.895 0.000 18.815 0.700 ;
        RECT 21.150 0.000 27.070 0.700 ;
        RECT 29.405 0.000 35.325 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.720 ;
        RECT 39.300 177.560 39.870 184.900 ;
        RECT 39.300 171.540 39.870 176.885 ;
        RECT 39.300 162.140 39.870 169.985 ;
        RECT 39.300 154.840 39.870 160.555 ;
        RECT 39.300 86.045 39.870 87.905 ;
        RECT 39.300 79.535 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 74.335 ;
        RECT 39.625 0.000 40.000 78.155 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.130 185.345 0.700 187.720 ;
        RECT 0.130 177.560 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.885 ;
        RECT 0.130 162.140 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 87.905 ;
        RECT 0.130 79.535 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.720 ;
        RECT 39.300 177.560 39.870 184.955 ;
        RECT 39.300 171.540 39.870 176.885 ;
        RECT 39.300 162.140 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 87.905 ;
        RECT 39.300 79.535 39.870 84.480 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 74.280 ;
        RECT 39.300 0.000 40.000 74.280 ;
        RECT 0.000 0.000 0.345 78.095 ;
        RECT 0.000 77.765 0.700 78.095 ;
        RECT 39.625 0.000 40.000 78.100 ;
  END 
END PSVSSO

MACRO PSVSSH
  CLASS  PAD ;
  FOREIGN PSVSSH 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN VSSH
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 4.210 188.300 35.790 189.000 ;
      LAYER V3 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M3 ;
        RECT 4.210 188.300 35.790 189.000 ;
      LAYER V2 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M2 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V1 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M1 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER M6 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V5 ;
        RECT 4.555 188.510 4.915 188.870 ;
        RECT 5.265 188.510 5.625 188.870 ;
        RECT 5.975 188.510 6.335 188.870 ;
        RECT 6.685 188.510 7.045 188.870 ;
        RECT 7.395 188.510 7.755 188.870 ;
        RECT 8.105 188.510 8.465 188.870 ;
        RECT 8.815 188.510 9.175 188.870 ;
        RECT 9.525 188.510 9.885 188.870 ;
        RECT 10.235 188.510 10.595 188.870 ;
        RECT 10.945 188.510 11.305 188.870 ;
        RECT 11.655 188.510 12.015 188.870 ;
        RECT 12.365 188.510 12.725 188.870 ;
        RECT 13.075 188.510 13.435 188.870 ;
        RECT 13.785 188.510 14.145 188.870 ;
        RECT 14.495 188.510 14.855 188.870 ;
        RECT 15.205 188.510 15.565 188.870 ;
        RECT 15.915 188.510 16.275 188.870 ;
        RECT 16.625 188.510 16.985 188.870 ;
        RECT 17.335 188.510 17.695 188.870 ;
        RECT 18.045 188.510 18.405 188.870 ;
        RECT 18.755 188.510 19.115 188.870 ;
        RECT 19.465 188.510 19.825 188.870 ;
        RECT 20.175 188.510 20.535 188.870 ;
        RECT 20.885 188.510 21.245 188.870 ;
        RECT 21.595 188.510 21.955 188.870 ;
        RECT 22.305 188.510 22.665 188.870 ;
        RECT 23.015 188.510 23.375 188.870 ;
        RECT 23.725 188.510 24.085 188.870 ;
        RECT 24.435 188.510 24.795 188.870 ;
        RECT 25.145 188.510 25.505 188.870 ;
        RECT 25.855 188.510 26.215 188.870 ;
        RECT 26.565 188.510 26.925 188.870 ;
        RECT 27.275 188.510 27.635 188.870 ;
        RECT 27.985 188.510 28.345 188.870 ;
        RECT 28.695 188.510 29.055 188.870 ;
        RECT 29.405 188.510 29.765 188.870 ;
        RECT 30.115 188.510 30.475 188.870 ;
        RECT 30.825 188.510 31.185 188.870 ;
        RECT 31.535 188.510 31.895 188.870 ;
        RECT 32.245 188.510 32.605 188.870 ;
        RECT 32.955 188.510 33.315 188.870 ;
        RECT 33.665 188.510 34.025 188.870 ;
        RECT 34.375 188.510 34.735 188.870 ;
        RECT 35.085 188.510 35.445 188.870 ;
      LAYER M5 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V4 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
    END
  END VSSH
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.700 187.720 ;
        RECT 0.130 177.560 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.885 ;
        RECT 0.130 162.085 0.700 170.040 ;
        RECT 0.130 154.785 0.700 160.610 ;
        RECT 0.130 86.045 0.700 87.905 ;
        RECT 0.130 79.535 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 74.280 ;
        RECT 0.000 0.000 0.345 78.095 ;
        RECT 0.000 77.765 0.700 78.095 ;
        RECT 4.680 0.000 10.595 0.700 ;
        RECT 12.895 0.000 18.815 0.700 ;
        RECT 21.150 0.000 27.070 0.700 ;
        RECT 29.405 0.000 35.325 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.720 ;
        RECT 39.300 177.560 39.870 184.900 ;
        RECT 39.300 171.540 39.870 176.885 ;
        RECT 39.300 162.140 39.870 169.985 ;
        RECT 39.300 154.840 39.870 160.555 ;
        RECT 39.300 86.045 39.870 87.905 ;
        RECT 39.300 79.535 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 74.280 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.700 187.775 ;
        RECT 0.000 177.565 0.700 184.480 ;
        RECT 0.000 171.540 0.700 176.885 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 40.000 187.775 ;
        RECT 39.300 177.565 40.000 184.480 ;
        RECT 39.300 171.540 40.000 176.885 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 85.980 40.000 160.610 ;
        RECT 39.300 79.600 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 74.280 ;
        RECT 0.000 0.000 0.700 76.370 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 39.625 0.000 40.000 78.100 ;
        RECT 39.300 77.770 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.700 187.720 ;
        RECT 0.130 177.560 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.885 ;
        RECT 0.130 162.085 0.700 170.040 ;
        RECT 0.130 154.785 0.700 160.610 ;
        RECT 0.130 86.045 0.700 87.905 ;
        RECT 0.130 79.535 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 74.280 ;
        RECT 0.000 0.000 0.345 78.095 ;
        RECT 0.000 77.765 0.700 78.095 ;
        RECT 4.680 0.000 10.595 0.700 ;
        RECT 12.895 0.000 18.815 0.700 ;
        RECT 21.150 0.000 27.070 0.700 ;
        RECT 29.405 0.000 35.325 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.720 ;
        RECT 39.300 177.560 39.870 184.900 ;
        RECT 39.300 171.540 39.870 176.885 ;
        RECT 39.300 162.140 39.870 169.985 ;
        RECT 39.300 154.840 39.870 160.555 ;
        RECT 39.300 86.045 39.870 87.905 ;
        RECT 39.300 79.535 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 74.335 ;
        RECT 39.625 0.000 40.000 78.155 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.130 185.345 0.700 187.720 ;
        RECT 0.130 177.560 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.885 ;
        RECT 0.130 162.140 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 87.905 ;
        RECT 0.130 79.535 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.720 ;
        RECT 39.300 177.560 39.870 184.955 ;
        RECT 39.300 171.540 39.870 176.885 ;
        RECT 39.300 162.140 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 87.905 ;
        RECT 39.300 79.535 39.870 84.480 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 74.280 ;
        RECT 39.300 0.000 40.000 74.280 ;
        RECT 0.000 0.000 0.345 78.095 ;
        RECT 0.000 77.765 0.700 78.095 ;
        RECT 39.625 0.000 40.000 78.100 ;
  END 
END PSVSSH

MACRO PSVSSC
  CLASS  PAD ;
  FOREIGN PSVSSC 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    CLASS CORE ;
      LAYER M4 ;
        RECT 12.895 0.000 18.815 0.700 ;
        RECT 4.210 188.300 35.790 189.000 ;
      LAYER V3 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M3 ;
        RECT 12.895 0.000 18.815 0.700 ;
        RECT 4.210 188.300 35.790 189.000 ;
      LAYER V2 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M2 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V1 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M1 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER M6 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V5 ;
        RECT 4.555 188.510 4.915 188.870 ;
        RECT 5.265 188.510 5.625 188.870 ;
        RECT 5.975 188.510 6.335 188.870 ;
        RECT 6.685 188.510 7.045 188.870 ;
        RECT 7.395 188.510 7.755 188.870 ;
        RECT 8.105 188.510 8.465 188.870 ;
        RECT 8.815 188.510 9.175 188.870 ;
        RECT 9.525 188.510 9.885 188.870 ;
        RECT 10.235 188.510 10.595 188.870 ;
        RECT 10.945 188.510 11.305 188.870 ;
        RECT 11.655 188.510 12.015 188.870 ;
        RECT 12.365 188.510 12.725 188.870 ;
        RECT 13.075 188.510 13.435 188.870 ;
        RECT 13.785 188.510 14.145 188.870 ;
        RECT 14.495 188.510 14.855 188.870 ;
        RECT 15.205 188.510 15.565 188.870 ;
        RECT 15.915 188.510 16.275 188.870 ;
        RECT 16.625 188.510 16.985 188.870 ;
        RECT 17.335 188.510 17.695 188.870 ;
        RECT 18.045 188.510 18.405 188.870 ;
        RECT 18.755 188.510 19.115 188.870 ;
        RECT 19.465 188.510 19.825 188.870 ;
        RECT 20.175 188.510 20.535 188.870 ;
        RECT 20.885 188.510 21.245 188.870 ;
        RECT 21.595 188.510 21.955 188.870 ;
        RECT 22.305 188.510 22.665 188.870 ;
        RECT 23.015 188.510 23.375 188.870 ;
        RECT 23.725 188.510 24.085 188.870 ;
        RECT 24.435 188.510 24.795 188.870 ;
        RECT 25.145 188.510 25.505 188.870 ;
        RECT 25.855 188.510 26.215 188.870 ;
        RECT 26.565 188.510 26.925 188.870 ;
        RECT 27.275 188.510 27.635 188.870 ;
        RECT 27.985 188.510 28.345 188.870 ;
        RECT 28.695 188.510 29.055 188.870 ;
        RECT 29.405 188.510 29.765 188.870 ;
        RECT 30.115 188.510 30.475 188.870 ;
        RECT 30.825 188.510 31.185 188.870 ;
        RECT 31.535 188.510 31.895 188.870 ;
        RECT 32.245 188.510 32.605 188.870 ;
        RECT 32.955 188.510 33.315 188.870 ;
        RECT 33.665 188.510 34.025 188.870 ;
        RECT 34.375 188.510 34.735 188.870 ;
        RECT 35.085 188.510 35.445 188.870 ;
      LAYER M5 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V4 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
    END
  END GND
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.700 187.720 ;
        RECT 0.130 177.560 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.885 ;
        RECT 0.130 162.085 0.700 170.040 ;
        RECT 0.130 154.785 0.700 160.610 ;
        RECT 0.130 86.045 0.700 87.905 ;
        RECT 0.130 79.535 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 74.280 ;
        RECT 0.000 0.000 0.345 78.095 ;
        RECT 0.000 77.765 0.700 78.095 ;
        RECT 4.680 0.000 10.595 0.700 ;
        RECT 21.150 0.000 27.070 0.700 ;
        RECT 29.405 0.000 35.325 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.720 ;
        RECT 39.300 177.560 39.870 184.900 ;
        RECT 39.300 171.540 39.870 176.885 ;
        RECT 39.300 162.140 39.870 169.985 ;
        RECT 39.300 154.840 39.870 160.555 ;
        RECT 39.300 86.045 39.870 87.905 ;
        RECT 39.300 79.535 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 74.280 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.700 187.775 ;
        RECT 0.000 177.565 0.700 184.480 ;
        RECT 0.000 171.540 0.700 176.885 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 40.000 187.775 ;
        RECT 39.300 177.565 40.000 184.480 ;
        RECT 39.300 171.540 40.000 176.885 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 85.980 40.000 160.610 ;
        RECT 39.300 79.600 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 74.280 ;
        RECT 0.000 0.000 0.700 76.370 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 39.625 0.000 40.000 78.100 ;
        RECT 39.300 77.770 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.700 187.720 ;
        RECT 0.130 177.560 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.885 ;
        RECT 0.130 162.085 0.700 170.040 ;
        RECT 0.130 154.785 0.700 160.610 ;
        RECT 0.130 86.045 0.700 87.905 ;
        RECT 0.130 79.535 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 74.280 ;
        RECT 0.000 0.000 0.345 78.095 ;
        RECT 0.000 77.765 0.700 78.095 ;
        RECT 4.680 0.000 10.595 0.700 ;
        RECT 21.150 0.000 27.070 0.700 ;
        RECT 29.405 0.000 35.325 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.720 ;
        RECT 39.300 177.560 39.870 184.900 ;
        RECT 39.300 171.540 39.870 176.885 ;
        RECT 39.300 162.140 39.870 169.985 ;
        RECT 39.300 154.840 39.870 160.555 ;
        RECT 39.300 86.045 39.870 87.905 ;
        RECT 39.300 79.535 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 74.335 ;
        RECT 39.625 0.000 40.000 78.155 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.130 185.345 0.700 187.720 ;
        RECT 0.130 177.560 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.885 ;
        RECT 0.130 162.140 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 87.905 ;
        RECT 0.130 79.535 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.720 ;
        RECT 39.300 177.560 39.870 184.955 ;
        RECT 39.300 171.540 39.870 176.885 ;
        RECT 39.300 162.140 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 87.905 ;
        RECT 39.300 79.535 39.870 84.480 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 74.280 ;
        RECT 39.300 0.000 40.000 74.280 ;
        RECT 0.000 0.000 0.345 78.095 ;
        RECT 0.000 77.765 0.700 78.095 ;
        RECT 39.625 0.000 40.000 78.100 ;
  END 
END PSVSSC

MACRO PSVDDO
  CLASS  PAD ;
  FOREIGN PSVDDO 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN VDDO
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
        RECT 4.210 188.300 35.790 189.000 ;
      LAYER V3 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
        RECT 4.210 188.300 35.790 189.000 ;
      LAYER V2 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M2 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V1 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M1 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER M6 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V5 ;
        RECT 4.555 188.510 4.915 188.870 ;
        RECT 5.265 188.510 5.625 188.870 ;
        RECT 5.975 188.510 6.335 188.870 ;
        RECT 6.685 188.510 7.045 188.870 ;
        RECT 7.395 188.510 7.755 188.870 ;
        RECT 8.105 188.510 8.465 188.870 ;
        RECT 8.815 188.510 9.175 188.870 ;
        RECT 9.525 188.510 9.885 188.870 ;
        RECT 10.235 188.510 10.595 188.870 ;
        RECT 10.945 188.510 11.305 188.870 ;
        RECT 11.655 188.510 12.015 188.870 ;
        RECT 12.365 188.510 12.725 188.870 ;
        RECT 13.075 188.510 13.435 188.870 ;
        RECT 13.785 188.510 14.145 188.870 ;
        RECT 14.495 188.510 14.855 188.870 ;
        RECT 15.205 188.510 15.565 188.870 ;
        RECT 15.915 188.510 16.275 188.870 ;
        RECT 16.625 188.510 16.985 188.870 ;
        RECT 17.335 188.510 17.695 188.870 ;
        RECT 18.045 188.510 18.405 188.870 ;
        RECT 18.755 188.510 19.115 188.870 ;
        RECT 19.465 188.510 19.825 188.870 ;
        RECT 20.175 188.510 20.535 188.870 ;
        RECT 20.885 188.510 21.245 188.870 ;
        RECT 21.595 188.510 21.955 188.870 ;
        RECT 22.305 188.510 22.665 188.870 ;
        RECT 23.015 188.510 23.375 188.870 ;
        RECT 23.725 188.510 24.085 188.870 ;
        RECT 24.435 188.510 24.795 188.870 ;
        RECT 25.145 188.510 25.505 188.870 ;
        RECT 25.855 188.510 26.215 188.870 ;
        RECT 26.565 188.510 26.925 188.870 ;
        RECT 27.275 188.510 27.635 188.870 ;
        RECT 27.985 188.510 28.345 188.870 ;
        RECT 28.695 188.510 29.055 188.870 ;
        RECT 29.405 188.510 29.765 188.870 ;
        RECT 30.115 188.510 30.475 188.870 ;
        RECT 30.825 188.510 31.185 188.870 ;
        RECT 31.535 188.510 31.895 188.870 ;
        RECT 32.245 188.510 32.605 188.870 ;
        RECT 32.955 188.510 33.315 188.870 ;
        RECT 33.665 188.510 34.025 188.870 ;
        RECT 34.375 188.510 34.735 188.870 ;
        RECT 35.085 188.510 35.445 188.870 ;
      LAYER M5 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V4 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
    END
  END VDDO
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.700 187.720 ;
        RECT 0.130 177.560 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.885 ;
        RECT 0.130 162.085 0.700 170.040 ;
        RECT 0.130 154.785 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.720 ;
        RECT 39.300 177.560 39.870 184.900 ;
        RECT 39.300 171.540 39.870 176.885 ;
        RECT 39.300 162.140 39.870 169.985 ;
        RECT 39.300 154.840 39.870 160.555 ;
        RECT 39.300 85.080 39.870 87.960 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.700 187.775 ;
        RECT 0.000 177.565 0.700 184.480 ;
        RECT 0.000 171.540 0.700 176.885 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 74.720 39.320 77.020 ;
        RECT 39.300 185.345 40.000 187.775 ;
        RECT 39.300 177.565 40.000 184.480 ;
        RECT 39.300 171.540 40.000 176.885 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 85.980 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 74.280 ;
        RECT 0.000 0.000 0.700 76.470 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.800 0.700 78.100 ;
        RECT 39.625 0.000 40.000 78.100 ;
        RECT 39.300 77.800 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.700 187.720 ;
        RECT 0.130 177.560 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.885 ;
        RECT 0.130 162.085 0.700 170.040 ;
        RECT 0.130 154.785 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.720 ;
        RECT 39.300 177.560 39.870 184.900 ;
        RECT 39.300 171.540 39.870 176.885 ;
        RECT 39.300 162.140 39.870 169.985 ;
        RECT 39.300 154.840 39.870 160.555 ;
        RECT 39.300 85.080 39.870 88.860 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.130 185.345 0.700 187.720 ;
        RECT 0.130 177.560 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.885 ;
        RECT 0.130 162.140 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.100 0.700 87.960 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 74.280 ;
        RECT 0.000 72.380 0.700 74.280 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.720 ;
        RECT 39.300 177.560 39.870 184.955 ;
        RECT 39.300 171.540 39.870 176.885 ;
        RECT 39.300 162.140 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.980 39.870 88.860 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 74.280 ;
        RECT 39.300 72.300 40.000 74.280 ;
        RECT 39.625 0.000 40.000 78.100 ;
  END 
END PSVDDO

MACRO PSVDDC
  CLASS  PAD ;
  FOREIGN PSVDDC 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    CLASS CORE ;
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
        RECT 4.210 188.300 35.790 189.000 ;
      LAYER V3 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
        RECT 4.210 188.300 35.790 189.000 ;
      LAYER V2 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M2 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V1 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M1 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER M6 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V5 ;
        RECT 4.555 188.510 4.915 188.870 ;
        RECT 5.265 188.510 5.625 188.870 ;
        RECT 5.975 188.510 6.335 188.870 ;
        RECT 6.685 188.510 7.045 188.870 ;
        RECT 7.395 188.510 7.755 188.870 ;
        RECT 8.105 188.510 8.465 188.870 ;
        RECT 8.815 188.510 9.175 188.870 ;
        RECT 9.525 188.510 9.885 188.870 ;
        RECT 10.235 188.510 10.595 188.870 ;
        RECT 10.945 188.510 11.305 188.870 ;
        RECT 11.655 188.510 12.015 188.870 ;
        RECT 12.365 188.510 12.725 188.870 ;
        RECT 13.075 188.510 13.435 188.870 ;
        RECT 13.785 188.510 14.145 188.870 ;
        RECT 14.495 188.510 14.855 188.870 ;
        RECT 15.205 188.510 15.565 188.870 ;
        RECT 15.915 188.510 16.275 188.870 ;
        RECT 16.625 188.510 16.985 188.870 ;
        RECT 17.335 188.510 17.695 188.870 ;
        RECT 18.045 188.510 18.405 188.870 ;
        RECT 18.755 188.510 19.115 188.870 ;
        RECT 19.465 188.510 19.825 188.870 ;
        RECT 20.175 188.510 20.535 188.870 ;
        RECT 20.885 188.510 21.245 188.870 ;
        RECT 21.595 188.510 21.955 188.870 ;
        RECT 22.305 188.510 22.665 188.870 ;
        RECT 23.015 188.510 23.375 188.870 ;
        RECT 23.725 188.510 24.085 188.870 ;
        RECT 24.435 188.510 24.795 188.870 ;
        RECT 25.145 188.510 25.505 188.870 ;
        RECT 25.855 188.510 26.215 188.870 ;
        RECT 26.565 188.510 26.925 188.870 ;
        RECT 27.275 188.510 27.635 188.870 ;
        RECT 27.985 188.510 28.345 188.870 ;
        RECT 28.695 188.510 29.055 188.870 ;
        RECT 29.405 188.510 29.765 188.870 ;
        RECT 30.115 188.510 30.475 188.870 ;
        RECT 30.825 188.510 31.185 188.870 ;
        RECT 31.535 188.510 31.895 188.870 ;
        RECT 32.245 188.510 32.605 188.870 ;
        RECT 32.955 188.510 33.315 188.870 ;
        RECT 33.665 188.510 34.025 188.870 ;
        RECT 34.375 188.510 34.735 188.870 ;
        RECT 35.085 188.510 35.445 188.870 ;
      LAYER M5 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V4 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
    END
  END VDD
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.700 187.720 ;
        RECT 0.130 177.560 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.885 ;
        RECT 0.130 162.085 0.700 170.040 ;
        RECT 0.130 154.785 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.720 ;
        RECT 39.300 177.560 39.870 184.900 ;
        RECT 39.300 171.540 39.870 176.885 ;
        RECT 39.300 162.140 39.870 169.985 ;
        RECT 39.300 154.840 39.870 160.555 ;
        RECT 39.300 85.080 39.870 87.960 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.700 187.775 ;
        RECT 0.000 177.565 0.700 184.480 ;
        RECT 0.000 171.540 0.700 176.885 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 74.720 39.320 77.020 ;
        RECT 39.300 185.345 40.000 187.775 ;
        RECT 39.300 177.565 40.000 184.480 ;
        RECT 39.300 171.540 40.000 176.885 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 85.980 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 74.280 ;
        RECT 0.000 0.000 0.700 76.470 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.800 0.700 78.100 ;
        RECT 39.625 0.000 40.000 78.100 ;
        RECT 39.300 77.800 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.700 187.720 ;
        RECT 0.130 177.560 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.885 ;
        RECT 0.130 162.085 0.700 170.040 ;
        RECT 0.130 154.785 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.720 ;
        RECT 39.300 177.560 39.870 184.900 ;
        RECT 39.300 171.540 39.870 176.885 ;
        RECT 39.300 162.140 39.870 169.985 ;
        RECT 39.300 154.840 39.870 160.555 ;
        RECT 39.300 85.080 39.870 88.860 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.130 185.345 0.700 187.720 ;
        RECT 0.130 177.560 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.885 ;
        RECT 0.130 162.140 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.100 0.700 87.960 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 74.280 ;
        RECT 0.000 72.380 0.700 74.280 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.720 ;
        RECT 39.300 177.560 39.870 184.955 ;
        RECT 39.300 171.540 39.870 176.885 ;
        RECT 39.300 162.140 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.980 39.870 88.860 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 74.280 ;
        RECT 39.300 72.300 40.000 74.280 ;
        RECT 39.625 0.000 40.000 78.100 ;
  END 
END PSVDDC

MACRO PSVDDH
  CLASS  PAD ;
  FOREIGN PSVDDH 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN VDDH
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
        RECT 4.210 188.300 35.790 189.000 ;
      LAYER V3 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
        RECT 4.210 188.300 35.790 189.000 ;
      LAYER V2 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M2 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V1 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M1 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER M6 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V5 ;
        RECT 4.555 188.510 4.915 188.870 ;
        RECT 5.265 188.510 5.625 188.870 ;
        RECT 5.975 188.510 6.335 188.870 ;
        RECT 6.685 188.510 7.045 188.870 ;
        RECT 7.395 188.510 7.755 188.870 ;
        RECT 8.105 188.510 8.465 188.870 ;
        RECT 8.815 188.510 9.175 188.870 ;
        RECT 9.525 188.510 9.885 188.870 ;
        RECT 10.235 188.510 10.595 188.870 ;
        RECT 10.945 188.510 11.305 188.870 ;
        RECT 11.655 188.510 12.015 188.870 ;
        RECT 12.365 188.510 12.725 188.870 ;
        RECT 13.075 188.510 13.435 188.870 ;
        RECT 13.785 188.510 14.145 188.870 ;
        RECT 14.495 188.510 14.855 188.870 ;
        RECT 15.205 188.510 15.565 188.870 ;
        RECT 15.915 188.510 16.275 188.870 ;
        RECT 16.625 188.510 16.985 188.870 ;
        RECT 17.335 188.510 17.695 188.870 ;
        RECT 18.045 188.510 18.405 188.870 ;
        RECT 18.755 188.510 19.115 188.870 ;
        RECT 19.465 188.510 19.825 188.870 ;
        RECT 20.175 188.510 20.535 188.870 ;
        RECT 20.885 188.510 21.245 188.870 ;
        RECT 21.595 188.510 21.955 188.870 ;
        RECT 22.305 188.510 22.665 188.870 ;
        RECT 23.015 188.510 23.375 188.870 ;
        RECT 23.725 188.510 24.085 188.870 ;
        RECT 24.435 188.510 24.795 188.870 ;
        RECT 25.145 188.510 25.505 188.870 ;
        RECT 25.855 188.510 26.215 188.870 ;
        RECT 26.565 188.510 26.925 188.870 ;
        RECT 27.275 188.510 27.635 188.870 ;
        RECT 27.985 188.510 28.345 188.870 ;
        RECT 28.695 188.510 29.055 188.870 ;
        RECT 29.405 188.510 29.765 188.870 ;
        RECT 30.115 188.510 30.475 188.870 ;
        RECT 30.825 188.510 31.185 188.870 ;
        RECT 31.535 188.510 31.895 188.870 ;
        RECT 32.245 188.510 32.605 188.870 ;
        RECT 32.955 188.510 33.315 188.870 ;
        RECT 33.665 188.510 34.025 188.870 ;
        RECT 34.375 188.510 34.735 188.870 ;
        RECT 35.085 188.510 35.445 188.870 ;
      LAYER M5 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V4 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
    END
  END VDDH
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.700 187.720 ;
        RECT 0.130 177.560 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.885 ;
        RECT 0.130 162.085 0.700 170.040 ;
        RECT 0.130 154.785 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.720 ;
        RECT 39.300 177.560 39.870 184.900 ;
        RECT 39.300 171.540 39.870 176.885 ;
        RECT 39.300 162.140 39.870 169.985 ;
        RECT 39.300 154.840 39.870 160.555 ;
        RECT 39.300 85.080 39.870 87.960 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.700 187.775 ;
        RECT 0.000 177.565 0.700 184.480 ;
        RECT 0.000 171.540 0.700 176.885 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 74.720 39.320 77.020 ;
        RECT 39.300 185.345 40.000 187.775 ;
        RECT 39.300 177.565 40.000 184.480 ;
        RECT 39.300 171.540 40.000 176.885 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 85.980 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 74.280 ;
        RECT 0.000 0.000 0.700 76.470 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.800 0.700 78.100 ;
        RECT 39.625 0.000 40.000 78.100 ;
        RECT 39.300 77.800 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.700 187.720 ;
        RECT 0.130 177.560 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.885 ;
        RECT 0.130 162.085 0.700 170.040 ;
        RECT 0.130 154.785 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.720 ;
        RECT 39.300 177.560 39.870 184.900 ;
        RECT 39.300 171.540 39.870 176.885 ;
        RECT 39.300 162.140 39.870 169.985 ;
        RECT 39.300 154.840 39.870 160.555 ;
        RECT 39.300 85.080 39.870 88.860 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.130 185.345 0.700 187.720 ;
        RECT 0.130 177.560 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.885 ;
        RECT 0.130 162.140 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.100 0.700 87.960 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 74.280 ;
        RECT 0.000 72.380 0.700 74.280 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.720 ;
        RECT 39.300 177.560 39.870 184.955 ;
        RECT 39.300 171.540 39.870 176.885 ;
        RECT 39.300 162.140 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.980 39.870 88.860 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 74.280 ;
        RECT 39.300 72.300 40.000 74.280 ;
        RECT 39.625 0.000 40.000 78.100 ;
  END 
END PSVDDH

MACRO PSOSCR14M
  CLASS  PAD ;
  FOREIGN PSOSCR14M 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 115.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN XTALIN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 47.530 0.000 53.450 0.700 ;
      LAYER M3 ;
        RECT 47.530 0.000 53.450 0.700 ;
    END
  END XTALIN
  PIN EI
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 16.680 188.380 17.680 189.000 ;
      LAYER V3 ;
        RECT 16.880 188.800 17.070 188.990 ;
        RECT 16.880 188.390 17.070 188.580 ;
        RECT 17.290 188.800 17.480 188.990 ;
        RECT 17.290 188.390 17.480 188.580 ;
      LAYER M3 ;
        RECT 16.680 188.380 17.680 189.000 ;
      LAYER V2 ;
        RECT 16.880 188.800 17.070 188.990 ;
        RECT 16.880 188.390 17.070 188.580 ;
        RECT 17.290 188.800 17.480 188.990 ;
        RECT 17.290 188.390 17.480 188.580 ;
      LAYER M2 ;
        RECT 17.075 188.300 17.285 189.000 ;
        RECT 16.680 188.380 17.680 189.000 ;
      LAYER V1 ;
        RECT 16.880 188.800 17.070 188.990 ;
        RECT 16.880 188.390 17.070 188.580 ;
        RECT 17.290 188.800 17.480 188.990 ;
        RECT 17.290 188.390 17.480 188.580 ;
      LAYER M1 ;
        RECT 16.680 188.380 17.680 189.000 ;
      LAYER M6 ;
        RECT 16.680 188.380 17.680 189.000 ;
      LAYER V5 ;
        RECT 17.000 188.510 17.360 188.870 ;
      LAYER M5 ;
        RECT 16.680 188.380 17.680 189.000 ;
      LAYER V4 ;
        RECT 16.880 188.800 17.070 188.990 ;
        RECT 16.880 188.390 17.070 188.580 ;
        RECT 17.290 188.800 17.480 188.990 ;
        RECT 17.290 188.390 17.480 188.580 ;
    END
  END EI
  PIN XTALOUT
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 96.550 0.000 102.470 0.700 ;
      LAYER M3 ;
        RECT 96.550 0.000 102.470 0.700 ;
    END
  END XTALOUT
  PIN EO
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 97.085 188.380 98.085 189.000 ;
      LAYER V3 ;
        RECT 97.285 188.800 97.475 188.990 ;
        RECT 97.285 188.390 97.475 188.580 ;
        RECT 97.695 188.800 97.885 188.990 ;
        RECT 97.695 188.390 97.885 188.580 ;
      LAYER M3 ;
        RECT 97.085 188.380 98.085 189.000 ;
      LAYER V2 ;
        RECT 97.285 188.800 97.475 188.990 ;
        RECT 97.285 188.390 97.475 188.580 ;
        RECT 97.695 188.800 97.885 188.990 ;
        RECT 97.695 188.390 97.885 188.580 ;
      LAYER M2 ;
        RECT 97.480 188.300 97.690 189.000 ;
        RECT 97.085 188.380 98.085 189.000 ;
      LAYER V1 ;
        RECT 97.285 188.800 97.475 188.990 ;
        RECT 97.285 188.390 97.475 188.580 ;
        RECT 97.695 188.800 97.885 188.990 ;
        RECT 97.695 188.390 97.885 188.580 ;
      LAYER M1 ;
        RECT 97.085 188.380 98.085 189.000 ;
      LAYER M6 ;
        RECT 97.085 188.380 98.085 189.000 ;
      LAYER V5 ;
        RECT 97.405 188.510 97.765 188.870 ;
      LAYER M5 ;
        RECT 97.085 188.380 98.085 189.000 ;
      LAYER V4 ;
        RECT 97.285 188.800 97.475 188.990 ;
        RECT 97.285 188.390 97.475 188.580 ;
        RECT 97.695 188.800 97.885 188.990 ;
        RECT 97.695 188.390 97.885 188.580 ;
    END
  END EO
  PIN CK
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 56.005 188.380 64.005 189.000 ;
      LAYER V3 ;
        RECT 56.220 188.800 56.410 188.990 ;
        RECT 56.220 188.390 56.410 188.580 ;
        RECT 56.630 188.800 56.820 188.990 ;
        RECT 56.630 188.390 56.820 188.580 ;
        RECT 57.040 188.800 57.230 188.990 ;
        RECT 57.040 188.390 57.230 188.580 ;
        RECT 57.450 188.800 57.640 188.990 ;
        RECT 57.450 188.390 57.640 188.580 ;
        RECT 57.860 188.800 58.050 188.990 ;
        RECT 57.860 188.390 58.050 188.580 ;
        RECT 58.270 188.800 58.460 188.990 ;
        RECT 58.270 188.390 58.460 188.580 ;
        RECT 58.680 188.800 58.870 188.990 ;
        RECT 58.680 188.390 58.870 188.580 ;
        RECT 59.090 188.800 59.280 188.990 ;
        RECT 59.090 188.390 59.280 188.580 ;
        RECT 59.500 188.800 59.690 188.990 ;
        RECT 59.500 188.390 59.690 188.580 ;
        RECT 59.910 188.800 60.100 188.990 ;
        RECT 59.910 188.390 60.100 188.580 ;
        RECT 60.320 188.800 60.510 188.990 ;
        RECT 60.320 188.390 60.510 188.580 ;
        RECT 60.730 188.800 60.920 188.990 ;
        RECT 60.730 188.390 60.920 188.580 ;
        RECT 61.140 188.800 61.330 188.990 ;
        RECT 61.140 188.390 61.330 188.580 ;
        RECT 61.550 188.800 61.740 188.990 ;
        RECT 61.550 188.390 61.740 188.580 ;
        RECT 61.960 188.800 62.150 188.990 ;
        RECT 61.960 188.390 62.150 188.580 ;
        RECT 62.370 188.800 62.560 188.990 ;
        RECT 62.370 188.390 62.560 188.580 ;
        RECT 62.780 188.800 62.970 188.990 ;
        RECT 62.780 188.390 62.970 188.580 ;
        RECT 63.190 188.800 63.380 188.990 ;
        RECT 63.190 188.390 63.380 188.580 ;
        RECT 63.600 188.800 63.790 188.990 ;
        RECT 63.600 188.390 63.790 188.580 ;
      LAYER M3 ;
        RECT 56.005 188.380 64.005 189.000 ;
      LAYER V2 ;
        RECT 56.220 188.800 56.410 188.990 ;
        RECT 56.220 188.390 56.410 188.580 ;
        RECT 56.630 188.800 56.820 188.990 ;
        RECT 56.630 188.390 56.820 188.580 ;
        RECT 57.040 188.800 57.230 188.990 ;
        RECT 57.040 188.390 57.230 188.580 ;
        RECT 57.450 188.800 57.640 188.990 ;
        RECT 57.450 188.390 57.640 188.580 ;
        RECT 57.860 188.800 58.050 188.990 ;
        RECT 57.860 188.390 58.050 188.580 ;
        RECT 58.270 188.800 58.460 188.990 ;
        RECT 58.270 188.390 58.460 188.580 ;
        RECT 58.680 188.800 58.870 188.990 ;
        RECT 58.680 188.390 58.870 188.580 ;
        RECT 59.090 188.800 59.280 188.990 ;
        RECT 59.090 188.390 59.280 188.580 ;
        RECT 59.500 188.800 59.690 188.990 ;
        RECT 59.500 188.390 59.690 188.580 ;
        RECT 59.910 188.800 60.100 188.990 ;
        RECT 59.910 188.390 60.100 188.580 ;
        RECT 60.320 188.800 60.510 188.990 ;
        RECT 60.320 188.390 60.510 188.580 ;
        RECT 60.730 188.800 60.920 188.990 ;
        RECT 60.730 188.390 60.920 188.580 ;
        RECT 61.140 188.800 61.330 188.990 ;
        RECT 61.140 188.390 61.330 188.580 ;
        RECT 61.550 188.800 61.740 188.990 ;
        RECT 61.550 188.390 61.740 188.580 ;
        RECT 61.960 188.800 62.150 188.990 ;
        RECT 61.960 188.390 62.150 188.580 ;
        RECT 62.370 188.800 62.560 188.990 ;
        RECT 62.370 188.390 62.560 188.580 ;
        RECT 62.780 188.800 62.970 188.990 ;
        RECT 62.780 188.390 62.970 188.580 ;
        RECT 63.190 188.800 63.380 188.990 ;
        RECT 63.190 188.390 63.380 188.580 ;
        RECT 63.600 188.800 63.790 188.990 ;
        RECT 63.600 188.390 63.790 188.580 ;
      LAYER M2 ;
        RECT 56.005 188.300 64.005 189.000 ;
      LAYER V1 ;
        RECT 56.220 188.800 56.410 188.990 ;
        RECT 56.220 188.390 56.410 188.580 ;
        RECT 56.630 188.800 56.820 188.990 ;
        RECT 56.630 188.390 56.820 188.580 ;
        RECT 57.040 188.800 57.230 188.990 ;
        RECT 57.040 188.390 57.230 188.580 ;
        RECT 57.450 188.800 57.640 188.990 ;
        RECT 57.450 188.390 57.640 188.580 ;
        RECT 57.860 188.800 58.050 188.990 ;
        RECT 57.860 188.390 58.050 188.580 ;
        RECT 58.270 188.800 58.460 188.990 ;
        RECT 58.270 188.390 58.460 188.580 ;
        RECT 58.680 188.800 58.870 188.990 ;
        RECT 58.680 188.390 58.870 188.580 ;
        RECT 59.090 188.800 59.280 188.990 ;
        RECT 59.090 188.390 59.280 188.580 ;
        RECT 59.500 188.800 59.690 188.990 ;
        RECT 59.500 188.390 59.690 188.580 ;
        RECT 59.910 188.800 60.100 188.990 ;
        RECT 59.910 188.390 60.100 188.580 ;
        RECT 60.320 188.800 60.510 188.990 ;
        RECT 60.320 188.390 60.510 188.580 ;
        RECT 60.730 188.800 60.920 188.990 ;
        RECT 60.730 188.390 60.920 188.580 ;
        RECT 61.140 188.800 61.330 188.990 ;
        RECT 61.140 188.390 61.330 188.580 ;
        RECT 61.550 188.800 61.740 188.990 ;
        RECT 61.550 188.390 61.740 188.580 ;
        RECT 61.960 188.800 62.150 188.990 ;
        RECT 61.960 188.390 62.150 188.580 ;
        RECT 62.370 188.800 62.560 188.990 ;
        RECT 62.370 188.390 62.560 188.580 ;
        RECT 62.780 188.800 62.970 188.990 ;
        RECT 62.780 188.390 62.970 188.580 ;
        RECT 63.190 188.800 63.380 188.990 ;
        RECT 63.190 188.390 63.380 188.580 ;
        RECT 63.600 188.800 63.790 188.990 ;
        RECT 63.600 188.390 63.790 188.580 ;
      LAYER M1 ;
        RECT 56.005 188.380 64.005 189.000 ;
      LAYER M6 ;
        RECT 56.005 188.380 64.005 189.000 ;
      LAYER V5 ;
        RECT 56.275 188.510 56.635 188.870 ;
        RECT 56.985 188.510 57.345 188.870 ;
        RECT 57.695 188.510 58.055 188.870 ;
        RECT 58.405 188.510 58.765 188.870 ;
        RECT 59.115 188.510 59.475 188.870 ;
        RECT 59.825 188.510 60.185 188.870 ;
        RECT 60.535 188.510 60.895 188.870 ;
        RECT 61.245 188.510 61.605 188.870 ;
        RECT 61.955 188.510 62.315 188.870 ;
        RECT 62.665 188.510 63.025 188.870 ;
        RECT 63.375 188.510 63.735 188.870 ;
      LAYER M5 ;
        RECT 56.005 188.380 64.005 189.000 ;
      LAYER V4 ;
        RECT 56.220 188.800 56.410 188.990 ;
        RECT 56.220 188.390 56.410 188.580 ;
        RECT 56.630 188.800 56.820 188.990 ;
        RECT 56.630 188.390 56.820 188.580 ;
        RECT 57.040 188.800 57.230 188.990 ;
        RECT 57.040 188.390 57.230 188.580 ;
        RECT 57.450 188.800 57.640 188.990 ;
        RECT 57.450 188.390 57.640 188.580 ;
        RECT 57.860 188.800 58.050 188.990 ;
        RECT 57.860 188.390 58.050 188.580 ;
        RECT 58.270 188.800 58.460 188.990 ;
        RECT 58.270 188.390 58.460 188.580 ;
        RECT 58.680 188.800 58.870 188.990 ;
        RECT 58.680 188.390 58.870 188.580 ;
        RECT 59.090 188.800 59.280 188.990 ;
        RECT 59.090 188.390 59.280 188.580 ;
        RECT 59.500 188.800 59.690 188.990 ;
        RECT 59.500 188.390 59.690 188.580 ;
        RECT 59.910 188.800 60.100 188.990 ;
        RECT 59.910 188.390 60.100 188.580 ;
        RECT 60.320 188.800 60.510 188.990 ;
        RECT 60.320 188.390 60.510 188.580 ;
        RECT 60.730 188.800 60.920 188.990 ;
        RECT 60.730 188.390 60.920 188.580 ;
        RECT 61.140 188.800 61.330 188.990 ;
        RECT 61.140 188.390 61.330 188.580 ;
        RECT 61.550 188.800 61.740 188.990 ;
        RECT 61.550 188.390 61.740 188.580 ;
        RECT 61.960 188.800 62.150 188.990 ;
        RECT 61.960 188.390 62.150 188.580 ;
        RECT 62.370 188.800 62.560 188.990 ;
        RECT 62.370 188.390 62.560 188.580 ;
        RECT 62.780 188.800 62.970 188.990 ;
        RECT 62.780 188.390 62.970 188.580 ;
        RECT 63.190 188.800 63.380 188.990 ;
        RECT 63.190 188.390 63.380 188.580 ;
        RECT 63.600 188.800 63.790 188.990 ;
        RECT 63.600 188.390 63.790 188.580 ;
    END
  END CK
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.700 187.775 ;
        RECT 0.130 177.610 0.700 184.950 ;
        RECT 0.130 171.540 0.700 176.940 ;
        RECT 0.130 162.140 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 35.000 0.000 36.500 0.700 ;
        RECT 38.510 0.000 44.430 0.700 ;
        RECT 56.550 0.000 62.470 0.700 ;
        RECT 65.570 0.000 71.490 0.700 ;
        RECT 73.500 0.000 76.500 0.700 ;
        RECT 78.510 0.000 84.430 0.700 ;
        RECT 87.530 0.000 93.450 0.700 ;
        RECT 105.570 0.000 111.490 0.700 ;
        RECT 1.100 1.100 113.900 187.900 ;
        RECT 114.300 185.345 114.870 187.775 ;
        RECT 114.300 177.615 114.870 184.950 ;
        RECT 114.300 171.540 114.870 176.940 ;
        RECT 114.300 162.140 114.870 170.040 ;
        RECT 114.300 155.265 114.870 160.610 ;
        RECT 114.300 86.205 114.870 87.960 ;
        RECT 114.665 79.590 114.870 84.480 ;
        RECT 114.300 83.585 114.870 84.480 ;
        RECT 113.500 0.000 115.000 0.700 ;
        RECT 114.300 0.000 115.000 1.820 ;
        RECT 114.500 0.000 115.000 78.100 ;
        RECT 114.300 72.380 115.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.700 187.775 ;
        RECT 0.000 171.540 0.700 177.145 ;
        RECT 0.000 171.540 0.330 184.975 ;
        RECT 0.000 177.580 0.700 184.975 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.600 0.700 160.610 ;
        RECT 1.100 1.100 113.900 187.900 ;
        RECT 114.300 185.345 115.000 187.775 ;
        RECT 114.300 171.540 115.000 176.980 ;
        RECT 114.670 171.540 115.000 184.975 ;
        RECT 114.300 177.580 115.000 184.975 ;
        RECT 114.300 162.140 115.000 170.040 ;
        RECT 114.300 85.980 115.000 160.610 ;
        RECT 114.665 79.590 115.000 84.480 ;
        RECT 114.300 83.590 115.000 84.480 ;
        RECT 35.000 0.000 115.000 0.400 ;
        RECT 35.000 0.000 36.500 0.700 ;
        RECT 73.500 0.000 76.500 0.700 ;
        RECT 113.500 0.000 115.000 0.700 ;
        RECT 114.300 0.000 115.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.700 187.775 ;
        RECT 0.130 177.610 0.700 185.015 ;
        RECT 0.130 171.540 0.700 176.940 ;
        RECT 0.130 162.140 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 35.000 0.000 36.500 0.700 ;
        RECT 38.510 0.000 44.430 0.700 ;
        RECT 56.550 0.000 62.470 0.700 ;
        RECT 65.570 0.000 71.490 0.700 ;
        RECT 73.500 0.000 76.500 0.700 ;
        RECT 78.510 0.000 84.430 0.700 ;
        RECT 87.530 0.000 93.450 0.700 ;
        RECT 105.570 0.000 111.490 0.700 ;
        RECT 1.100 1.100 113.900 187.900 ;
        RECT 114.300 185.345 114.870 187.775 ;
        RECT 114.300 177.615 114.870 184.950 ;
        RECT 114.300 171.540 114.870 176.940 ;
        RECT 114.300 162.140 114.870 170.040 ;
        RECT 114.300 155.265 114.870 160.610 ;
        RECT 114.300 86.205 114.870 87.960 ;
        RECT 114.665 79.590 114.870 84.480 ;
        RECT 114.300 83.585 114.870 84.480 ;
        RECT 113.500 0.000 115.000 0.700 ;
        RECT 114.300 0.000 115.000 1.820 ;
        RECT 114.500 0.000 115.000 78.100 ;
        RECT 114.300 72.380 115.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 113.900 187.900 ;
        RECT 114.300 185.015 115.000 187.775 ;
        RECT 114.300 177.615 115.000 184.415 ;
        RECT 114.300 170.640 115.000 176.940 ;
        RECT 114.300 162.140 115.000 170.040 ;
        RECT 114.300 154.840 115.000 161.540 ;
        RECT 114.300 139.530 115.000 150.030 ;
        RECT 114.300 127.890 115.000 136.030 ;
        RECT 114.300 116.930 115.000 124.390 ;
        RECT 114.300 105.930 115.000 113.930 ;
        RECT 114.300 94.290 115.000 102.430 ;
        RECT 114.300 90.340 115.000 92.340 ;
        RECT 114.300 85.080 115.000 87.960 ;
        RECT 114.300 79.590 115.000 84.480 ;
        RECT 114.300 71.440 115.000 79.110 ;
        RECT 114.300 57.770 115.000 68.270 ;
        RECT 114.300 45.630 115.000 54.270 ;
        RECT 114.300 32.770 115.000 42.130 ;
        RECT 114.300 20.470 115.000 28.910 ;
        RECT 114.300 9.130 115.000 16.970 ;
        RECT 114.300 3.610 115.000 5.630 ;
        RECT 0.000 0.000 115.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 114.300 0.000 115.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 113.900 187.900 ;
        RECT 114.300 185.400 115.000 187.775 ;
        RECT 114.300 177.615 115.000 184.955 ;
        RECT 114.300 170.640 115.000 176.940 ;
        RECT 114.300 162.140 115.000 170.040 ;
        RECT 114.300 154.840 115.000 161.540 ;
        RECT 114.300 145.030 115.000 150.030 ;
        RECT 114.300 133.390 115.000 141.530 ;
        RECT 114.300 122.170 115.000 129.890 ;
        RECT 114.300 111.430 115.000 119.170 ;
        RECT 114.300 99.790 115.000 107.930 ;
        RECT 114.300 90.340 115.000 96.290 ;
        RECT 114.300 85.080 115.000 87.960 ;
        RECT 114.300 79.590 115.000 84.480 ;
        RECT 114.300 71.440 115.000 79.110 ;
        RECT 114.300 63.270 115.000 68.270 ;
        RECT 114.300 51.630 115.000 59.770 ;
        RECT 114.300 39.130 115.000 48.130 ;
        RECT 114.300 26.270 115.000 35.270 ;
        RECT 114.300 14.630 115.000 22.770 ;
        RECT 114.300 3.610 115.000 11.130 ;
        RECT 0.000 0.000 115.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 114.300 0.000 115.000 2.960 ;
      LAYER M2 ;
        RECT 0.130 185.345 0.700 187.775 ;
        RECT 0.130 177.610 0.700 184.950 ;
        RECT 0.130 171.540 0.700 176.940 ;
        RECT 0.130 162.140 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 35.000 0.000 36.500 0.700 ;
        RECT 73.500 0.000 76.500 0.700 ;
        RECT 1.100 1.100 113.900 187.900 ;
        RECT 114.300 185.345 114.870 187.775 ;
        RECT 114.300 177.615 114.870 184.950 ;
        RECT 114.300 171.540 114.870 176.940 ;
        RECT 114.300 162.140 114.870 170.040 ;
        RECT 114.300 155.265 114.870 160.610 ;
        RECT 114.300 86.205 114.870 87.960 ;
        RECT 114.665 79.590 114.870 84.480 ;
        RECT 114.300 83.585 114.870 84.480 ;
        RECT 113.500 0.000 115.000 0.700 ;
        RECT 114.300 0.000 115.000 1.820 ;
        RECT 114.500 0.000 115.000 78.100 ;
        RECT 114.300 72.380 115.000 78.100 ;
  END 
END PSOSCR14M

MACRO PSOSC14M
  CLASS  PAD ;
  FOREIGN PSOSC14M 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN XTALIN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
    END
  END XTALIN
  PIN EI
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 8.130 188.380 9.130 189.000 ;
      LAYER V3 ;
        RECT 8.330 188.800 8.520 188.990 ;
        RECT 8.330 188.390 8.520 188.580 ;
        RECT 8.740 188.800 8.930 188.990 ;
        RECT 8.740 188.390 8.930 188.580 ;
      LAYER M3 ;
        RECT 8.130 188.380 9.130 189.000 ;
      LAYER V2 ;
        RECT 8.330 188.800 8.520 188.990 ;
        RECT 8.330 188.390 8.520 188.580 ;
        RECT 8.740 188.800 8.930 188.990 ;
        RECT 8.740 188.390 8.930 188.580 ;
      LAYER M2 ;
        RECT 8.525 188.300 8.735 189.000 ;
        RECT 8.130 188.380 9.130 189.000 ;
      LAYER V1 ;
        RECT 8.330 188.800 8.520 188.990 ;
        RECT 8.330 188.390 8.520 188.580 ;
        RECT 8.740 188.800 8.930 188.990 ;
        RECT 8.740 188.390 8.930 188.580 ;
      LAYER M1 ;
        RECT 8.130 188.380 9.130 189.000 ;
      LAYER M6 ;
        RECT 8.130 188.380 9.130 189.000 ;
      LAYER V5 ;
        RECT 8.450 188.510 8.810 188.870 ;
      LAYER M5 ;
        RECT 8.130 188.380 9.130 189.000 ;
      LAYER V4 ;
        RECT 8.330 188.800 8.520 188.990 ;
        RECT 8.330 188.390 8.520 188.580 ;
        RECT 8.740 188.800 8.930 188.990 ;
        RECT 8.740 188.390 8.930 188.580 ;
    END
  END EI
  PIN XTALOUT
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 61.550 0.000 67.470 0.700 ;
      LAYER M3 ;
        RECT 61.550 0.000 67.470 0.700 ;
    END
  END XTALOUT
  PIN EO
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 70.970 188.380 71.970 189.000 ;
      LAYER V3 ;
        RECT 71.170 188.800 71.360 188.990 ;
        RECT 71.170 188.390 71.360 188.580 ;
        RECT 71.580 188.800 71.770 188.990 ;
        RECT 71.580 188.390 71.770 188.580 ;
      LAYER M3 ;
        RECT 70.970 188.380 71.970 189.000 ;
      LAYER V2 ;
        RECT 71.170 188.800 71.360 188.990 ;
        RECT 71.170 188.390 71.360 188.580 ;
        RECT 71.580 188.800 71.770 188.990 ;
        RECT 71.580 188.390 71.770 188.580 ;
      LAYER M2 ;
        RECT 71.365 188.300 71.575 189.000 ;
        RECT 70.970 188.380 71.970 189.000 ;
      LAYER V1 ;
        RECT 71.170 188.800 71.360 188.990 ;
        RECT 71.170 188.390 71.360 188.580 ;
        RECT 71.580 188.800 71.770 188.990 ;
        RECT 71.580 188.390 71.770 188.580 ;
      LAYER M1 ;
        RECT 70.970 188.380 71.970 189.000 ;
      LAYER M6 ;
        RECT 70.970 188.380 71.970 189.000 ;
      LAYER V5 ;
        RECT 71.290 188.510 71.650 188.870 ;
      LAYER M5 ;
        RECT 70.970 188.380 71.970 189.000 ;
      LAYER V4 ;
        RECT 71.170 188.800 71.360 188.990 ;
        RECT 71.170 188.390 71.360 188.580 ;
        RECT 71.580 188.800 71.770 188.990 ;
        RECT 71.580 188.390 71.770 188.580 ;
    END
  END EO
  PIN CK
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 37.400 188.380 45.400 189.000 ;
      LAYER V3 ;
        RECT 37.615 188.800 37.805 188.990 ;
        RECT 37.615 188.390 37.805 188.580 ;
        RECT 38.025 188.800 38.215 188.990 ;
        RECT 38.025 188.390 38.215 188.580 ;
        RECT 38.435 188.800 38.625 188.990 ;
        RECT 38.435 188.390 38.625 188.580 ;
        RECT 38.845 188.800 39.035 188.990 ;
        RECT 38.845 188.390 39.035 188.580 ;
        RECT 39.255 188.800 39.445 188.990 ;
        RECT 39.255 188.390 39.445 188.580 ;
        RECT 39.665 188.800 39.855 188.990 ;
        RECT 39.665 188.390 39.855 188.580 ;
        RECT 40.075 188.800 40.265 188.990 ;
        RECT 40.075 188.390 40.265 188.580 ;
        RECT 40.485 188.800 40.675 188.990 ;
        RECT 40.485 188.390 40.675 188.580 ;
        RECT 40.895 188.800 41.085 188.990 ;
        RECT 40.895 188.390 41.085 188.580 ;
        RECT 41.305 188.800 41.495 188.990 ;
        RECT 41.305 188.390 41.495 188.580 ;
        RECT 41.715 188.800 41.905 188.990 ;
        RECT 41.715 188.390 41.905 188.580 ;
        RECT 42.125 188.800 42.315 188.990 ;
        RECT 42.125 188.390 42.315 188.580 ;
        RECT 42.535 188.800 42.725 188.990 ;
        RECT 42.535 188.390 42.725 188.580 ;
        RECT 42.945 188.800 43.135 188.990 ;
        RECT 42.945 188.390 43.135 188.580 ;
        RECT 43.355 188.800 43.545 188.990 ;
        RECT 43.355 188.390 43.545 188.580 ;
        RECT 43.765 188.800 43.955 188.990 ;
        RECT 43.765 188.390 43.955 188.580 ;
        RECT 44.175 188.800 44.365 188.990 ;
        RECT 44.175 188.390 44.365 188.580 ;
        RECT 44.585 188.800 44.775 188.990 ;
        RECT 44.585 188.390 44.775 188.580 ;
        RECT 44.995 188.800 45.185 188.990 ;
        RECT 44.995 188.390 45.185 188.580 ;
      LAYER M3 ;
        RECT 37.400 188.380 45.400 189.000 ;
      LAYER V2 ;
        RECT 37.615 188.800 37.805 188.990 ;
        RECT 37.615 188.390 37.805 188.580 ;
        RECT 38.025 188.800 38.215 188.990 ;
        RECT 38.025 188.390 38.215 188.580 ;
        RECT 38.435 188.800 38.625 188.990 ;
        RECT 38.435 188.390 38.625 188.580 ;
        RECT 38.845 188.800 39.035 188.990 ;
        RECT 38.845 188.390 39.035 188.580 ;
        RECT 39.255 188.800 39.445 188.990 ;
        RECT 39.255 188.390 39.445 188.580 ;
        RECT 39.665 188.800 39.855 188.990 ;
        RECT 39.665 188.390 39.855 188.580 ;
        RECT 40.075 188.800 40.265 188.990 ;
        RECT 40.075 188.390 40.265 188.580 ;
        RECT 40.485 188.800 40.675 188.990 ;
        RECT 40.485 188.390 40.675 188.580 ;
        RECT 40.895 188.800 41.085 188.990 ;
        RECT 40.895 188.390 41.085 188.580 ;
        RECT 41.305 188.800 41.495 188.990 ;
        RECT 41.305 188.390 41.495 188.580 ;
        RECT 41.715 188.800 41.905 188.990 ;
        RECT 41.715 188.390 41.905 188.580 ;
        RECT 42.125 188.800 42.315 188.990 ;
        RECT 42.125 188.390 42.315 188.580 ;
        RECT 42.535 188.800 42.725 188.990 ;
        RECT 42.535 188.390 42.725 188.580 ;
        RECT 42.945 188.800 43.135 188.990 ;
        RECT 42.945 188.390 43.135 188.580 ;
        RECT 43.355 188.800 43.545 188.990 ;
        RECT 43.355 188.390 43.545 188.580 ;
        RECT 43.765 188.800 43.955 188.990 ;
        RECT 43.765 188.390 43.955 188.580 ;
        RECT 44.175 188.800 44.365 188.990 ;
        RECT 44.175 188.390 44.365 188.580 ;
        RECT 44.585 188.800 44.775 188.990 ;
        RECT 44.585 188.390 44.775 188.580 ;
        RECT 44.995 188.800 45.185 188.990 ;
        RECT 44.995 188.390 45.185 188.580 ;
      LAYER M2 ;
        RECT 37.400 188.300 45.400 189.000 ;
      LAYER V1 ;
        RECT 37.615 188.800 37.805 188.990 ;
        RECT 37.615 188.390 37.805 188.580 ;
        RECT 38.025 188.800 38.215 188.990 ;
        RECT 38.025 188.390 38.215 188.580 ;
        RECT 38.435 188.800 38.625 188.990 ;
        RECT 38.435 188.390 38.625 188.580 ;
        RECT 38.845 188.800 39.035 188.990 ;
        RECT 38.845 188.390 39.035 188.580 ;
        RECT 39.255 188.800 39.445 188.990 ;
        RECT 39.255 188.390 39.445 188.580 ;
        RECT 39.665 188.800 39.855 188.990 ;
        RECT 39.665 188.390 39.855 188.580 ;
        RECT 40.075 188.800 40.265 188.990 ;
        RECT 40.075 188.390 40.265 188.580 ;
        RECT 40.485 188.800 40.675 188.990 ;
        RECT 40.485 188.390 40.675 188.580 ;
        RECT 40.895 188.800 41.085 188.990 ;
        RECT 40.895 188.390 41.085 188.580 ;
        RECT 41.305 188.800 41.495 188.990 ;
        RECT 41.305 188.390 41.495 188.580 ;
        RECT 41.715 188.800 41.905 188.990 ;
        RECT 41.715 188.390 41.905 188.580 ;
        RECT 42.125 188.800 42.315 188.990 ;
        RECT 42.125 188.390 42.315 188.580 ;
        RECT 42.535 188.800 42.725 188.990 ;
        RECT 42.535 188.390 42.725 188.580 ;
        RECT 42.945 188.800 43.135 188.990 ;
        RECT 42.945 188.390 43.135 188.580 ;
        RECT 43.355 188.800 43.545 188.990 ;
        RECT 43.355 188.390 43.545 188.580 ;
        RECT 43.765 188.800 43.955 188.990 ;
        RECT 43.765 188.390 43.955 188.580 ;
        RECT 44.175 188.800 44.365 188.990 ;
        RECT 44.175 188.390 44.365 188.580 ;
        RECT 44.585 188.800 44.775 188.990 ;
        RECT 44.585 188.390 44.775 188.580 ;
        RECT 44.995 188.800 45.185 188.990 ;
        RECT 44.995 188.390 45.185 188.580 ;
      LAYER M1 ;
        RECT 37.400 188.380 45.400 189.000 ;
      LAYER M6 ;
        RECT 37.400 188.380 45.400 189.000 ;
      LAYER V5 ;
        RECT 37.670 188.510 38.030 188.870 ;
        RECT 38.380 188.510 38.740 188.870 ;
        RECT 39.090 188.510 39.450 188.870 ;
        RECT 39.800 188.510 40.160 188.870 ;
        RECT 40.510 188.510 40.870 188.870 ;
        RECT 41.220 188.510 41.580 188.870 ;
        RECT 41.930 188.510 42.290 188.870 ;
        RECT 42.640 188.510 43.000 188.870 ;
        RECT 43.350 188.510 43.710 188.870 ;
        RECT 44.060 188.510 44.420 188.870 ;
        RECT 44.770 188.510 45.130 188.870 ;
      LAYER M5 ;
        RECT 37.400 188.380 45.400 189.000 ;
      LAYER V4 ;
        RECT 37.615 188.800 37.805 188.990 ;
        RECT 37.615 188.390 37.805 188.580 ;
        RECT 38.025 188.800 38.215 188.990 ;
        RECT 38.025 188.390 38.215 188.580 ;
        RECT 38.435 188.800 38.625 188.990 ;
        RECT 38.435 188.390 38.625 188.580 ;
        RECT 38.845 188.800 39.035 188.990 ;
        RECT 38.845 188.390 39.035 188.580 ;
        RECT 39.255 188.800 39.445 188.990 ;
        RECT 39.255 188.390 39.445 188.580 ;
        RECT 39.665 188.800 39.855 188.990 ;
        RECT 39.665 188.390 39.855 188.580 ;
        RECT 40.075 188.800 40.265 188.990 ;
        RECT 40.075 188.390 40.265 188.580 ;
        RECT 40.485 188.800 40.675 188.990 ;
        RECT 40.485 188.390 40.675 188.580 ;
        RECT 40.895 188.800 41.085 188.990 ;
        RECT 40.895 188.390 41.085 188.580 ;
        RECT 41.305 188.800 41.495 188.990 ;
        RECT 41.305 188.390 41.495 188.580 ;
        RECT 41.715 188.800 41.905 188.990 ;
        RECT 41.715 188.390 41.905 188.580 ;
        RECT 42.125 188.800 42.315 188.990 ;
        RECT 42.125 188.390 42.315 188.580 ;
        RECT 42.535 188.800 42.725 188.990 ;
        RECT 42.535 188.390 42.725 188.580 ;
        RECT 42.945 188.800 43.135 188.990 ;
        RECT 42.945 188.390 43.135 188.580 ;
        RECT 43.355 188.800 43.545 188.990 ;
        RECT 43.355 188.390 43.545 188.580 ;
        RECT 43.765 188.800 43.955 188.990 ;
        RECT 43.765 188.390 43.955 188.580 ;
        RECT 44.175 188.800 44.365 188.990 ;
        RECT 44.175 188.390 44.365 188.580 ;
        RECT 44.585 188.800 44.775 188.990 ;
        RECT 44.585 188.390 44.775 188.580 ;
        RECT 44.995 188.800 45.185 188.990 ;
        RECT 44.995 188.390 45.185 188.580 ;
    END
  END CK
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.700 187.775 ;
        RECT 0.130 177.615 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.940 ;
        RECT 0.130 162.140 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 87.910 ;
        RECT 0.130 79.590 0.335 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 78.100 ;
        RECT 0.000 72.380 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 38.500 0.000 41.500 0.700 ;
        RECT 43.510 0.000 49.430 0.700 ;
        RECT 52.530 0.000 58.450 0.700 ;
        RECT 70.570 0.000 76.490 0.700 ;
        RECT 1.100 1.100 78.900 187.900 ;
        RECT 79.300 185.345 79.870 187.775 ;
        RECT 79.300 177.615 79.870 184.955 ;
        RECT 79.300 171.540 79.870 176.940 ;
        RECT 79.300 162.140 79.870 170.040 ;
        RECT 79.300 154.840 79.870 160.610 ;
        RECT 79.300 86.205 79.870 87.960 ;
        RECT 79.665 79.590 79.870 84.480 ;
        RECT 79.300 83.585 79.870 84.480 ;
        RECT 78.500 0.000 80.000 0.700 ;
        RECT 79.300 0.000 80.000 1.820 ;
        RECT 79.500 0.000 80.000 78.100 ;
        RECT 79.300 72.380 80.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.700 187.775 ;
        RECT 0.000 171.540 0.700 176.975 ;
        RECT 0.000 171.540 0.330 184.975 ;
        RECT 0.000 177.580 0.700 184.975 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.335 84.480 ;
        RECT 0.000 84.180 0.700 84.480 ;
        RECT 1.100 1.100 78.900 187.900 ;
        RECT 79.300 185.345 80.000 187.775 ;
        RECT 79.300 171.540 80.000 176.975 ;
        RECT 79.670 171.540 80.000 184.975 ;
        RECT 79.300 177.580 80.000 184.975 ;
        RECT 79.300 162.140 80.000 170.040 ;
        RECT 79.300 85.980 80.000 160.610 ;
        RECT 79.665 79.590 80.000 84.480 ;
        RECT 79.300 83.590 80.000 84.480 ;
        RECT 0.000 0.000 80.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 41.500 0.700 ;
        RECT 78.500 0.000 80.000 0.700 ;
        RECT 0.000 0.000 0.700 78.100 ;
        RECT 79.300 0.000 80.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.700 187.775 ;
        RECT 0.130 177.615 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.940 ;
        RECT 0.130 162.140 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 87.905 ;
        RECT 0.130 79.590 0.335 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 78.100 ;
        RECT 0.000 72.380 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 38.500 0.000 41.500 0.700 ;
        RECT 43.510 0.000 49.430 0.700 ;
        RECT 52.530 0.000 58.450 0.700 ;
        RECT 70.570 0.000 76.490 0.700 ;
        RECT 1.100 1.100 78.900 187.900 ;
        RECT 79.300 185.345 79.870 187.775 ;
        RECT 79.300 177.615 79.870 184.955 ;
        RECT 79.300 171.540 79.870 176.940 ;
        RECT 79.300 162.140 79.870 170.040 ;
        RECT 79.300 154.840 79.870 160.610 ;
        RECT 79.300 86.205 79.870 87.960 ;
        RECT 79.665 79.590 79.870 84.480 ;
        RECT 79.300 83.585 79.870 84.480 ;
        RECT 78.500 0.000 80.000 0.700 ;
        RECT 79.300 0.000 80.000 1.820 ;
        RECT 79.500 0.000 80.000 78.100 ;
        RECT 79.300 72.380 80.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 78.900 187.900 ;
        RECT 79.300 185.015 80.000 187.775 ;
        RECT 79.300 177.615 80.000 184.415 ;
        RECT 79.300 170.640 80.000 176.940 ;
        RECT 79.300 162.140 80.000 170.040 ;
        RECT 79.300 154.840 80.000 161.540 ;
        RECT 79.300 139.530 80.000 150.030 ;
        RECT 79.300 127.890 80.000 136.030 ;
        RECT 79.300 116.930 80.000 124.390 ;
        RECT 79.300 105.930 80.000 113.930 ;
        RECT 79.300 94.290 80.000 102.430 ;
        RECT 79.300 90.340 80.000 92.340 ;
        RECT 79.300 85.080 80.000 87.960 ;
        RECT 79.300 79.590 80.000 84.480 ;
        RECT 79.300 71.440 80.000 79.110 ;
        RECT 79.300 57.770 80.000 68.270 ;
        RECT 79.300 45.630 80.000 54.270 ;
        RECT 79.300 32.770 80.000 42.130 ;
        RECT 79.300 20.470 80.000 28.910 ;
        RECT 79.300 9.130 80.000 16.970 ;
        RECT 79.300 3.610 80.000 5.630 ;
        RECT 0.000 0.000 80.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 79.300 0.000 80.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 78.900 187.900 ;
        RECT 79.300 185.400 80.000 187.775 ;
        RECT 79.300 177.615 80.000 184.955 ;
        RECT 79.300 170.640 80.000 176.940 ;
        RECT 79.300 162.140 80.000 170.040 ;
        RECT 79.300 154.840 80.000 161.540 ;
        RECT 79.300 145.030 80.000 150.030 ;
        RECT 79.300 133.390 80.000 141.530 ;
        RECT 79.300 122.170 80.000 129.890 ;
        RECT 79.300 111.430 80.000 119.170 ;
        RECT 79.300 99.790 80.000 107.930 ;
        RECT 79.300 90.340 80.000 96.290 ;
        RECT 79.300 85.080 80.000 87.960 ;
        RECT 79.300 79.590 80.000 84.780 ;
        RECT 79.300 71.440 80.000 79.110 ;
        RECT 79.300 63.270 80.000 68.270 ;
        RECT 79.300 51.630 80.000 59.770 ;
        RECT 79.300 39.130 80.000 48.130 ;
        RECT 79.300 26.270 80.000 35.270 ;
        RECT 79.300 14.630 80.000 22.770 ;
        RECT 79.300 3.610 80.000 11.130 ;
        RECT 0.000 0.000 80.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 79.300 0.000 80.000 2.960 ;
      LAYER M2 ;
        RECT 0.130 185.345 0.700 187.775 ;
        RECT 0.130 177.615 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.940 ;
        RECT 0.130 162.140 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 87.910 ;
        RECT 0.130 79.590 0.335 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 78.100 ;
        RECT 0.000 72.380 0.700 78.100 ;
        RECT 38.500 0.000 41.500 0.700 ;
        RECT 1.100 1.100 78.900 187.900 ;
        RECT 79.300 185.345 79.870 187.775 ;
        RECT 79.300 177.615 79.870 184.955 ;
        RECT 79.300 171.540 79.870 176.940 ;
        RECT 79.300 162.140 79.870 170.040 ;
        RECT 79.300 154.840 79.870 160.610 ;
        RECT 79.300 86.205 79.870 87.960 ;
        RECT 79.665 79.590 79.870 84.480 ;
        RECT 79.300 83.585 79.870 84.480 ;
        RECT 78.500 0.000 80.000 0.700 ;
        RECT 79.300 0.000 80.000 1.820 ;
        RECT 79.500 0.000 80.000 78.100 ;
        RECT 79.300 72.380 80.000 78.100 ;
  END 
END PSOSC14M

MACRO PSBIAR
  CLASS  PAD ;
  FOREIGN PSBIAR 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
    END
  END P
  PIN AI
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 4.210 188.300 35.790 189.000 ;
      LAYER V3 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M3 ;
        RECT 4.210 188.300 35.790 189.000 ;
      LAYER V2 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M2 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V1 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M1 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER M6 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V5 ;
        RECT 4.555 188.510 4.915 188.870 ;
        RECT 5.265 188.510 5.625 188.870 ;
        RECT 5.975 188.510 6.335 188.870 ;
        RECT 6.685 188.510 7.045 188.870 ;
        RECT 7.395 188.510 7.755 188.870 ;
        RECT 8.105 188.510 8.465 188.870 ;
        RECT 8.815 188.510 9.175 188.870 ;
        RECT 9.525 188.510 9.885 188.870 ;
        RECT 10.235 188.510 10.595 188.870 ;
        RECT 10.945 188.510 11.305 188.870 ;
        RECT 11.655 188.510 12.015 188.870 ;
        RECT 12.365 188.510 12.725 188.870 ;
        RECT 13.075 188.510 13.435 188.870 ;
        RECT 13.785 188.510 14.145 188.870 ;
        RECT 14.495 188.510 14.855 188.870 ;
        RECT 15.205 188.510 15.565 188.870 ;
        RECT 15.915 188.510 16.275 188.870 ;
        RECT 16.625 188.510 16.985 188.870 ;
        RECT 17.335 188.510 17.695 188.870 ;
        RECT 18.045 188.510 18.405 188.870 ;
        RECT 18.755 188.510 19.115 188.870 ;
        RECT 19.465 188.510 19.825 188.870 ;
        RECT 20.175 188.510 20.535 188.870 ;
        RECT 20.885 188.510 21.245 188.870 ;
        RECT 21.595 188.510 21.955 188.870 ;
        RECT 22.305 188.510 22.665 188.870 ;
        RECT 23.015 188.510 23.375 188.870 ;
        RECT 23.725 188.510 24.085 188.870 ;
        RECT 24.435 188.510 24.795 188.870 ;
        RECT 25.145 188.510 25.505 188.870 ;
        RECT 25.855 188.510 26.215 188.870 ;
        RECT 26.565 188.510 26.925 188.870 ;
        RECT 27.275 188.510 27.635 188.870 ;
        RECT 27.985 188.510 28.345 188.870 ;
        RECT 28.695 188.510 29.055 188.870 ;
        RECT 29.405 188.510 29.765 188.870 ;
        RECT 30.115 188.510 30.475 188.870 ;
        RECT 30.825 188.510 31.185 188.870 ;
        RECT 31.535 188.510 31.895 188.870 ;
        RECT 32.245 188.510 32.605 188.870 ;
        RECT 32.955 188.510 33.315 188.870 ;
        RECT 33.665 188.510 34.025 188.870 ;
        RECT 34.375 188.510 34.735 188.870 ;
        RECT 35.085 188.510 35.445 188.870 ;
      LAYER M5 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V4 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
    END
  END AI
  OBS 
      LAYER M4 ;
        RECT 0.130 185.015 0.700 187.775 ;
        RECT 0.130 177.615 0.700 184.415 ;
        RECT 0.130 171.540 0.700 176.940 ;
        RECT 0.130 162.140 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 39.870 187.775 ;
        RECT 39.300 177.615 39.870 184.415 ;
        RECT 39.300 171.540 39.870 176.940 ;
        RECT 39.300 162.140 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.960 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.700 187.775 ;
        RECT 0.000 177.565 0.700 184.975 ;
        RECT 0.000 171.540 0.700 176.885 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 74.720 39.320 77.020 ;
        RECT 39.300 185.345 40.000 187.775 ;
        RECT 39.300 177.565 40.000 184.975 ;
        RECT 39.300 171.540 40.000 176.885 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 85.980 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 74.280 ;
        RECT 0.000 0.000 0.700 76.470 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.800 0.700 78.100 ;
        RECT 39.625 0.000 40.000 78.100 ;
        RECT 39.300 77.800 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.015 0.700 187.775 ;
        RECT 0.130 177.615 0.700 184.415 ;
        RECT 0.130 171.540 0.700 176.940 ;
        RECT 0.130 162.140 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 39.870 187.775 ;
        RECT 39.300 177.615 39.870 184.415 ;
        RECT 39.300 171.540 39.870 176.940 ;
        RECT 39.300 162.140 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 88.860 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.130 185.345 0.700 187.775 ;
        RECT 0.130 177.615 0.700 184.415 ;
        RECT 0.130 171.540 0.700 176.940 ;
        RECT 0.130 162.140 0.700 170.040 ;
        RECT 0.130 153.910 0.700 160.610 ;
        RECT 0.130 86.100 0.700 87.960 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 74.280 ;
        RECT 0.000 72.380 0.700 74.280 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.775 ;
        RECT 39.300 177.615 39.870 184.415 ;
        RECT 39.300 171.540 39.870 176.940 ;
        RECT 39.300 162.140 39.870 170.040 ;
        RECT 39.300 153.915 39.870 160.610 ;
        RECT 39.300 85.980 39.870 88.860 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 74.280 ;
        RECT 39.300 72.300 40.000 74.280 ;
        RECT 39.625 0.000 40.000 78.100 ;
  END 
END PSBIAR

MACRO PSBIA
  CLASS  PAD ;
  FOREIGN PSBIA 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
        RECT 4.210 188.300 35.790 189.000 ;
      LAYER V3 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
        RECT 4.210 188.300 35.790 189.000 ;
      LAYER V2 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M2 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V1 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
      LAYER M1 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER M6 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V5 ;
        RECT 4.555 188.510 4.915 188.870 ;
        RECT 5.265 188.510 5.625 188.870 ;
        RECT 5.975 188.510 6.335 188.870 ;
        RECT 6.685 188.510 7.045 188.870 ;
        RECT 7.395 188.510 7.755 188.870 ;
        RECT 8.105 188.510 8.465 188.870 ;
        RECT 8.815 188.510 9.175 188.870 ;
        RECT 9.525 188.510 9.885 188.870 ;
        RECT 10.235 188.510 10.595 188.870 ;
        RECT 10.945 188.510 11.305 188.870 ;
        RECT 11.655 188.510 12.015 188.870 ;
        RECT 12.365 188.510 12.725 188.870 ;
        RECT 13.075 188.510 13.435 188.870 ;
        RECT 13.785 188.510 14.145 188.870 ;
        RECT 14.495 188.510 14.855 188.870 ;
        RECT 15.205 188.510 15.565 188.870 ;
        RECT 15.915 188.510 16.275 188.870 ;
        RECT 16.625 188.510 16.985 188.870 ;
        RECT 17.335 188.510 17.695 188.870 ;
        RECT 18.045 188.510 18.405 188.870 ;
        RECT 18.755 188.510 19.115 188.870 ;
        RECT 19.465 188.510 19.825 188.870 ;
        RECT 20.175 188.510 20.535 188.870 ;
        RECT 20.885 188.510 21.245 188.870 ;
        RECT 21.595 188.510 21.955 188.870 ;
        RECT 22.305 188.510 22.665 188.870 ;
        RECT 23.015 188.510 23.375 188.870 ;
        RECT 23.725 188.510 24.085 188.870 ;
        RECT 24.435 188.510 24.795 188.870 ;
        RECT 25.145 188.510 25.505 188.870 ;
        RECT 25.855 188.510 26.215 188.870 ;
        RECT 26.565 188.510 26.925 188.870 ;
        RECT 27.275 188.510 27.635 188.870 ;
        RECT 27.985 188.510 28.345 188.870 ;
        RECT 28.695 188.510 29.055 188.870 ;
        RECT 29.405 188.510 29.765 188.870 ;
        RECT 30.115 188.510 30.475 188.870 ;
        RECT 30.825 188.510 31.185 188.870 ;
        RECT 31.535 188.510 31.895 188.870 ;
        RECT 32.245 188.510 32.605 188.870 ;
        RECT 32.955 188.510 33.315 188.870 ;
        RECT 33.665 188.510 34.025 188.870 ;
        RECT 34.375 188.510 34.735 188.870 ;
        RECT 35.085 188.510 35.445 188.870 ;
      LAYER M5 ;
        RECT 4.210 188.380 35.790 189.000 ;
      LAYER V4 ;
        RECT 4.545 188.595 4.735 188.785 ;
        RECT 5.025 188.595 5.215 188.785 ;
        RECT 5.505 188.595 5.695 188.785 ;
        RECT 5.985 188.595 6.175 188.785 ;
        RECT 6.465 188.595 6.655 188.785 ;
        RECT 6.945 188.595 7.135 188.785 ;
        RECT 7.425 188.595 7.615 188.785 ;
        RECT 7.905 188.595 8.095 188.785 ;
        RECT 8.385 188.595 8.575 188.785 ;
        RECT 8.865 188.595 9.055 188.785 ;
        RECT 9.345 188.595 9.535 188.785 ;
        RECT 9.825 188.595 10.015 188.785 ;
        RECT 10.305 188.595 10.495 188.785 ;
        RECT 10.785 188.595 10.975 188.785 ;
        RECT 11.265 188.595 11.455 188.785 ;
        RECT 11.745 188.595 11.935 188.785 ;
        RECT 12.225 188.595 12.415 188.785 ;
        RECT 12.705 188.595 12.895 188.785 ;
        RECT 13.185 188.595 13.375 188.785 ;
        RECT 13.665 188.595 13.855 188.785 ;
        RECT 14.145 188.595 14.335 188.785 ;
        RECT 14.625 188.595 14.815 188.785 ;
        RECT 15.105 188.595 15.295 188.785 ;
        RECT 15.585 188.595 15.775 188.785 ;
        RECT 16.065 188.595 16.255 188.785 ;
        RECT 16.545 188.595 16.735 188.785 ;
        RECT 17.025 188.595 17.215 188.785 ;
        RECT 17.505 188.595 17.695 188.785 ;
        RECT 17.985 188.595 18.175 188.785 ;
        RECT 18.465 188.595 18.655 188.785 ;
        RECT 18.945 188.595 19.135 188.785 ;
        RECT 19.425 188.595 19.615 188.785 ;
        RECT 19.905 188.595 20.095 188.785 ;
        RECT 20.385 188.595 20.575 188.785 ;
        RECT 20.865 188.595 21.055 188.785 ;
        RECT 21.345 188.595 21.535 188.785 ;
        RECT 21.825 188.595 22.015 188.785 ;
        RECT 22.305 188.595 22.495 188.785 ;
        RECT 22.785 188.595 22.975 188.785 ;
        RECT 23.265 188.595 23.455 188.785 ;
        RECT 23.745 188.595 23.935 188.785 ;
        RECT 24.225 188.595 24.415 188.785 ;
        RECT 24.705 188.595 24.895 188.785 ;
        RECT 25.185 188.595 25.375 188.785 ;
        RECT 25.665 188.595 25.855 188.785 ;
        RECT 26.145 188.595 26.335 188.785 ;
        RECT 26.625 188.595 26.815 188.785 ;
        RECT 27.105 188.595 27.295 188.785 ;
        RECT 27.585 188.595 27.775 188.785 ;
        RECT 28.065 188.595 28.255 188.785 ;
        RECT 28.545 188.595 28.735 188.785 ;
        RECT 29.025 188.595 29.215 188.785 ;
        RECT 29.505 188.595 29.695 188.785 ;
        RECT 29.985 188.595 30.175 188.785 ;
        RECT 30.465 188.595 30.655 188.785 ;
        RECT 30.945 188.595 31.135 188.785 ;
        RECT 31.425 188.595 31.615 188.785 ;
        RECT 31.905 188.595 32.095 188.785 ;
        RECT 32.385 188.595 32.575 188.785 ;
        RECT 32.865 188.595 33.055 188.785 ;
        RECT 33.345 188.595 33.535 188.785 ;
        RECT 33.825 188.595 34.015 188.785 ;
        RECT 34.305 188.595 34.495 188.785 ;
        RECT 34.785 188.595 34.975 188.785 ;
        RECT 35.265 188.595 35.455 188.785 ;
    END
  END P
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.700 187.775 ;
        RECT 0.130 177.615 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.940 ;
        RECT 0.130 162.140 0.700 170.040 ;
        RECT 0.130 153.940 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.775 ;
        RECT 39.300 177.615 39.870 184.955 ;
        RECT 39.300 171.540 39.870 176.940 ;
        RECT 39.300 162.140 39.870 170.040 ;
        RECT 39.300 153.910 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.960 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.700 187.775 ;
        RECT 0.000 177.565 0.700 184.975 ;
        RECT 0.000 171.540 0.700 176.885 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 74.720 39.320 77.020 ;
        RECT 39.300 185.345 40.000 187.775 ;
        RECT 39.300 177.565 40.000 184.975 ;
        RECT 39.300 171.540 40.000 176.885 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 85.980 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 74.280 ;
        RECT 0.000 0.000 0.700 76.470 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.800 0.700 78.100 ;
        RECT 39.625 0.000 40.000 78.100 ;
        RECT 39.300 77.800 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.700 187.775 ;
        RECT 0.130 177.615 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.940 ;
        RECT 0.130 162.140 0.700 170.040 ;
        RECT 0.130 153.940 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.775 ;
        RECT 39.300 177.615 39.870 184.955 ;
        RECT 39.300 171.540 39.870 176.940 ;
        RECT 39.300 162.140 39.870 170.040 ;
        RECT 39.300 153.910 39.870 160.610 ;
        RECT 39.300 85.080 39.870 88.860 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.130 185.345 0.700 187.775 ;
        RECT 0.130 177.615 0.700 184.955 ;
        RECT 0.130 171.540 0.700 176.940 ;
        RECT 0.130 162.140 0.700 170.040 ;
        RECT 0.130 153.940 0.700 160.610 ;
        RECT 0.130 86.100 0.700 87.960 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 74.280 ;
        RECT 0.000 72.380 0.700 74.280 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.870 187.775 ;
        RECT 39.300 177.615 39.870 184.955 ;
        RECT 39.300 171.540 39.870 176.940 ;
        RECT 39.300 162.140 39.870 170.040 ;
        RECT 39.300 153.910 39.870 160.610 ;
        RECT 39.300 85.980 39.870 88.860 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 74.280 ;
        RECT 39.300 72.300 40.000 74.280 ;
        RECT 39.625 0.000 40.000 78.100 ;
  END 
END PSBIA

MACRO PSBI24S
  CLASS  PAD ;
  FOREIGN PSBI24S 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V3 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M3 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V2 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M2 ;
        RECT 6.495 188.300 6.695 189.000 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V1 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M1 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER M6 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V5 ;
        RECT 6.435 188.510 6.795 188.870 ;
      LAYER M5 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V4 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V3 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M3 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V2 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M2 ;
        RECT 20.165 188.300 20.775 189.000 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V1 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M1 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER M6 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V5 ;
        RECT 20.310 188.510 20.670 188.870 ;
      LAYER M5 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V4 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V3 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M3 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V2 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M2 ;
        RECT 10.080 188.300 10.280 189.000 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V1 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M1 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER M6 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V5 ;
        RECT 10.020 188.510 10.380 188.870 ;
      LAYER M5 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V4 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V3 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M3 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V2 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M2 ;
        RECT 37.945 188.300 38.145 189.000 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V1 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M1 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER M6 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V5 ;
        RECT 37.885 188.510 38.245 188.870 ;
      LAYER M5 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V4 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V3 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M3 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V2 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M2 ;
        RECT 12.010 188.300 12.210 189.000 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V1 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M1 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER M6 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V5 ;
        RECT 11.950 188.510 12.310 188.870 ;
      LAYER M5 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V4 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V3 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M3 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V2 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M2 ;
        RECT 8.270 188.300 8.470 189.000 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V1 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M1 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER M6 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V5 ;
        RECT 8.190 188.510 8.550 188.870 ;
      LAYER M5 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V4 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V3 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M3 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V2 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M2 ;
        RECT 13.680 188.300 13.880 189.000 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V1 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M1 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER M6 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V5 ;
        RECT 13.620 188.510 13.980 188.870 ;
      LAYER M5 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V4 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V3 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M3 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V2 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M2 ;
        RECT 36.230 188.300 36.430 189.000 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V1 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M1 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER M6 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V5 ;
        RECT 36.170 188.510 36.530 188.870 ;
      LAYER M5 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V4 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.345 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.600 0.700 79.900 ;
        RECT 0.130 79.600 0.330 84.480 ;
        RECT 0.130 84.190 0.700 84.480 ;
        RECT 0.000 0.000 0.500 74.300 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.480 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.375 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 87.960 ;
        RECT 39.670 79.600 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 74.300 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.620 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.000 187.475 0.700 187.775 ;
        RECT 0.000 171.540 0.700 171.805 ;
        RECT 0.000 171.540 0.335 184.975 ;
        RECT 0.000 184.725 0.700 184.975 ;
        RECT 0.590 165.170 0.700 169.020 ;
        RECT 0.000 162.140 0.700 162.440 ;
        RECT 0.000 162.140 0.335 170.040 ;
        RECT 0.000 169.795 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 79.900 ;
        RECT 0.000 79.600 0.335 84.480 ;
        RECT 0.000 81.040 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 74.735 39.400 77.335 ;
        RECT 39.300 74.725 39.390 77.345 ;
        RECT 39.300 74.715 39.380 77.355 ;
        RECT 39.300 74.705 39.370 77.365 ;
        RECT 39.300 74.695 39.360 77.375 ;
        RECT 39.300 74.685 39.350 77.385 ;
        RECT 39.300 74.675 39.340 77.395 ;
        RECT 39.300 74.665 39.330 77.405 ;
        RECT 39.300 74.655 39.320 77.415 ;
        RECT 39.300 74.645 39.310 77.425 ;
        RECT 39.300 186.355 39.340 187.775 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 40.000 187.775 ;
        RECT 39.300 187.475 40.000 187.775 ;
        RECT 39.300 171.540 40.000 171.805 ;
        RECT 39.300 171.540 39.340 180.590 ;
        RECT 39.300 171.540 39.330 181.440 ;
        RECT 39.665 171.540 40.000 184.975 ;
        RECT 39.300 184.725 40.000 184.975 ;
        RECT 39.300 162.140 40.000 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 162.140 39.320 165.910 ;
        RECT 39.300 167.375 39.325 170.040 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.665 162.140 40.000 170.040 ;
        RECT 39.300 169.795 40.000 170.040 ;
        RECT 39.300 85.980 40.000 154.360 ;
        RECT 39.310 85.980 40.000 154.370 ;
        RECT 39.320 85.980 40.000 154.380 ;
        RECT 39.300 156.960 40.000 157.560 ;
        RECT 39.310 156.950 40.000 157.570 ;
        RECT 39.320 156.940 40.000 157.580 ;
        RECT 39.320 160.140 40.000 160.610 ;
        RECT 39.310 160.150 40.000 160.610 ;
        RECT 39.330 85.980 40.000 160.610 ;
        RECT 39.300 160.160 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 74.280 ;
        RECT 0.000 0.000 0.700 74.300 ;
        RECT 0.585 0.000 0.700 76.475 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 39.620 0.000 40.000 78.100 ;
        RECT 39.300 77.770 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.600 0.700 79.900 ;
        RECT 0.130 79.600 0.330 84.480 ;
        RECT 0.130 84.190 0.700 84.480 ;
        RECT 0.000 0.000 0.500 74.300 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.480 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 87.960 ;
        RECT 39.670 79.600 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 74.300 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.620 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.100 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.100 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.335 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.600 0.700 79.900 ;
        RECT 0.130 79.600 0.330 84.480 ;
        RECT 0.130 84.190 0.700 84.480 ;
        RECT 0.000 0.000 0.500 74.300 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.305 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.935 39.330 181.400 ;
        RECT 39.300 74.735 39.400 77.335 ;
        RECT 39.300 74.725 39.390 77.345 ;
        RECT 39.300 74.715 39.380 77.355 ;
        RECT 39.300 74.705 39.370 77.365 ;
        RECT 39.300 74.695 39.360 77.375 ;
        RECT 39.300 74.685 39.350 77.385 ;
        RECT 39.300 74.675 39.340 77.395 ;
        RECT 39.300 74.665 39.330 77.405 ;
        RECT 39.300 74.655 39.320 77.415 ;
        RECT 39.300 74.645 39.310 77.425 ;
        RECT 39.665 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.430 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 87.960 ;
        RECT 39.670 79.600 39.870 84.480 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.900 187.775 ;
        RECT 39.300 187.475 39.900 187.775 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.430 0.000 40.000 74.300 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.625 0.000 40.000 78.100 ;
  END 
END PSBI24S

MACRO PSBI24N
  CLASS  PAD ;
  FOREIGN PSBI24N 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V3 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M3 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V2 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M2 ;
        RECT 6.495 188.300 6.695 189.000 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V1 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M1 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER M6 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V5 ;
        RECT 6.435 188.510 6.795 188.870 ;
      LAYER M5 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V4 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V3 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M3 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V2 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M2 ;
        RECT 20.165 188.300 20.775 189.000 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V1 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M1 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER M6 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V5 ;
        RECT 20.310 188.510 20.670 188.870 ;
      LAYER M5 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V4 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V3 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M3 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V2 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M2 ;
        RECT 10.080 188.300 10.280 189.000 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V1 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M1 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER M6 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V5 ;
        RECT 10.020 188.510 10.380 188.870 ;
      LAYER M5 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V4 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V3 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M3 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V2 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M2 ;
        RECT 37.945 188.300 38.145 189.000 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V1 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M1 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER M6 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V5 ;
        RECT 37.885 188.510 38.245 188.870 ;
      LAYER M5 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V4 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V3 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M3 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V2 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M2 ;
        RECT 12.010 188.300 12.210 189.000 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V1 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M1 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER M6 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V5 ;
        RECT 11.950 188.510 12.310 188.870 ;
      LAYER M5 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V4 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V3 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M3 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V2 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M2 ;
        RECT 8.270 188.300 8.470 189.000 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V1 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M1 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER M6 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V5 ;
        RECT 8.190 188.510 8.550 188.870 ;
      LAYER M5 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V4 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V3 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M3 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V2 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M2 ;
        RECT 13.680 188.300 13.880 189.000 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V1 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M1 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER M6 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V5 ;
        RECT 13.620 188.510 13.980 188.870 ;
      LAYER M5 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V4 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V3 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M3 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V2 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M2 ;
        RECT 36.230 188.300 36.430 189.000 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V1 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M1 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER M6 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V5 ;
        RECT 36.170 188.510 36.530 188.870 ;
      LAYER M5 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V4 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.345 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.600 0.700 79.900 ;
        RECT 0.130 79.600 0.330 84.480 ;
        RECT 0.130 84.190 0.700 84.480 ;
        RECT 0.000 0.000 0.500 74.300 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.480 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.375 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 87.960 ;
        RECT 39.670 79.600 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 74.300 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.620 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.000 187.475 0.700 187.775 ;
        RECT 0.000 171.540 0.700 171.805 ;
        RECT 0.000 171.540 0.335 184.975 ;
        RECT 0.000 184.725 0.700 184.975 ;
        RECT 0.590 163.670 0.700 169.020 ;
        RECT 0.000 162.140 0.700 162.440 ;
        RECT 0.000 162.140 0.335 170.040 ;
        RECT 0.000 169.795 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 79.900 ;
        RECT 0.000 79.600 0.335 84.480 ;
        RECT 0.000 81.040 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 74.735 39.400 77.335 ;
        RECT 39.300 74.725 39.390 77.345 ;
        RECT 39.300 74.715 39.380 77.355 ;
        RECT 39.300 74.705 39.370 77.365 ;
        RECT 39.300 74.695 39.360 77.375 ;
        RECT 39.300 74.685 39.350 77.385 ;
        RECT 39.300 74.675 39.340 77.395 ;
        RECT 39.300 74.665 39.330 77.405 ;
        RECT 39.300 74.655 39.320 77.415 ;
        RECT 39.300 74.645 39.310 77.425 ;
        RECT 39.300 186.355 39.340 187.775 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 40.000 187.775 ;
        RECT 39.300 187.475 40.000 187.775 ;
        RECT 39.300 171.540 40.000 171.805 ;
        RECT 39.300 171.540 39.340 180.590 ;
        RECT 39.300 171.540 39.330 181.440 ;
        RECT 39.665 171.540 40.000 184.975 ;
        RECT 39.300 184.725 40.000 184.975 ;
        RECT 39.300 162.140 40.000 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 162.140 39.320 165.910 ;
        RECT 39.300 167.375 39.325 170.040 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.665 162.140 40.000 170.040 ;
        RECT 39.300 169.795 40.000 170.040 ;
        RECT 39.300 85.980 40.000 154.360 ;
        RECT 39.310 85.980 40.000 154.370 ;
        RECT 39.320 85.980 40.000 154.380 ;
        RECT 39.300 156.960 40.000 157.560 ;
        RECT 39.310 156.950 40.000 157.570 ;
        RECT 39.320 156.940 40.000 157.580 ;
        RECT 39.320 160.140 40.000 160.610 ;
        RECT 39.310 160.150 40.000 160.610 ;
        RECT 39.330 85.980 40.000 160.610 ;
        RECT 39.300 160.160 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 74.280 ;
        RECT 0.000 0.000 0.700 74.300 ;
        RECT 0.585 0.000 0.700 76.475 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 39.620 0.000 40.000 78.100 ;
        RECT 39.300 77.770 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.600 0.700 79.900 ;
        RECT 0.130 79.600 0.330 84.480 ;
        RECT 0.130 84.190 0.700 84.480 ;
        RECT 0.000 0.000 0.500 74.300 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.480 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 87.960 ;
        RECT 39.670 79.600 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 74.300 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.620 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.100 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.100 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.335 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.600 0.700 79.900 ;
        RECT 0.130 79.600 0.330 84.480 ;
        RECT 0.130 84.190 0.700 84.480 ;
        RECT 0.000 0.000 0.500 74.300 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.305 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.935 39.330 181.400 ;
        RECT 39.300 74.735 39.400 77.335 ;
        RECT 39.300 74.725 39.390 77.345 ;
        RECT 39.300 74.715 39.380 77.355 ;
        RECT 39.300 74.705 39.370 77.365 ;
        RECT 39.300 74.695 39.360 77.375 ;
        RECT 39.300 74.685 39.350 77.385 ;
        RECT 39.300 74.675 39.340 77.395 ;
        RECT 39.300 74.665 39.330 77.405 ;
        RECT 39.300 74.655 39.320 77.415 ;
        RECT 39.300 74.645 39.310 77.425 ;
        RECT 39.665 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.430 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 87.960 ;
        RECT 39.670 79.600 39.870 84.480 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.900 187.775 ;
        RECT 39.300 187.475 39.900 187.775 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.430 0.000 40.000 74.300 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.625 0.000 40.000 78.100 ;
  END 
END PSBI24N

MACRO PSBI24F
  CLASS  PAD ;
  FOREIGN PSBI24F 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V3 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M3 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V2 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M2 ;
        RECT 6.495 188.300 6.695 189.000 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V1 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M1 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER M6 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V5 ;
        RECT 6.435 188.510 6.795 188.870 ;
      LAYER M5 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V4 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V3 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M3 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V2 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M2 ;
        RECT 20.165 188.300 20.775 189.000 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V1 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M1 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER M6 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V5 ;
        RECT 20.310 188.510 20.670 188.870 ;
      LAYER M5 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V4 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V3 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M3 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V2 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M2 ;
        RECT 10.080 188.300 10.280 189.000 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V1 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M1 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER M6 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V5 ;
        RECT 10.020 188.510 10.380 188.870 ;
      LAYER M5 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V4 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V3 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M3 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V2 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M2 ;
        RECT 37.945 188.300 38.145 189.000 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V1 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M1 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER M6 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V5 ;
        RECT 37.885 188.510 38.245 188.870 ;
      LAYER M5 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V4 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V3 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M3 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V2 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M2 ;
        RECT 12.010 188.300 12.210 189.000 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V1 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M1 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER M6 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V5 ;
        RECT 11.950 188.510 12.310 188.870 ;
      LAYER M5 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V4 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V3 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M3 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V2 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M2 ;
        RECT 8.270 188.300 8.470 189.000 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V1 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M1 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER M6 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V5 ;
        RECT 8.190 188.510 8.550 188.870 ;
      LAYER M5 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V4 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V3 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M3 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V2 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M2 ;
        RECT 13.680 188.300 13.880 189.000 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V1 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M1 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER M6 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V5 ;
        RECT 13.620 188.510 13.980 188.870 ;
      LAYER M5 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V4 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V3 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M3 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V2 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M2 ;
        RECT 36.230 188.300 36.430 189.000 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V1 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M1 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER M6 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V5 ;
        RECT 36.170 188.510 36.530 188.870 ;
      LAYER M5 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V4 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.345 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.600 0.700 79.900 ;
        RECT 0.130 79.600 0.330 84.480 ;
        RECT 0.130 84.190 0.700 84.480 ;
        RECT 0.000 0.000 0.500 74.300 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.480 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.375 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 87.960 ;
        RECT 39.670 79.600 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 74.300 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.620 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.000 187.475 0.700 187.775 ;
        RECT 0.000 171.540 0.700 171.805 ;
        RECT 0.000 171.540 0.335 184.975 ;
        RECT 0.000 184.725 0.700 184.975 ;
        RECT 0.590 163.110 0.700 169.020 ;
        RECT 0.000 162.140 0.700 162.440 ;
        RECT 0.000 162.140 0.335 170.040 ;
        RECT 0.000 169.795 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 79.900 ;
        RECT 0.000 79.600 0.335 84.480 ;
        RECT 0.000 81.040 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 74.735 39.400 77.335 ;
        RECT 39.300 74.725 39.390 77.345 ;
        RECT 39.300 74.715 39.380 77.355 ;
        RECT 39.300 74.705 39.370 77.365 ;
        RECT 39.300 74.695 39.360 77.375 ;
        RECT 39.300 74.685 39.350 77.385 ;
        RECT 39.300 74.675 39.340 77.395 ;
        RECT 39.300 74.665 39.330 77.405 ;
        RECT 39.300 74.655 39.320 77.415 ;
        RECT 39.300 74.645 39.310 77.425 ;
        RECT 39.300 186.355 39.340 187.775 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 40.000 187.775 ;
        RECT 39.300 187.475 40.000 187.775 ;
        RECT 39.300 171.540 40.000 171.805 ;
        RECT 39.300 171.540 39.340 180.590 ;
        RECT 39.300 171.540 39.330 181.440 ;
        RECT 39.665 171.540 40.000 184.975 ;
        RECT 39.300 184.725 40.000 184.975 ;
        RECT 39.300 162.140 40.000 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 162.140 39.320 165.910 ;
        RECT 39.300 167.375 39.325 170.040 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.665 162.140 40.000 170.040 ;
        RECT 39.300 169.795 40.000 170.040 ;
        RECT 39.300 85.980 40.000 154.360 ;
        RECT 39.310 85.980 40.000 154.370 ;
        RECT 39.320 85.980 40.000 154.380 ;
        RECT 39.300 156.960 40.000 157.560 ;
        RECT 39.310 156.950 40.000 157.570 ;
        RECT 39.320 156.940 40.000 157.580 ;
        RECT 39.320 160.140 40.000 160.610 ;
        RECT 39.310 160.150 40.000 160.610 ;
        RECT 39.330 85.980 40.000 160.610 ;
        RECT 39.300 160.160 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 74.280 ;
        RECT 0.000 0.000 0.700 74.300 ;
        RECT 0.585 0.000 0.700 76.475 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 39.620 0.000 40.000 78.100 ;
        RECT 39.300 77.770 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.600 0.700 79.900 ;
        RECT 0.130 79.600 0.330 84.480 ;
        RECT 0.130 84.190 0.700 84.480 ;
        RECT 0.000 0.000 0.500 74.300 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.480 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 87.960 ;
        RECT 39.670 79.600 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 74.300 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.620 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.100 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.100 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.335 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.040 0.700 87.960 ;
        RECT 0.130 79.600 0.700 79.900 ;
        RECT 0.130 79.600 0.330 84.480 ;
        RECT 0.130 84.190 0.700 84.480 ;
        RECT 0.000 0.000 0.500 74.300 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.305 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.935 39.330 181.400 ;
        RECT 39.300 74.735 39.400 77.335 ;
        RECT 39.300 74.725 39.390 77.345 ;
        RECT 39.300 74.715 39.380 77.355 ;
        RECT 39.300 74.705 39.370 77.365 ;
        RECT 39.300 74.695 39.360 77.375 ;
        RECT 39.300 74.685 39.350 77.385 ;
        RECT 39.300 74.675 39.340 77.395 ;
        RECT 39.300 74.665 39.330 77.405 ;
        RECT 39.300 74.655 39.320 77.415 ;
        RECT 39.300 74.645 39.310 77.425 ;
        RECT 39.665 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.430 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 87.960 ;
        RECT 39.670 79.600 39.870 84.480 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.900 187.775 ;
        RECT 39.300 187.475 39.900 187.775 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.430 0.000 40.000 74.300 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.625 0.000 40.000 78.100 ;
  END 
END PSBI24F

MACRO PSBI16S
  CLASS  PAD ;
  FOREIGN PSBI16S 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V3 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M3 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V2 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M2 ;
        RECT 6.495 188.300 6.695 189.000 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V1 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M1 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER M6 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V5 ;
        RECT 6.435 188.510 6.795 188.870 ;
      LAYER M5 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V4 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V3 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M3 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V2 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M2 ;
        RECT 20.165 188.300 20.775 189.000 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V1 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M1 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER M6 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V5 ;
        RECT 20.310 188.510 20.670 188.870 ;
      LAYER M5 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V4 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V3 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M3 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V2 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M2 ;
        RECT 10.080 188.300 10.280 189.000 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V1 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M1 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER M6 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V5 ;
        RECT 10.020 188.510 10.380 188.870 ;
      LAYER M5 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V4 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V3 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M3 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V2 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M2 ;
        RECT 37.945 188.300 38.145 189.000 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V1 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M1 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER M6 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V5 ;
        RECT 37.885 188.510 38.245 188.870 ;
      LAYER M5 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V4 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V3 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M3 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V2 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M2 ;
        RECT 12.010 188.300 12.210 189.000 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V1 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M1 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER M6 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V5 ;
        RECT 11.950 188.510 12.310 188.870 ;
      LAYER M5 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V4 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V3 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M3 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V2 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M2 ;
        RECT 8.270 188.300 8.470 189.000 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V1 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M1 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER M6 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V5 ;
        RECT 8.190 188.510 8.550 188.870 ;
      LAYER M5 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V4 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V3 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M3 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V2 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M2 ;
        RECT 13.680 188.300 13.880 189.000 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V1 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M1 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER M6 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V5 ;
        RECT 13.620 188.510 13.980 188.870 ;
      LAYER M5 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V4 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V3 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M3 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V2 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M2 ;
        RECT 36.230 188.300 36.430 189.000 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V1 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M1 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER M6 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V5 ;
        RECT 36.170 188.510 36.530 188.870 ;
      LAYER M5 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V4 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.345 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.025 0.700 88.720 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.585 72.380 0.700 77.200 ;
        RECT 0.000 0.000 0.345 78.090 ;
        RECT 0.000 77.760 0.700 78.090 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.375 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 89.160 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.000 187.475 0.700 187.775 ;
        RECT 0.000 171.540 0.700 171.805 ;
        RECT 0.000 171.540 0.335 184.975 ;
        RECT 0.000 184.725 0.700 184.975 ;
        RECT 0.590 165.170 0.700 169.020 ;
        RECT 0.000 162.140 0.700 162.440 ;
        RECT 0.000 162.140 0.335 170.040 ;
        RECT 0.000 169.795 0.700 170.040 ;
        RECT 0.000 85.980 0.700 86.720 ;
        RECT 0.000 85.980 0.330 160.610 ;
        RECT 0.000 154.360 0.700 160.610 ;
        RECT 0.000 79.600 0.700 79.900 ;
        RECT 0.000 79.600 0.335 84.480 ;
        RECT 0.000 81.030 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 74.760 39.400 77.360 ;
        RECT 39.300 74.750 39.390 77.370 ;
        RECT 39.300 74.740 39.380 77.380 ;
        RECT 39.300 74.730 39.370 77.390 ;
        RECT 39.300 74.720 39.360 77.400 ;
        RECT 39.300 74.710 39.350 77.410 ;
        RECT 39.300 74.700 39.340 77.420 ;
        RECT 39.300 74.690 39.330 77.430 ;
        RECT 39.300 74.680 39.320 77.440 ;
        RECT 39.300 74.670 39.310 77.450 ;
        RECT 39.300 186.355 39.340 187.775 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 40.000 187.775 ;
        RECT 39.300 187.475 40.000 187.775 ;
        RECT 39.300 171.540 40.000 171.805 ;
        RECT 39.300 171.540 39.340 180.590 ;
        RECT 39.300 171.540 39.330 181.440 ;
        RECT 39.665 171.540 40.000 184.975 ;
        RECT 39.300 184.725 40.000 184.975 ;
        RECT 39.300 162.140 40.000 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 162.140 39.320 165.910 ;
        RECT 39.300 167.375 39.325 170.040 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.665 162.140 40.000 170.040 ;
        RECT 39.300 169.795 40.000 170.040 ;
        RECT 39.300 85.980 40.000 86.720 ;
        RECT 39.300 153.910 40.000 154.360 ;
        RECT 39.310 153.910 40.000 154.370 ;
        RECT 39.320 153.910 40.000 154.380 ;
        RECT 39.300 156.960 40.000 157.560 ;
        RECT 39.310 156.950 40.000 157.570 ;
        RECT 39.320 156.940 40.000 157.580 ;
        RECT 39.320 160.140 40.000 160.610 ;
        RECT 39.310 160.150 40.000 160.610 ;
        RECT 39.330 85.980 40.000 160.610 ;
        RECT 39.300 160.160 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 74.300 ;
        RECT 39.300 0.000 40.000 74.300 ;
        RECT 0.585 0.000 0.700 76.655 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.800 0.700 78.100 ;
        RECT 39.630 0.000 40.000 78.100 ;
        RECT 39.300 77.800 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.025 0.700 88.720 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.585 72.380 0.700 77.200 ;
        RECT 0.000 0.000 0.345 78.090 ;
        RECT 0.000 77.760 0.700 78.090 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 89.160 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 74.300 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.100 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.100 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.335 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.025 0.700 86.645 ;
        RECT 0.120 86.400 0.700 86.645 ;
        RECT 0.130 86.025 0.610 88.720 ;
        RECT 0.120 86.400 0.610 88.720 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 74.300 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.420 ;
        RECT 0.000 0.000 0.345 78.090 ;
        RECT 0.000 77.760 0.700 78.090 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.935 39.330 181.400 ;
        RECT 39.300 74.760 39.400 77.360 ;
        RECT 39.300 74.750 39.390 77.370 ;
        RECT 39.300 74.740 39.380 77.380 ;
        RECT 39.300 74.730 39.370 77.390 ;
        RECT 39.300 74.720 39.360 77.400 ;
        RECT 39.300 74.710 39.350 77.410 ;
        RECT 39.300 74.700 39.340 77.420 ;
        RECT 39.300 74.690 39.330 77.430 ;
        RECT 39.300 74.680 39.320 77.440 ;
        RECT 39.300 74.670 39.310 77.450 ;
        RECT 39.665 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.430 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 89.160 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.900 187.775 ;
        RECT 39.300 187.475 39.900 187.775 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 74.300 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.640 0.000 40.000 78.100 ;
  END 
END PSBI16S

MACRO PSBI16N
  CLASS  PAD ;
  FOREIGN PSBI16N 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V3 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M3 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V2 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M2 ;
        RECT 6.495 188.300 6.695 189.000 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V1 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M1 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER M6 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V5 ;
        RECT 6.435 188.510 6.795 188.870 ;
      LAYER M5 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V4 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V3 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M3 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V2 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M2 ;
        RECT 20.165 188.300 20.775 189.000 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V1 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M1 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER M6 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V5 ;
        RECT 20.310 188.510 20.670 188.870 ;
      LAYER M5 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V4 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V3 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M3 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V2 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M2 ;
        RECT 10.080 188.300 10.280 189.000 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V1 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M1 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER M6 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V5 ;
        RECT 10.020 188.510 10.380 188.870 ;
      LAYER M5 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V4 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V3 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M3 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V2 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M2 ;
        RECT 37.945 188.300 38.145 189.000 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V1 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M1 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER M6 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V5 ;
        RECT 37.885 188.510 38.245 188.870 ;
      LAYER M5 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V4 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V3 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M3 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V2 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M2 ;
        RECT 12.010 188.300 12.210 189.000 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V1 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M1 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER M6 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V5 ;
        RECT 11.950 188.510 12.310 188.870 ;
      LAYER M5 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V4 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V3 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M3 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V2 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M2 ;
        RECT 8.270 188.300 8.470 189.000 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V1 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M1 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER M6 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V5 ;
        RECT 8.190 188.510 8.550 188.870 ;
      LAYER M5 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V4 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V3 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M3 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V2 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M2 ;
        RECT 13.680 188.300 13.880 189.000 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V1 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M1 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER M6 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V5 ;
        RECT 13.620 188.510 13.980 188.870 ;
      LAYER M5 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V4 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V3 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M3 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V2 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M2 ;
        RECT 36.230 188.300 36.430 189.000 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V1 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M1 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER M6 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V5 ;
        RECT 36.170 188.510 36.530 188.870 ;
      LAYER M5 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V4 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.345 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.025 0.700 88.720 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.585 72.380 0.700 77.200 ;
        RECT 0.000 0.000 0.345 78.090 ;
        RECT 0.000 77.760 0.700 78.090 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.375 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 89.160 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.000 187.475 0.700 187.775 ;
        RECT 0.000 171.540 0.700 171.805 ;
        RECT 0.000 171.540 0.335 184.975 ;
        RECT 0.000 184.725 0.700 184.975 ;
        RECT 0.590 163.670 0.700 169.020 ;
        RECT 0.000 162.140 0.700 162.440 ;
        RECT 0.000 162.140 0.335 170.040 ;
        RECT 0.000 169.795 0.700 170.040 ;
        RECT 0.000 85.980 0.700 86.720 ;
        RECT 0.000 85.980 0.330 160.610 ;
        RECT 0.000 154.360 0.700 160.610 ;
        RECT 0.000 79.600 0.700 79.900 ;
        RECT 0.000 79.600 0.335 84.480 ;
        RECT 0.000 81.030 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 74.760 39.400 77.360 ;
        RECT 39.300 74.750 39.390 77.370 ;
        RECT 39.300 74.740 39.380 77.380 ;
        RECT 39.300 74.730 39.370 77.390 ;
        RECT 39.300 74.720 39.360 77.400 ;
        RECT 39.300 74.710 39.350 77.410 ;
        RECT 39.300 74.700 39.340 77.420 ;
        RECT 39.300 74.690 39.330 77.430 ;
        RECT 39.300 74.680 39.320 77.440 ;
        RECT 39.300 74.670 39.310 77.450 ;
        RECT 39.300 186.355 39.340 187.775 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 40.000 187.775 ;
        RECT 39.300 187.475 40.000 187.775 ;
        RECT 39.300 171.540 40.000 171.805 ;
        RECT 39.300 171.540 39.340 180.590 ;
        RECT 39.300 171.540 39.330 181.440 ;
        RECT 39.665 171.540 40.000 184.975 ;
        RECT 39.300 184.725 40.000 184.975 ;
        RECT 39.300 162.140 40.000 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 162.140 39.320 165.910 ;
        RECT 39.300 167.375 39.325 170.040 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.665 162.140 40.000 170.040 ;
        RECT 39.300 169.795 40.000 170.040 ;
        RECT 39.300 85.980 40.000 86.720 ;
        RECT 39.300 153.910 40.000 154.360 ;
        RECT 39.310 153.910 40.000 154.370 ;
        RECT 39.320 153.910 40.000 154.380 ;
        RECT 39.300 156.960 40.000 157.560 ;
        RECT 39.310 156.950 40.000 157.570 ;
        RECT 39.320 156.940 40.000 157.580 ;
        RECT 39.320 160.140 40.000 160.610 ;
        RECT 39.310 160.150 40.000 160.610 ;
        RECT 39.330 85.980 40.000 160.610 ;
        RECT 39.300 160.160 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 74.300 ;
        RECT 39.300 0.000 40.000 74.300 ;
        RECT 0.585 0.000 0.700 76.655 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.800 0.700 78.100 ;
        RECT 39.630 0.000 40.000 78.100 ;
        RECT 39.300 77.800 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.025 0.700 88.720 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.585 72.380 0.700 77.200 ;
        RECT 0.000 0.000 0.345 78.090 ;
        RECT 0.000 77.760 0.700 78.090 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 89.160 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 74.300 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.100 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.100 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.335 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.025 0.700 86.645 ;
        RECT 0.120 86.400 0.700 86.645 ;
        RECT 0.130 86.025 0.610 88.720 ;
        RECT 0.120 86.400 0.610 88.720 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 74.300 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.420 ;
        RECT 0.000 0.000 0.345 78.090 ;
        RECT 0.000 77.760 0.700 78.090 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.935 39.330 181.400 ;
        RECT 39.300 74.760 39.400 77.360 ;
        RECT 39.300 74.750 39.390 77.370 ;
        RECT 39.300 74.740 39.380 77.380 ;
        RECT 39.300 74.730 39.370 77.390 ;
        RECT 39.300 74.720 39.360 77.400 ;
        RECT 39.300 74.710 39.350 77.410 ;
        RECT 39.300 74.700 39.340 77.420 ;
        RECT 39.300 74.690 39.330 77.430 ;
        RECT 39.300 74.680 39.320 77.440 ;
        RECT 39.300 74.670 39.310 77.450 ;
        RECT 39.665 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.430 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 89.160 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.900 187.775 ;
        RECT 39.300 187.475 39.900 187.775 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 74.300 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.640 0.000 40.000 78.100 ;
  END 
END PSBI16N

MACRO PSBI16F
  CLASS  PAD ;
  FOREIGN PSBI16F 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V3 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M3 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V2 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M2 ;
        RECT 6.495 188.300 6.695 189.000 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V1 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M1 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER M6 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V5 ;
        RECT 6.435 188.510 6.795 188.870 ;
      LAYER M5 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V4 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V3 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M3 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V2 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M2 ;
        RECT 20.165 188.300 20.775 189.000 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V1 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M1 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER M6 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V5 ;
        RECT 20.310 188.510 20.670 188.870 ;
      LAYER M5 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V4 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V3 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M3 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V2 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M2 ;
        RECT 10.080 188.300 10.280 189.000 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V1 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M1 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER M6 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V5 ;
        RECT 10.020 188.510 10.380 188.870 ;
      LAYER M5 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V4 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V3 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M3 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V2 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M2 ;
        RECT 37.945 188.300 38.145 189.000 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V1 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M1 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER M6 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V5 ;
        RECT 37.885 188.510 38.245 188.870 ;
      LAYER M5 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V4 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V3 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M3 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V2 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M2 ;
        RECT 12.010 188.300 12.210 189.000 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V1 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M1 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER M6 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V5 ;
        RECT 11.950 188.510 12.310 188.870 ;
      LAYER M5 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V4 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V3 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M3 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V2 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M2 ;
        RECT 8.270 188.300 8.470 189.000 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V1 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M1 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER M6 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V5 ;
        RECT 8.190 188.510 8.550 188.870 ;
      LAYER M5 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V4 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V3 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M3 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V2 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M2 ;
        RECT 13.680 188.300 13.880 189.000 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V1 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M1 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER M6 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V5 ;
        RECT 13.620 188.510 13.980 188.870 ;
      LAYER M5 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V4 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V3 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M3 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V2 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M2 ;
        RECT 36.230 188.300 36.430 189.000 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V1 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M1 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER M6 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V5 ;
        RECT 36.170 188.510 36.530 188.870 ;
      LAYER M5 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V4 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.345 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.025 0.700 88.720 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.585 72.380 0.700 77.200 ;
        RECT 0.000 0.000 0.345 78.090 ;
        RECT 0.000 77.760 0.700 78.090 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.375 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 89.160 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.000 187.475 0.700 187.775 ;
        RECT 0.000 171.540 0.700 171.805 ;
        RECT 0.000 171.540 0.335 184.975 ;
        RECT 0.000 184.725 0.700 184.975 ;
        RECT 0.590 163.110 0.700 169.020 ;
        RECT 0.000 162.140 0.700 162.440 ;
        RECT 0.000 162.140 0.335 170.040 ;
        RECT 0.000 169.795 0.700 170.040 ;
        RECT 0.000 85.980 0.700 86.720 ;
        RECT 0.000 85.980 0.330 160.610 ;
        RECT 0.000 154.360 0.700 160.610 ;
        RECT 0.000 79.600 0.700 79.900 ;
        RECT 0.000 79.600 0.335 84.480 ;
        RECT 0.000 81.030 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 74.760 39.400 77.360 ;
        RECT 39.300 74.750 39.390 77.370 ;
        RECT 39.300 74.740 39.380 77.380 ;
        RECT 39.300 74.730 39.370 77.390 ;
        RECT 39.300 74.720 39.360 77.400 ;
        RECT 39.300 74.710 39.350 77.410 ;
        RECT 39.300 74.700 39.340 77.420 ;
        RECT 39.300 74.690 39.330 77.430 ;
        RECT 39.300 74.680 39.320 77.440 ;
        RECT 39.300 74.670 39.310 77.450 ;
        RECT 39.300 186.355 39.340 187.775 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 40.000 187.775 ;
        RECT 39.300 187.475 40.000 187.775 ;
        RECT 39.300 171.540 40.000 171.805 ;
        RECT 39.300 171.540 39.340 180.590 ;
        RECT 39.300 171.540 39.330 181.440 ;
        RECT 39.665 171.540 40.000 184.975 ;
        RECT 39.300 184.725 40.000 184.975 ;
        RECT 39.300 162.140 40.000 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 162.140 39.320 165.910 ;
        RECT 39.300 167.375 39.325 170.040 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.665 162.140 40.000 170.040 ;
        RECT 39.300 169.795 40.000 170.040 ;
        RECT 39.300 85.980 40.000 86.720 ;
        RECT 39.300 153.910 40.000 154.360 ;
        RECT 39.310 153.910 40.000 154.370 ;
        RECT 39.320 153.910 40.000 154.380 ;
        RECT 39.300 156.960 40.000 157.560 ;
        RECT 39.310 156.950 40.000 157.570 ;
        RECT 39.320 156.940 40.000 157.580 ;
        RECT 39.320 160.140 40.000 160.610 ;
        RECT 39.310 160.150 40.000 160.610 ;
        RECT 39.330 85.980 40.000 160.610 ;
        RECT 39.300 160.160 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 74.300 ;
        RECT 39.300 0.000 40.000 74.300 ;
        RECT 0.585 0.000 0.700 76.655 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.800 0.700 78.100 ;
        RECT 39.630 0.000 40.000 78.100 ;
        RECT 39.300 77.800 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.025 0.700 88.720 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.585 72.380 0.700 77.200 ;
        RECT 0.000 0.000 0.345 78.090 ;
        RECT 0.000 77.760 0.700 78.090 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 89.160 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 74.300 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.100 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.100 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.335 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.025 0.700 86.645 ;
        RECT 0.120 86.400 0.700 86.645 ;
        RECT 0.130 86.025 0.610 88.720 ;
        RECT 0.120 86.400 0.610 88.720 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 74.300 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.420 ;
        RECT 0.000 0.000 0.345 78.090 ;
        RECT 0.000 77.760 0.700 78.090 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.935 39.330 181.400 ;
        RECT 39.300 74.760 39.400 77.360 ;
        RECT 39.300 74.750 39.390 77.370 ;
        RECT 39.300 74.740 39.380 77.380 ;
        RECT 39.300 74.730 39.370 77.390 ;
        RECT 39.300 74.720 39.360 77.400 ;
        RECT 39.300 74.710 39.350 77.410 ;
        RECT 39.300 74.700 39.340 77.420 ;
        RECT 39.300 74.690 39.330 77.430 ;
        RECT 39.300 74.680 39.320 77.440 ;
        RECT 39.300 74.670 39.310 77.450 ;
        RECT 39.665 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.430 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 89.160 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.900 187.775 ;
        RECT 39.300 187.475 39.900 187.775 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 74.300 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.640 0.000 40.000 78.100 ;
  END 
END PSBI16F

MACRO PSBI8N
  CLASS  PAD ;
  FOREIGN PSBI8N 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V3 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M3 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V2 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M2 ;
        RECT 6.495 188.300 6.695 189.000 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V1 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M1 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER M6 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V5 ;
        RECT 6.435 188.510 6.795 188.870 ;
      LAYER M5 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V4 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V3 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M3 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V2 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M2 ;
        RECT 20.165 188.300 20.775 189.000 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V1 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M1 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER M6 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V5 ;
        RECT 20.310 188.510 20.670 188.870 ;
      LAYER M5 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V4 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V3 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M3 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V2 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M2 ;
        RECT 10.080 188.300 10.280 189.000 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V1 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M1 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER M6 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V5 ;
        RECT 10.020 188.510 10.380 188.870 ;
      LAYER M5 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V4 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V3 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M3 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V2 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M2 ;
        RECT 37.945 188.300 38.145 189.000 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V1 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M1 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER M6 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V5 ;
        RECT 37.885 188.510 38.245 188.870 ;
      LAYER M5 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V4 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V3 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M3 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V2 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M2 ;
        RECT 12.010 188.300 12.210 189.000 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V1 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M1 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER M6 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V5 ;
        RECT 11.950 188.510 12.310 188.870 ;
      LAYER M5 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V4 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V3 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M3 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V2 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M2 ;
        RECT 8.270 188.300 8.470 189.000 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V1 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M1 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER M6 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V5 ;
        RECT 8.190 188.510 8.550 188.870 ;
      LAYER M5 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V4 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V3 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M3 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V2 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M2 ;
        RECT 13.680 188.300 13.880 189.000 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V1 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M1 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER M6 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V5 ;
        RECT 13.620 188.510 13.980 188.870 ;
      LAYER M5 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V4 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V3 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M3 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V2 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M2 ;
        RECT 36.230 188.300 36.430 189.000 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V1 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M1 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER M6 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V5 ;
        RECT 36.170 188.510 36.530 188.870 ;
      LAYER M5 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V4 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.345 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 86.665 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.585 72.380 0.700 77.200 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.375 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.830 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.000 187.475 0.700 187.775 ;
        RECT 0.000 171.540 0.700 171.805 ;
        RECT 0.000 171.540 0.335 184.975 ;
        RECT 0.000 184.725 0.700 184.975 ;
        RECT 0.590 163.670 0.700 169.020 ;
        RECT 0.000 162.140 0.700 162.440 ;
        RECT 0.000 162.140 0.335 170.040 ;
        RECT 0.000 169.795 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 79.900 ;
        RECT 0.000 79.600 0.335 84.480 ;
        RECT 0.000 81.030 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 186.355 39.340 187.775 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 40.000 187.775 ;
        RECT 39.300 187.475 40.000 187.775 ;
        RECT 39.300 171.540 40.000 171.805 ;
        RECT 39.300 171.540 39.340 180.590 ;
        RECT 39.300 171.540 39.330 181.440 ;
        RECT 39.665 171.540 40.000 184.975 ;
        RECT 39.300 184.725 40.000 184.975 ;
        RECT 39.300 162.140 40.000 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 162.140 39.320 165.910 ;
        RECT 39.300 167.375 39.325 170.040 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.665 162.140 40.000 170.040 ;
        RECT 39.300 169.795 40.000 170.040 ;
        RECT 39.300 85.980 40.000 86.720 ;
        RECT 39.300 153.910 40.000 154.360 ;
        RECT 39.310 153.910 40.000 154.370 ;
        RECT 39.320 153.910 40.000 154.380 ;
        RECT 39.300 156.960 40.000 157.560 ;
        RECT 39.310 156.950 40.000 157.570 ;
        RECT 39.320 156.940 40.000 157.580 ;
        RECT 39.320 160.140 40.000 160.610 ;
        RECT 39.310 160.150 40.000 160.610 ;
        RECT 39.330 85.980 40.000 160.610 ;
        RECT 39.300 160.160 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 74.300 ;
        RECT 39.300 0.000 40.000 74.300 ;
        RECT 0.585 0.000 0.700 76.635 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.800 0.700 78.100 ;
        RECT 39.630 0.000 40.000 78.100 ;
        RECT 39.300 77.800 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 86.665 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.585 75.065 0.700 77.200 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.000 0.000 0.360 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.830 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.100 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.100 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.335 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 92.335 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.940 ;
        RECT 0.000 0.000 0.365 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.935 39.330 181.400 ;
        RECT 39.665 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.430 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 92.335 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.900 187.775 ;
        RECT 39.300 187.475 39.900 187.775 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.630 0.000 40.000 75.080 ;
        RECT 39.635 0.000 40.000 78.100 ;
  END 
END PSBI8N

MACRO PSBI8S
  CLASS  PAD ;
  FOREIGN PSBI8S 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V3 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M3 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V2 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M2 ;
        RECT 6.495 188.300 6.695 189.000 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V1 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M1 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER M6 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V5 ;
        RECT 6.435 188.510 6.795 188.870 ;
      LAYER M5 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V4 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V3 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M3 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V2 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M2 ;
        RECT 20.165 188.300 20.775 189.000 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V1 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M1 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER M6 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V5 ;
        RECT 20.310 188.510 20.670 188.870 ;
      LAYER M5 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V4 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V3 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M3 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V2 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M2 ;
        RECT 10.080 188.300 10.280 189.000 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V1 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M1 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER M6 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V5 ;
        RECT 10.020 188.510 10.380 188.870 ;
      LAYER M5 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V4 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V3 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M3 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V2 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M2 ;
        RECT 37.945 188.300 38.145 189.000 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V1 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M1 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER M6 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V5 ;
        RECT 37.885 188.510 38.245 188.870 ;
      LAYER M5 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V4 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V3 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M3 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V2 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M2 ;
        RECT 12.010 188.300 12.210 189.000 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V1 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M1 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER M6 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V5 ;
        RECT 11.950 188.510 12.310 188.870 ;
      LAYER M5 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V4 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V3 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M3 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V2 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M2 ;
        RECT 8.270 188.300 8.470 189.000 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V1 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M1 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER M6 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V5 ;
        RECT 8.190 188.510 8.550 188.870 ;
      LAYER M5 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V4 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V3 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M3 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V2 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M2 ;
        RECT 13.680 188.300 13.880 189.000 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V1 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M1 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER M6 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V5 ;
        RECT 13.620 188.510 13.980 188.870 ;
      LAYER M5 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V4 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V3 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M3 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V2 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M2 ;
        RECT 36.230 188.300 36.430 189.000 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V1 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M1 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER M6 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V5 ;
        RECT 36.170 188.510 36.530 188.870 ;
      LAYER M5 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V4 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.345 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 86.665 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.585 72.380 0.700 77.200 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.375 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.830 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.000 187.475 0.700 187.775 ;
        RECT 0.000 171.540 0.700 171.805 ;
        RECT 0.000 171.540 0.335 184.975 ;
        RECT 0.000 184.725 0.700 184.975 ;
        RECT 0.590 165.170 0.700 169.020 ;
        RECT 0.000 162.140 0.700 162.440 ;
        RECT 0.000 162.140 0.335 170.040 ;
        RECT 0.000 169.795 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 79.900 ;
        RECT 0.000 79.600 0.335 84.480 ;
        RECT 0.000 81.030 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 186.355 39.340 187.775 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 40.000 187.775 ;
        RECT 39.300 187.475 40.000 187.775 ;
        RECT 39.300 171.540 40.000 171.805 ;
        RECT 39.300 171.540 39.340 180.590 ;
        RECT 39.300 171.540 39.330 181.440 ;
        RECT 39.665 171.540 40.000 184.975 ;
        RECT 39.300 184.725 40.000 184.975 ;
        RECT 39.300 162.140 40.000 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 162.140 39.320 165.910 ;
        RECT 39.300 167.375 39.325 170.040 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.665 162.140 40.000 170.040 ;
        RECT 39.300 169.795 40.000 170.040 ;
        RECT 39.300 85.980 40.000 86.720 ;
        RECT 39.300 153.910 40.000 154.360 ;
        RECT 39.310 153.910 40.000 154.370 ;
        RECT 39.320 153.910 40.000 154.380 ;
        RECT 39.300 156.960 40.000 157.560 ;
        RECT 39.310 156.950 40.000 157.570 ;
        RECT 39.320 156.940 40.000 157.580 ;
        RECT 39.320 160.140 40.000 160.610 ;
        RECT 39.310 160.150 40.000 160.610 ;
        RECT 39.330 85.980 40.000 160.610 ;
        RECT 39.300 160.160 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 74.300 ;
        RECT 39.300 0.000 40.000 74.300 ;
        RECT 0.585 0.000 0.700 76.635 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.800 0.700 78.100 ;
        RECT 39.630 0.000 40.000 78.100 ;
        RECT 39.300 77.800 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 86.665 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.585 75.065 0.700 77.200 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.000 0.000 0.360 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.830 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.100 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.100 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.335 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 92.335 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.940 ;
        RECT 0.000 0.000 0.365 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.935 39.330 181.400 ;
        RECT 39.665 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.430 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 92.335 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.900 187.775 ;
        RECT 39.300 187.475 39.900 187.775 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.630 0.000 40.000 75.080 ;
        RECT 39.635 0.000 40.000 78.100 ;
  END 
END PSBI8S

MACRO PSBI8F
  CLASS  PAD ;
  FOREIGN PSBI8F 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V3 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M3 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V2 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M2 ;
        RECT 6.495 188.300 6.695 189.000 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V1 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M1 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER M6 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V5 ;
        RECT 6.435 188.510 6.795 188.870 ;
      LAYER M5 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V4 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V3 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M3 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V2 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M2 ;
        RECT 20.165 188.300 20.775 189.000 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V1 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M1 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER M6 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V5 ;
        RECT 20.310 188.510 20.670 188.870 ;
      LAYER M5 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V4 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V3 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M3 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V2 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M2 ;
        RECT 10.080 188.300 10.280 189.000 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V1 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M1 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER M6 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V5 ;
        RECT 10.020 188.510 10.380 188.870 ;
      LAYER M5 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V4 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V3 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M3 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V2 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M2 ;
        RECT 37.945 188.300 38.145 189.000 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V1 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M1 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER M6 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V5 ;
        RECT 37.885 188.510 38.245 188.870 ;
      LAYER M5 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V4 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V3 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M3 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V2 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M2 ;
        RECT 12.010 188.300 12.210 189.000 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V1 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M1 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER M6 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V5 ;
        RECT 11.950 188.510 12.310 188.870 ;
      LAYER M5 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V4 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V3 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M3 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V2 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M2 ;
        RECT 8.270 188.300 8.470 189.000 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V1 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M1 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER M6 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V5 ;
        RECT 8.190 188.510 8.550 188.870 ;
      LAYER M5 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V4 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V3 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M3 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V2 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M2 ;
        RECT 13.680 188.300 13.880 189.000 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V1 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M1 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER M6 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V5 ;
        RECT 13.620 188.510 13.980 188.870 ;
      LAYER M5 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V4 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V3 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M3 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V2 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M2 ;
        RECT 36.230 188.300 36.430 189.000 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V1 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M1 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER M6 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V5 ;
        RECT 36.170 188.510 36.530 188.870 ;
      LAYER M5 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V4 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.345 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 86.665 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.585 72.380 0.700 77.200 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.375 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.830 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.000 187.475 0.700 187.775 ;
        RECT 0.000 171.540 0.700 171.805 ;
        RECT 0.000 171.540 0.335 184.975 ;
        RECT 0.000 184.725 0.700 184.975 ;
        RECT 0.590 163.110 0.700 169.020 ;
        RECT 0.000 162.140 0.700 162.440 ;
        RECT 0.000 162.140 0.335 170.040 ;
        RECT 0.000 169.795 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 79.900 ;
        RECT 0.000 79.600 0.335 84.480 ;
        RECT 0.000 81.030 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 186.355 39.340 187.775 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 40.000 187.775 ;
        RECT 39.300 187.475 40.000 187.775 ;
        RECT 39.300 171.540 40.000 171.805 ;
        RECT 39.300 171.540 39.340 180.590 ;
        RECT 39.300 171.540 39.330 181.440 ;
        RECT 39.665 171.540 40.000 184.975 ;
        RECT 39.300 184.725 40.000 184.975 ;
        RECT 39.300 162.140 40.000 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 162.140 39.320 165.910 ;
        RECT 39.300 167.375 39.325 170.040 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.665 162.140 40.000 170.040 ;
        RECT 39.300 169.795 40.000 170.040 ;
        RECT 39.300 85.980 40.000 86.720 ;
        RECT 39.300 153.910 40.000 154.360 ;
        RECT 39.310 153.910 40.000 154.370 ;
        RECT 39.320 153.910 40.000 154.380 ;
        RECT 39.300 156.960 40.000 157.560 ;
        RECT 39.310 156.950 40.000 157.570 ;
        RECT 39.320 156.940 40.000 157.580 ;
        RECT 39.320 160.140 40.000 160.610 ;
        RECT 39.310 160.150 40.000 160.610 ;
        RECT 39.330 85.980 40.000 160.610 ;
        RECT 39.300 160.160 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 74.300 ;
        RECT 39.300 0.000 40.000 74.300 ;
        RECT 0.585 0.000 0.700 76.635 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.800 0.700 78.100 ;
        RECT 39.630 0.000 40.000 78.100 ;
        RECT 39.300 77.800 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 86.665 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.585 75.065 0.700 77.200 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.000 0.000 0.360 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.830 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.100 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.100 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.335 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 92.335 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.940 ;
        RECT 0.000 0.000 0.365 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.935 39.330 181.400 ;
        RECT 39.665 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.430 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 92.335 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.900 187.775 ;
        RECT 39.300 187.475 39.900 187.775 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.630 0.000 40.000 75.080 ;
        RECT 39.635 0.000 40.000 78.100 ;
  END 
END PSBI8F

MACRO PSBI4S
  CLASS  PAD ;
  FOREIGN PSBI4S 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V3 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M3 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V2 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M2 ;
        RECT 6.495 188.300 6.695 189.000 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V1 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M1 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER M6 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V5 ;
        RECT 6.435 188.510 6.795 188.870 ;
      LAYER M5 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V4 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V3 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M3 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V2 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M2 ;
        RECT 20.165 188.300 20.775 189.000 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V1 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M1 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER M6 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V5 ;
        RECT 20.310 188.510 20.670 188.870 ;
      LAYER M5 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V4 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V3 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M3 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V2 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M2 ;
        RECT 10.080 188.300 10.280 189.000 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V1 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M1 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER M6 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V5 ;
        RECT 10.020 188.510 10.380 188.870 ;
      LAYER M5 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V4 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V3 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M3 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V2 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M2 ;
        RECT 37.945 188.300 38.145 189.000 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V1 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M1 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER M6 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V5 ;
        RECT 37.885 188.510 38.245 188.870 ;
      LAYER M5 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V4 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V3 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M3 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V2 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M2 ;
        RECT 12.010 188.300 12.210 189.000 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V1 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M1 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER M6 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V5 ;
        RECT 11.950 188.510 12.310 188.870 ;
      LAYER M5 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V4 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V3 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M3 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V2 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M2 ;
        RECT 8.270 188.300 8.470 189.000 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V1 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M1 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER M6 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V5 ;
        RECT 8.190 188.510 8.550 188.870 ;
      LAYER M5 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V4 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V3 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M3 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V2 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M2 ;
        RECT 13.680 188.300 13.880 189.000 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V1 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M1 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER M6 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V5 ;
        RECT 13.620 188.510 13.980 188.870 ;
      LAYER M5 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V4 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V3 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M3 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V2 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M2 ;
        RECT 36.230 188.300 36.430 189.000 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V1 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M1 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER M6 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V5 ;
        RECT 36.170 188.510 36.530 188.870 ;
      LAYER M5 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V4 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.345 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 86.665 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.585 72.380 0.700 77.200 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.375 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.830 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.000 187.475 0.700 187.775 ;
        RECT 0.000 171.540 0.700 171.805 ;
        RECT 0.000 171.540 0.335 184.975 ;
        RECT 0.000 184.725 0.700 184.975 ;
        RECT 0.590 165.170 0.700 169.020 ;
        RECT 0.000 162.140 0.700 162.440 ;
        RECT 0.000 162.140 0.335 170.040 ;
        RECT 0.000 169.795 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 79.900 ;
        RECT 0.000 79.600 0.335 84.480 ;
        RECT 0.000 81.030 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 186.355 39.340 187.775 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 40.000 187.775 ;
        RECT 39.300 187.475 40.000 187.775 ;
        RECT 39.300 171.540 40.000 171.805 ;
        RECT 39.300 171.540 39.340 180.590 ;
        RECT 39.300 171.540 39.330 181.440 ;
        RECT 39.665 171.540 40.000 184.975 ;
        RECT 39.300 184.725 40.000 184.975 ;
        RECT 39.300 162.140 40.000 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 162.140 39.320 165.910 ;
        RECT 39.300 167.375 39.325 170.040 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.665 162.140 40.000 170.040 ;
        RECT 39.300 169.795 40.000 170.040 ;
        RECT 39.300 85.980 40.000 86.720 ;
        RECT 39.300 153.910 40.000 154.360 ;
        RECT 39.310 153.910 40.000 154.370 ;
        RECT 39.320 153.910 40.000 154.380 ;
        RECT 39.300 156.960 40.000 157.560 ;
        RECT 39.310 156.950 40.000 157.570 ;
        RECT 39.320 156.940 40.000 157.580 ;
        RECT 39.320 160.140 40.000 160.610 ;
        RECT 39.310 160.150 40.000 160.610 ;
        RECT 39.330 85.980 40.000 160.610 ;
        RECT 39.300 160.160 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 74.300 ;
        RECT 39.300 0.000 40.000 74.300 ;
        RECT 0.585 0.000 0.700 76.635 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.800 0.700 78.100 ;
        RECT 39.630 0.000 40.000 78.100 ;
        RECT 39.300 77.800 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 86.665 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.585 75.065 0.700 77.200 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.000 0.000 0.360 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.830 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.100 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.100 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.335 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 92.335 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.940 ;
        RECT 0.000 0.000 0.365 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.935 39.330 181.400 ;
        RECT 39.665 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.430 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 92.335 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.900 187.775 ;
        RECT 39.300 187.475 39.900 187.775 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.630 0.000 40.000 75.080 ;
        RECT 39.635 0.000 40.000 78.100 ;
  END 
END PSBI4S

MACRO PSSPLIT40CON
  CLASS  PAD ;
  FOREIGN PSSPLIT40CON 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 162.140 0.700 170.040 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.400 187.775 ;
        RECT 39.300 162.140 39.400 170.040 ;
        RECT 39.300 79.590 39.400 84.480 ;
      LAYER M1 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 162.140 0.700 170.040 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.400 187.775 ;
        RECT 39.300 162.140 39.400 170.040 ;
        RECT 39.300 79.590 39.400 84.480 ;
      LAYER M3 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 162.140 0.700 170.040 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.400 187.775 ;
        RECT 39.300 162.140 39.400 170.040 ;
        RECT 39.300 79.590 39.400 84.480 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 79.590 40.000 84.480 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 79.590 40.000 84.480 ;
      LAYER M2 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 162.140 0.700 170.040 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.400 187.775 ;
        RECT 39.300 162.140 39.400 170.040 ;
        RECT 39.300 79.590 39.400 84.480 ;
  END 
END PSSPLIT40CON

MACRO PSSPLIT40
  CLASS  PAD ;
  FOREIGN PSSPLIT40 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 0.600 162.140 0.700 170.040 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 162.140 39.400 170.040 ;
        RECT 39.300 79.590 39.400 84.480 ;
      LAYER M1 ;
        RECT 0.600 162.140 0.700 170.040 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 162.140 39.400 170.040 ;
        RECT 39.300 79.590 39.400 84.480 ;
      LAYER M3 ;
        RECT 0.600 162.140 0.700 170.040 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 162.140 39.400 170.040 ;
        RECT 39.300 79.590 39.400 84.480 ;
      LAYER M6 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 79.590 40.000 84.480 ;
      LAYER M5 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 79.590 40.000 84.480 ;
      LAYER M2 ;
        RECT 0.600 162.140 0.700 170.040 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 162.140 39.400 170.040 ;
        RECT 39.300 79.590 39.400 84.480 ;
  END 
END PSSPLIT40

MACRO PSFILLER40
  CLASS  PAD ;
  FOREIGN PSFILLER40 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.955 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 86.045 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 0.600 0.000 4.400 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 5.600 0.000 9.400 0.700 ;
        RECT 10.600 0.000 14.400 0.700 ;
        RECT 15.600 0.000 19.400 0.700 ;
        RECT 20.600 0.000 24.400 0.700 ;
        RECT 25.600 0.000 29.400 0.700 ;
        RECT 30.600 0.000 34.400 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.400 187.775 ;
        RECT 39.300 171.540 39.400 184.955 ;
        RECT 39.300 162.140 39.400 170.035 ;
        RECT 39.300 154.840 39.400 160.610 ;
        RECT 39.300 86.045 39.400 87.960 ;
        RECT 39.300 79.590 39.400 84.480 ;
        RECT 35.600 0.000 39.400 0.700 ;
        RECT 39.300 0.000 39.400 78.100 ;
      LAYER M1 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.975 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 85.980 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 0.600 0.000 4.400 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 5.600 0.000 9.400 0.700 ;
        RECT 10.600 0.000 14.400 0.700 ;
        RECT 15.600 0.000 19.400 0.700 ;
        RECT 20.600 0.000 24.400 0.700 ;
        RECT 25.600 0.000 29.400 0.700 ;
        RECT 30.600 0.000 34.400 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.400 187.775 ;
        RECT 39.300 171.540 39.400 184.975 ;
        RECT 39.300 162.140 39.400 170.035 ;
        RECT 39.300 154.840 39.400 160.610 ;
        RECT 39.300 85.980 39.400 87.960 ;
        RECT 39.300 79.590 39.400 84.480 ;
        RECT 35.600 0.000 39.400 0.700 ;
        RECT 39.300 0.000 39.400 78.100 ;
      LAYER M3 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.955 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 86.045 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 0.600 0.000 4.400 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 5.600 0.000 9.400 0.700 ;
        RECT 10.600 0.000 14.400 0.700 ;
        RECT 15.600 0.000 19.400 0.700 ;
        RECT 20.600 0.000 24.400 0.700 ;
        RECT 25.600 0.000 29.400 0.700 ;
        RECT 30.600 0.000 34.400 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.400 187.775 ;
        RECT 39.300 171.540 39.400 184.955 ;
        RECT 39.300 162.140 39.400 170.035 ;
        RECT 39.300 154.840 39.400 160.610 ;
        RECT 39.300 86.045 39.400 87.960 ;
        RECT 39.300 79.590 39.400 84.480 ;
        RECT 35.600 0.000 39.400 0.700 ;
        RECT 39.300 0.000 39.400 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.955 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 86.045 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 0.600 0.000 4.400 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 5.600 0.000 9.400 0.700 ;
        RECT 10.600 0.000 14.400 0.700 ;
        RECT 15.600 0.000 19.400 0.700 ;
        RECT 20.600 0.000 24.400 0.700 ;
        RECT 25.600 0.000 29.400 0.700 ;
        RECT 30.600 0.000 34.400 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.345 39.400 187.775 ;
        RECT 39.300 171.540 39.400 184.955 ;
        RECT 39.300 162.140 39.400 170.035 ;
        RECT 39.300 154.840 39.400 160.610 ;
        RECT 39.300 86.045 39.400 87.960 ;
        RECT 39.300 79.590 39.400 84.480 ;
        RECT 35.600 0.000 39.400 0.700 ;
        RECT 39.300 0.000 39.400 78.100 ;
  END 
END PSFILLER40

MACRO PSFILLER20
  CLASS  PAD ;
  FOREIGN PSFILLER20 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.955 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 86.045 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 0.600 0.000 4.400 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 5.600 0.000 9.400 0.700 ;
        RECT 10.600 0.000 14.400 0.700 ;
        RECT 1.100 1.100 18.900 187.900 ;
        RECT 19.300 185.345 19.400 187.775 ;
        RECT 19.300 171.540 19.400 184.955 ;
        RECT 19.300 162.140 19.400 170.035 ;
        RECT 19.300 154.840 19.400 160.610 ;
        RECT 19.300 86.045 19.400 87.960 ;
        RECT 19.300 79.590 19.400 84.480 ;
        RECT 15.600 0.000 19.400 0.700 ;
        RECT 19.300 0.000 19.400 78.100 ;
      LAYER M1 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.975 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 85.980 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 0.600 0.000 4.400 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 5.600 0.000 9.400 0.700 ;
        RECT 10.600 0.000 14.400 0.700 ;
        RECT 1.100 1.100 18.900 187.900 ;
        RECT 19.300 185.345 19.400 187.775 ;
        RECT 19.300 171.540 19.400 184.975 ;
        RECT 19.300 162.140 19.400 170.035 ;
        RECT 19.300 154.840 19.400 160.610 ;
        RECT 19.300 85.980 19.400 87.960 ;
        RECT 19.300 79.590 19.400 84.480 ;
        RECT 15.600 0.000 19.400 0.700 ;
        RECT 19.300 0.000 19.400 78.100 ;
      LAYER M3 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.955 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 86.045 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 0.600 0.000 4.400 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 5.600 0.000 9.400 0.700 ;
        RECT 10.600 0.000 14.400 0.700 ;
        RECT 1.100 1.100 18.900 187.900 ;
        RECT 19.300 185.345 19.400 187.775 ;
        RECT 19.300 171.540 19.400 184.955 ;
        RECT 19.300 162.140 19.400 170.035 ;
        RECT 19.300 154.840 19.400 160.610 ;
        RECT 19.300 86.045 19.400 87.960 ;
        RECT 19.300 79.590 19.400 84.480 ;
        RECT 15.600 0.000 19.400 0.700 ;
        RECT 19.300 0.000 19.400 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 18.900 187.900 ;
        RECT 19.300 185.015 20.000 187.775 ;
        RECT 19.300 177.615 20.000 184.415 ;
        RECT 19.300 170.640 20.000 176.940 ;
        RECT 19.300 162.140 20.000 170.040 ;
        RECT 19.300 154.840 20.000 161.540 ;
        RECT 19.300 139.530 20.000 150.030 ;
        RECT 19.300 127.890 20.000 136.030 ;
        RECT 19.300 116.930 20.000 124.390 ;
        RECT 19.300 105.930 20.000 113.930 ;
        RECT 19.300 94.290 20.000 102.430 ;
        RECT 19.300 90.340 20.000 92.340 ;
        RECT 19.300 85.080 20.000 87.960 ;
        RECT 19.300 79.590 20.000 84.480 ;
        RECT 19.300 71.440 20.000 79.110 ;
        RECT 19.300 57.770 20.000 68.270 ;
        RECT 19.300 45.630 20.000 54.270 ;
        RECT 19.300 32.770 20.000 42.130 ;
        RECT 19.300 20.470 20.000 28.910 ;
        RECT 19.300 9.130 20.000 16.970 ;
        RECT 19.300 3.610 20.000 5.630 ;
        RECT 0.000 0.000 20.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 19.300 0.000 20.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 18.900 187.900 ;
        RECT 19.300 185.400 20.000 187.775 ;
        RECT 19.300 177.615 20.000 184.955 ;
        RECT 19.300 170.640 20.000 176.940 ;
        RECT 19.300 162.140 20.000 170.040 ;
        RECT 19.300 154.840 20.000 161.540 ;
        RECT 19.300 145.030 20.000 150.030 ;
        RECT 19.300 133.390 20.000 141.530 ;
        RECT 19.300 122.170 20.000 129.890 ;
        RECT 19.300 111.430 20.000 119.170 ;
        RECT 19.300 99.790 20.000 107.930 ;
        RECT 19.300 90.340 20.000 96.290 ;
        RECT 19.300 85.080 20.000 87.960 ;
        RECT 19.300 79.590 20.000 84.480 ;
        RECT 19.300 71.440 20.000 79.110 ;
        RECT 19.300 63.270 20.000 68.270 ;
        RECT 19.300 51.630 20.000 59.770 ;
        RECT 19.300 39.130 20.000 48.130 ;
        RECT 19.300 26.270 20.000 35.270 ;
        RECT 19.300 14.630 20.000 22.770 ;
        RECT 19.300 3.610 20.000 11.130 ;
        RECT 0.000 0.000 20.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 19.300 0.000 20.000 2.960 ;
      LAYER M2 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.955 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 86.045 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 0.600 0.000 4.400 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 5.600 0.000 9.400 0.700 ;
        RECT 10.600 0.000 14.400 0.700 ;
        RECT 1.100 1.100 18.900 187.900 ;
        RECT 19.300 185.345 19.400 187.775 ;
        RECT 19.300 171.540 19.400 184.955 ;
        RECT 19.300 162.140 19.400 170.035 ;
        RECT 19.300 154.840 19.400 160.610 ;
        RECT 19.300 86.045 19.400 87.960 ;
        RECT 19.300 79.590 19.400 84.480 ;
        RECT 15.600 0.000 19.400 0.700 ;
        RECT 19.300 0.000 19.400 78.100 ;
  END 
END PSFILLER20

MACRO PSBI4N
  CLASS  PAD ;
  FOREIGN PSBI4N 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V3 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M3 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V2 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M2 ;
        RECT 6.495 188.300 6.695 189.000 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V1 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M1 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER M6 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V5 ;
        RECT 6.435 188.510 6.795 188.870 ;
      LAYER M5 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V4 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V3 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M3 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V2 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M2 ;
        RECT 20.165 188.300 20.775 189.000 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V1 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M1 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER M6 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V5 ;
        RECT 20.310 188.510 20.670 188.870 ;
      LAYER M5 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V4 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V3 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M3 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V2 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M2 ;
        RECT 10.080 188.300 10.280 189.000 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V1 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M1 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER M6 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V5 ;
        RECT 10.020 188.510 10.380 188.870 ;
      LAYER M5 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V4 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V3 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M3 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V2 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M2 ;
        RECT 37.945 188.300 38.145 189.000 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V1 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M1 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER M6 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V5 ;
        RECT 37.885 188.510 38.245 188.870 ;
      LAYER M5 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V4 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V3 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M3 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V2 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M2 ;
        RECT 12.010 188.300 12.210 189.000 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V1 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M1 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER M6 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V5 ;
        RECT 11.950 188.510 12.310 188.870 ;
      LAYER M5 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V4 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V3 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M3 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V2 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M2 ;
        RECT 8.270 188.300 8.470 189.000 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V1 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M1 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER M6 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V5 ;
        RECT 8.190 188.510 8.550 188.870 ;
      LAYER M5 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V4 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V3 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M3 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V2 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M2 ;
        RECT 13.680 188.300 13.880 189.000 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V1 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M1 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER M6 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V5 ;
        RECT 13.620 188.510 13.980 188.870 ;
      LAYER M5 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V4 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V3 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M3 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V2 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M2 ;
        RECT 36.230 188.300 36.430 189.000 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V1 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M1 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER M6 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V5 ;
        RECT 36.170 188.510 36.530 188.870 ;
      LAYER M5 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V4 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.345 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 86.665 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.585 72.380 0.700 77.200 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.375 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.830 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.000 187.475 0.700 187.775 ;
        RECT 0.000 171.540 0.700 171.805 ;
        RECT 0.000 171.540 0.335 184.975 ;
        RECT 0.000 184.725 0.700 184.975 ;
        RECT 0.590 163.670 0.700 169.020 ;
        RECT 0.000 162.140 0.700 162.440 ;
        RECT 0.000 162.140 0.335 170.040 ;
        RECT 0.000 169.795 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 79.900 ;
        RECT 0.000 79.600 0.335 84.480 ;
        RECT 0.000 81.030 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 186.355 39.340 187.775 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 40.000 187.775 ;
        RECT 39.300 187.475 40.000 187.775 ;
        RECT 39.300 171.540 40.000 171.805 ;
        RECT 39.300 171.540 39.340 180.590 ;
        RECT 39.300 171.540 39.330 181.440 ;
        RECT 39.665 171.540 40.000 184.975 ;
        RECT 39.300 184.725 40.000 184.975 ;
        RECT 39.300 162.140 40.000 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 162.140 39.320 165.910 ;
        RECT 39.300 167.375 39.325 170.040 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.665 162.140 40.000 170.040 ;
        RECT 39.300 169.795 40.000 170.040 ;
        RECT 39.300 85.980 40.000 86.720 ;
        RECT 39.300 153.910 40.000 154.360 ;
        RECT 39.310 153.910 40.000 154.370 ;
        RECT 39.320 153.910 40.000 154.380 ;
        RECT 39.300 156.960 40.000 157.560 ;
        RECT 39.310 156.950 40.000 157.570 ;
        RECT 39.320 156.940 40.000 157.580 ;
        RECT 39.320 160.140 40.000 160.610 ;
        RECT 39.310 160.150 40.000 160.610 ;
        RECT 39.330 85.980 40.000 160.610 ;
        RECT 39.300 160.160 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 74.300 ;
        RECT 39.300 0.000 40.000 74.300 ;
        RECT 0.585 0.000 0.700 76.635 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.800 0.700 78.100 ;
        RECT 39.630 0.000 40.000 78.100 ;
        RECT 39.300 77.800 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 86.665 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.585 75.065 0.700 77.200 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.000 0.000 0.360 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.830 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.100 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.100 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.335 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 92.335 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.940 ;
        RECT 0.000 0.000 0.365 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.935 39.330 181.400 ;
        RECT 39.665 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.430 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 92.335 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.900 187.775 ;
        RECT 39.300 187.475 39.900 187.775 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.630 0.000 40.000 75.080 ;
        RECT 39.635 0.000 40.000 78.100 ;
  END 
END PSBI4N

MACRO PSFILLER10
  CLASS  PAD ;
  FOREIGN PSFILLER10 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.955 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 86.045 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 0.600 0.000 4.400 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 1.100 1.100 8.900 187.900 ;
        RECT 9.300 185.345 9.400 187.775 ;
        RECT 9.300 171.540 9.400 184.955 ;
        RECT 9.300 162.140 9.400 170.035 ;
        RECT 9.300 154.840 9.400 160.610 ;
        RECT 9.300 86.045 9.400 87.960 ;
        RECT 9.300 79.590 9.400 84.480 ;
        RECT 5.600 0.000 9.400 0.700 ;
        RECT 9.300 0.000 9.400 78.100 ;
      LAYER M1 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.975 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 85.980 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 0.600 0.000 4.400 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 1.100 1.100 8.900 187.900 ;
        RECT 9.300 185.345 9.400 187.775 ;
        RECT 9.300 171.540 9.400 184.975 ;
        RECT 9.300 162.140 9.400 170.035 ;
        RECT 9.300 154.840 9.400 160.610 ;
        RECT 9.300 85.980 9.400 87.960 ;
        RECT 9.300 79.590 9.400 84.480 ;
        RECT 5.600 0.000 9.400 0.700 ;
        RECT 9.300 0.000 9.400 78.100 ;
      LAYER M3 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.955 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 86.045 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 0.600 0.000 4.400 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 1.100 1.100 8.900 187.900 ;
        RECT 9.300 185.345 9.400 187.775 ;
        RECT 9.300 171.540 9.400 184.955 ;
        RECT 9.300 162.140 9.400 170.035 ;
        RECT 9.300 154.840 9.400 160.610 ;
        RECT 9.300 86.045 9.400 87.960 ;
        RECT 9.300 79.590 9.400 84.480 ;
        RECT 5.600 0.000 9.400 0.700 ;
        RECT 9.300 0.000 9.400 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 8.900 187.900 ;
        RECT 9.300 185.015 10.000 187.775 ;
        RECT 9.300 177.615 10.000 184.415 ;
        RECT 9.300 170.640 10.000 176.940 ;
        RECT 9.300 162.140 10.000 170.040 ;
        RECT 9.300 154.840 10.000 161.540 ;
        RECT 9.300 90.340 10.000 150.030 ;
        RECT 9.300 85.080 10.000 87.960 ;
        RECT 9.300 79.590 10.000 84.480 ;
        RECT 9.300 71.440 10.000 79.110 ;
        RECT 9.300 3.610 10.000 68.270 ;
        RECT 0.000 0.000 10.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 9.300 0.000 10.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 8.900 187.900 ;
        RECT 9.300 185.400 10.000 187.775 ;
        RECT 9.300 177.615 10.000 184.955 ;
        RECT 9.300 170.640 10.000 176.940 ;
        RECT 9.300 162.140 10.000 170.040 ;
        RECT 9.300 154.840 10.000 161.540 ;
        RECT 9.300 90.340 10.000 150.030 ;
        RECT 9.300 85.080 10.000 87.960 ;
        RECT 9.300 79.590 10.000 84.480 ;
        RECT 9.300 71.440 10.000 79.110 ;
        RECT 9.300 3.610 10.000 68.270 ;
        RECT 0.000 0.000 10.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 9.300 0.000 10.000 2.960 ;
      LAYER M2 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.955 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 86.045 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 0.600 0.000 4.400 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 1.100 1.100 8.900 187.900 ;
        RECT 9.300 185.345 9.400 187.775 ;
        RECT 9.300 171.540 9.400 184.955 ;
        RECT 9.300 162.140 9.400 170.035 ;
        RECT 9.300 154.840 9.400 160.610 ;
        RECT 9.300 86.045 9.400 87.960 ;
        RECT 9.300 79.590 9.400 84.480 ;
        RECT 5.600 0.000 9.400 0.700 ;
        RECT 9.300 0.000 9.400 78.100 ;
  END 
END PSFILLER10

MACRO PSFILLER7_5
  CLASS  PAD ;
  FOREIGN PSFILLER7_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.975 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 85.980 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 1.100 1.100 6.400 187.900 ;
        RECT 6.800 185.345 6.900 187.775 ;
        RECT 6.800 171.540 6.900 184.975 ;
        RECT 6.800 162.140 6.900 170.035 ;
        RECT 6.800 154.840 6.900 160.610 ;
        RECT 6.800 85.980 6.900 87.960 ;
        RECT 6.800 79.590 6.900 84.480 ;
        RECT 0.600 0.000 6.900 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 6.800 0.000 6.900 78.100 ;
      LAYER M1 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.975 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 85.980 0.700 87.960 ;
        RECT 0.600 79.600 0.700 84.480 ;
        RECT 1.100 1.100 6.400 187.900 ;
        RECT 6.800 185.345 6.900 187.775 ;
        RECT 6.800 171.540 6.900 184.975 ;
        RECT 6.800 162.140 6.900 170.035 ;
        RECT 6.800 154.840 6.900 160.610 ;
        RECT 6.800 85.980 6.900 87.960 ;
        RECT 6.800 79.600 6.900 84.480 ;
        RECT 0.600 0.000 6.900 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 6.800 0.000 6.900 78.100 ;
      LAYER M3 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.975 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 85.980 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 1.100 1.100 6.400 187.900 ;
        RECT 6.800 185.345 6.900 187.775 ;
        RECT 6.800 171.540 6.900 184.975 ;
        RECT 6.800 162.140 6.900 170.035 ;
        RECT 6.800 154.840 6.900 160.610 ;
        RECT 6.800 85.980 6.900 87.960 ;
        RECT 6.800 79.590 6.900 84.480 ;
        RECT 0.600 0.000 6.900 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 6.800 0.000 6.900 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 6.400 187.900 ;
        RECT 6.800 185.015 7.500 187.775 ;
        RECT 6.800 177.615 7.500 184.415 ;
        RECT 6.800 170.640 7.500 176.940 ;
        RECT 6.800 162.140 7.500 170.040 ;
        RECT 6.800 154.840 7.500 161.540 ;
        RECT 6.800 139.530 7.500 150.030 ;
        RECT 6.800 127.890 7.500 136.030 ;
        RECT 6.800 116.930 7.500 124.390 ;
        RECT 6.800 105.930 7.500 113.930 ;
        RECT 6.800 94.290 7.500 102.430 ;
        RECT 6.800 90.340 7.500 92.340 ;
        RECT 6.800 85.080 7.500 87.960 ;
        RECT 6.800 79.590 7.500 84.480 ;
        RECT 6.800 71.440 7.500 79.110 ;
        RECT 6.800 57.770 7.500 68.270 ;
        RECT 6.800 45.630 7.500 54.270 ;
        RECT 6.800 32.770 7.500 42.130 ;
        RECT 6.800 20.470 7.500 28.910 ;
        RECT 6.800 9.130 7.500 16.970 ;
        RECT 6.800 3.610 7.500 5.630 ;
        RECT 0.000 0.000 7.500 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 6.800 0.000 7.500 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 6.400 187.900 ;
        RECT 6.800 185.400 7.500 187.775 ;
        RECT 6.800 177.615 7.500 184.955 ;
        RECT 6.800 170.640 7.500 176.940 ;
        RECT 6.800 162.140 7.500 170.040 ;
        RECT 6.800 154.840 7.500 161.540 ;
        RECT 6.800 145.030 7.500 150.030 ;
        RECT 6.800 133.390 7.500 141.530 ;
        RECT 6.800 122.170 7.500 129.890 ;
        RECT 6.800 111.430 7.500 119.170 ;
        RECT 6.800 99.790 7.500 107.930 ;
        RECT 6.800 90.340 7.500 96.290 ;
        RECT 6.800 85.080 7.500 87.960 ;
        RECT 6.800 79.590 7.500 84.480 ;
        RECT 6.800 71.440 7.500 79.110 ;
        RECT 6.800 63.270 7.500 68.270 ;
        RECT 6.800 51.630 7.500 59.770 ;
        RECT 6.800 39.130 7.500 48.130 ;
        RECT 6.800 26.270 7.500 35.270 ;
        RECT 6.800 14.630 7.500 22.770 ;
        RECT 6.800 3.610 7.500 11.130 ;
        RECT 0.000 0.000 7.500 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 6.800 0.000 7.500 2.960 ;
      LAYER M2 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.975 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 85.980 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 1.100 1.100 6.400 187.900 ;
        RECT 6.800 185.345 6.900 187.775 ;
        RECT 6.800 171.540 6.900 184.975 ;
        RECT 6.800 162.140 6.900 170.035 ;
        RECT 6.800 154.840 6.900 160.610 ;
        RECT 6.800 85.980 6.900 87.960 ;
        RECT 6.800 79.590 6.900 84.480 ;
        RECT 0.600 0.000 6.900 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 6.800 0.000 6.900 78.100 ;
  END 
END PSFILLER7_5

MACRO PSFILLER0005
  CLASS  PAD ;
  FOREIGN PSFILLER0005 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.005 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M6 ;
        RECT 0.000 185.015 0.005 187.775 ;
        RECT 0.000 177.615 0.005 184.415 ;
        RECT 0.000 170.640 0.005 176.940 ;
        RECT 0.000 162.140 0.005 170.040 ;
        RECT 0.000 154.840 0.005 161.540 ;
        RECT 0.000 139.530 0.005 150.030 ;
        RECT 0.000 127.890 0.005 136.030 ;
        RECT 0.000 116.930 0.005 124.390 ;
        RECT 0.000 105.930 0.005 113.930 ;
        RECT 0.000 94.290 0.005 102.430 ;
        RECT 0.000 90.340 0.005 92.340 ;
        RECT 0.000 85.080 0.005 87.960 ;
        RECT 0.000 79.590 0.005 84.480 ;
        RECT 0.000 71.440 0.005 79.110 ;
        RECT 0.000 57.770 0.005 68.270 ;
        RECT 0.000 45.630 0.005 54.270 ;
        RECT 0.000 32.770 0.005 42.130 ;
        RECT 0.000 20.470 0.005 28.910 ;
        RECT 0.000 9.130 0.005 16.970 ;
        RECT 0.000 3.610 0.005 5.630 ;
        RECT 0.000 0.000 0.005 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.005 187.775 ;
        RECT 0.000 177.615 0.005 184.955 ;
        RECT 0.000 170.640 0.005 176.940 ;
        RECT 0.000 162.140 0.005 170.040 ;
        RECT 0.000 154.840 0.005 161.540 ;
        RECT 0.000 145.030 0.005 150.030 ;
        RECT 0.000 133.390 0.005 141.530 ;
        RECT 0.000 122.170 0.005 129.890 ;
        RECT 0.000 111.430 0.005 119.170 ;
        RECT 0.000 99.790 0.005 107.930 ;
        RECT 0.000 90.340 0.005 96.290 ;
        RECT 0.000 85.080 0.005 87.960 ;
        RECT 0.000 79.590 0.005 84.480 ;
        RECT 0.000 71.440 0.005 79.110 ;
        RECT 0.000 63.270 0.005 68.270 ;
        RECT 0.000 51.630 0.005 59.770 ;
        RECT 0.000 39.130 0.005 48.130 ;
        RECT 0.000 26.270 0.005 35.270 ;
        RECT 0.000 14.630 0.005 22.770 ;
        RECT 0.000 3.610 0.005 11.130 ;
        RECT 0.000 0.000 0.005 2.960 ;
  END 
END PSFILLER0005

MACRO PSFILLER5
  CLASS  PAD ;
  FOREIGN PSFILLER5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M4 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.955 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 86.045 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 1.100 1.100 3.900 187.900 ;
        RECT 4.300 185.345 4.400 187.775 ;
        RECT 4.300 171.540 4.400 184.955 ;
        RECT 4.300 162.140 4.400 170.035 ;
        RECT 4.300 154.840 4.400 160.610 ;
        RECT 4.300 86.045 4.400 87.960 ;
        RECT 4.300 79.590 4.400 84.480 ;
        RECT 0.600 0.000 4.400 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 4.300 0.000 4.400 78.100 ;
      LAYER M1 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.975 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 85.980 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 1.100 1.100 3.900 187.900 ;
        RECT 4.300 185.345 4.400 187.775 ;
        RECT 4.300 171.540 4.400 184.975 ;
        RECT 4.300 162.140 4.400 170.035 ;
        RECT 4.300 154.840 4.400 160.610 ;
        RECT 4.300 85.980 4.400 87.960 ;
        RECT 4.300 79.590 4.400 84.480 ;
        RECT 0.600 0.000 4.400 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 4.300 0.000 4.400 78.100 ;
      LAYER M3 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.955 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 86.045 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 1.100 1.100 3.900 187.900 ;
        RECT 4.300 185.345 4.400 187.775 ;
        RECT 4.300 171.540 4.400 184.955 ;
        RECT 4.300 162.140 4.400 170.035 ;
        RECT 4.300 154.840 4.400 160.610 ;
        RECT 4.300 86.045 4.400 87.960 ;
        RECT 4.300 79.590 4.400 84.480 ;
        RECT 0.600 0.000 4.400 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 4.300 0.000 4.400 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 3.900 187.900 ;
        RECT 4.300 185.015 5.000 187.775 ;
        RECT 4.300 177.615 5.000 184.415 ;
        RECT 4.300 170.640 5.000 176.940 ;
        RECT 4.300 162.140 5.000 170.040 ;
        RECT 4.300 154.840 5.000 161.540 ;
        RECT 4.300 139.530 5.000 150.030 ;
        RECT 4.300 127.890 5.000 136.030 ;
        RECT 4.300 116.930 5.000 124.390 ;
        RECT 4.300 105.930 5.000 113.930 ;
        RECT 4.300 94.290 5.000 102.430 ;
        RECT 4.300 90.340 5.000 92.340 ;
        RECT 4.300 85.080 5.000 87.960 ;
        RECT 4.300 79.590 5.000 84.480 ;
        RECT 4.300 71.440 5.000 79.110 ;
        RECT 4.300 57.770 5.000 68.270 ;
        RECT 4.300 45.630 5.000 54.270 ;
        RECT 4.300 32.770 5.000 42.130 ;
        RECT 4.300 20.470 5.000 28.910 ;
        RECT 4.300 9.130 5.000 16.970 ;
        RECT 4.300 3.610 5.000 5.630 ;
        RECT 0.000 0.000 5.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 4.300 0.000 5.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 3.900 187.900 ;
        RECT 4.300 185.400 5.000 187.775 ;
        RECT 4.300 177.615 5.000 184.955 ;
        RECT 4.300 170.640 5.000 176.940 ;
        RECT 4.300 162.140 5.000 170.040 ;
        RECT 4.300 154.840 5.000 161.540 ;
        RECT 4.300 145.030 5.000 150.030 ;
        RECT 4.300 133.390 5.000 141.530 ;
        RECT 4.300 122.170 5.000 129.890 ;
        RECT 4.300 111.430 5.000 119.170 ;
        RECT 4.300 99.790 5.000 107.930 ;
        RECT 4.300 90.340 5.000 96.290 ;
        RECT 4.300 85.080 5.000 87.960 ;
        RECT 4.300 79.590 5.000 84.480 ;
        RECT 4.300 71.440 5.000 79.110 ;
        RECT 4.300 63.270 5.000 68.270 ;
        RECT 4.300 51.630 5.000 59.770 ;
        RECT 4.300 39.130 5.000 48.130 ;
        RECT 4.300 26.270 5.000 35.270 ;
        RECT 4.300 14.630 5.000 22.770 ;
        RECT 4.300 3.610 5.000 11.130 ;
        RECT 0.000 0.000 5.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 4.300 0.000 5.000 2.960 ;
      LAYER M2 ;
        RECT 0.600 185.345 0.700 187.775 ;
        RECT 0.600 171.540 0.700 184.955 ;
        RECT 0.600 162.140 0.700 170.035 ;
        RECT 0.600 154.840 0.700 160.610 ;
        RECT 0.600 86.045 0.700 87.960 ;
        RECT 0.600 79.590 0.700 84.480 ;
        RECT 1.100 1.100 3.900 187.900 ;
        RECT 4.300 185.345 4.400 187.775 ;
        RECT 4.300 171.540 4.400 184.955 ;
        RECT 4.300 162.140 4.400 170.035 ;
        RECT 4.300 154.840 4.400 160.610 ;
        RECT 4.300 86.045 4.400 87.960 ;
        RECT 4.300 79.590 4.400 84.480 ;
        RECT 0.600 0.000 4.400 0.700 ;
        RECT 0.600 0.000 0.700 78.100 ;
        RECT 4.300 0.000 4.400 78.100 ;
  END 
END PSFILLER5

MACRO PSFILLER1
  CLASS  PAD ;
  FOREIGN PSFILLER1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M6 ;
        RECT 0.000 185.015 1.000 187.775 ;
        RECT 0.000 177.615 1.000 184.415 ;
        RECT 0.000 170.640 1.000 176.940 ;
        RECT 0.000 162.140 1.000 170.040 ;
        RECT 0.000 154.840 1.000 161.540 ;
        RECT 0.000 139.530 1.000 150.030 ;
        RECT 0.000 127.890 1.000 136.030 ;
        RECT 0.000 116.930 1.000 124.390 ;
        RECT 0.000 105.930 1.000 113.930 ;
        RECT 0.000 94.290 1.000 102.430 ;
        RECT 0.000 90.340 1.000 92.340 ;
        RECT 0.000 85.080 1.000 87.960 ;
        RECT 0.000 79.590 1.000 84.480 ;
        RECT 0.000 71.440 1.000 79.110 ;
        RECT 0.000 57.770 1.000 68.270 ;
        RECT 0.000 45.630 1.000 54.270 ;
        RECT 0.000 32.770 1.000 42.130 ;
        RECT 0.000 20.470 1.000 28.910 ;
        RECT 0.000 9.130 1.000 16.970 ;
        RECT 0.000 3.610 1.000 5.630 ;
        RECT 0.000 0.000 1.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 1.000 187.775 ;
        RECT 0.000 177.615 1.000 184.955 ;
        RECT 0.000 170.640 1.000 176.940 ;
        RECT 0.000 162.140 1.000 170.040 ;
        RECT 0.000 154.840 1.000 161.540 ;
        RECT 0.000 145.030 1.000 150.030 ;
        RECT 0.000 133.390 1.000 141.530 ;
        RECT 0.000 122.170 1.000 129.890 ;
        RECT 0.000 111.430 1.000 119.170 ;
        RECT 0.000 99.790 1.000 107.930 ;
        RECT 0.000 90.340 1.000 96.290 ;
        RECT 0.000 85.080 1.000 87.960 ;
        RECT 0.000 79.590 1.000 84.480 ;
        RECT 0.000 71.440 1.000 79.110 ;
        RECT 0.000 63.270 1.000 68.270 ;
        RECT 0.000 51.630 1.000 59.770 ;
        RECT 0.000 39.130 1.000 48.130 ;
        RECT 0.000 26.270 1.000 35.270 ;
        RECT 0.000 14.630 1.000 22.770 ;
        RECT 0.000 3.610 1.000 11.130 ;
        RECT 0.000 0.000 1.000 2.960 ;
  END 
END PSFILLER1

MACRO PSFILLER01
  CLASS  PAD ;
  FOREIGN PSFILLER01 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.100 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M6 ;
        RECT 0.000 185.015 0.100 187.775 ;
        RECT 0.000 177.615 0.100 184.415 ;
        RECT 0.000 170.640 0.100 176.940 ;
        RECT 0.000 162.140 0.100 170.040 ;
        RECT 0.000 154.840 0.100 161.540 ;
        RECT 0.000 139.530 0.100 150.030 ;
        RECT 0.000 127.890 0.100 136.030 ;
        RECT 0.000 116.930 0.100 124.390 ;
        RECT 0.000 105.930 0.100 113.930 ;
        RECT 0.000 94.290 0.100 102.430 ;
        RECT 0.000 90.340 0.100 92.340 ;
        RECT 0.000 85.080 0.100 87.960 ;
        RECT 0.000 79.590 0.100 84.480 ;
        RECT 0.000 71.440 0.100 79.110 ;
        RECT 0.000 57.770 0.100 68.270 ;
        RECT 0.000 45.630 0.100 54.270 ;
        RECT 0.000 32.770 0.100 42.130 ;
        RECT 0.000 20.470 0.100 28.910 ;
        RECT 0.000 9.130 0.100 16.970 ;
        RECT 0.000 3.610 0.100 5.630 ;
        RECT 0.000 0.000 0.100 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.100 187.775 ;
        RECT 0.000 177.615 0.100 184.955 ;
        RECT 0.000 170.640 0.100 176.940 ;
        RECT 0.000 162.140 0.100 170.040 ;
        RECT 0.000 154.840 0.100 161.540 ;
        RECT 0.000 145.030 0.100 150.030 ;
        RECT 0.000 133.390 0.100 141.530 ;
        RECT 0.000 122.170 0.100 129.890 ;
        RECT 0.000 111.430 0.100 119.170 ;
        RECT 0.000 99.790 0.100 107.930 ;
        RECT 0.000 90.340 0.100 96.290 ;
        RECT 0.000 85.080 0.100 87.960 ;
        RECT 0.000 79.590 0.100 84.480 ;
        RECT 0.000 71.440 0.100 79.110 ;
        RECT 0.000 63.270 0.100 68.270 ;
        RECT 0.000 51.630 0.100 59.770 ;
        RECT 0.000 39.130 0.100 48.130 ;
        RECT 0.000 26.270 0.100 35.270 ;
        RECT 0.000 14.630 0.100 22.770 ;
        RECT 0.000 3.610 0.100 11.130 ;
        RECT 0.000 0.000 0.100 2.960 ;
  END 
END PSFILLER01

MACRO PSFILLER001
  CLASS  PAD ;
  FOREIGN PSFILLER001 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.010 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  OBS 
      LAYER M6 ;
        RECT 0.000 185.015 0.010 187.775 ;
        RECT 0.000 177.615 0.010 184.415 ;
        RECT 0.000 170.640 0.010 176.940 ;
        RECT 0.000 162.140 0.010 170.040 ;
        RECT 0.000 154.840 0.010 161.540 ;
        RECT 0.000 139.530 0.010 150.030 ;
        RECT 0.000 127.890 0.010 136.030 ;
        RECT 0.000 116.930 0.010 124.390 ;
        RECT 0.000 105.930 0.010 113.930 ;
        RECT 0.000 94.290 0.010 102.430 ;
        RECT 0.000 90.340 0.010 92.340 ;
        RECT 0.000 85.080 0.010 87.960 ;
        RECT 0.000 79.590 0.010 84.480 ;
        RECT 0.000 71.440 0.010 79.110 ;
        RECT 0.000 57.770 0.010 68.270 ;
        RECT 0.000 45.630 0.010 54.270 ;
        RECT 0.000 32.770 0.010 42.130 ;
        RECT 0.000 20.470 0.010 28.910 ;
        RECT 0.000 9.130 0.010 16.970 ;
        RECT 0.000 3.610 0.010 5.630 ;
        RECT 0.000 0.000 0.010 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.010 187.775 ;
        RECT 0.000 177.615 0.010 184.955 ;
        RECT 0.000 170.640 0.010 176.940 ;
        RECT 0.000 162.140 0.010 170.040 ;
        RECT 0.000 154.840 0.010 161.540 ;
        RECT 0.000 145.030 0.010 150.030 ;
        RECT 0.000 133.390 0.010 141.530 ;
        RECT 0.000 122.170 0.010 129.890 ;
        RECT 0.000 111.430 0.010 119.170 ;
        RECT 0.000 99.790 0.010 107.930 ;
        RECT 0.000 90.340 0.010 96.290 ;
        RECT 0.000 85.080 0.010 87.960 ;
        RECT 0.000 79.590 0.010 84.480 ;
        RECT 0.000 71.440 0.010 79.110 ;
        RECT 0.000 63.270 0.010 68.270 ;
        RECT 0.000 51.630 0.010 59.770 ;
        RECT 0.000 39.130 0.010 48.130 ;
        RECT 0.000 26.270 0.010 35.270 ;
        RECT 0.000 14.630 0.010 22.770 ;
        RECT 0.000 3.610 0.010 11.130 ;
        RECT 0.000 0.000 0.010 2.960 ;
  END 
END PSFILLER001

MACRO PSBI4F
  CLASS  PAD ;
  FOREIGN PSBI4F 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V3 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M3 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V2 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M2 ;
        RECT 6.495 188.300 6.695 189.000 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V1 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M1 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER M6 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V5 ;
        RECT 6.435 188.510 6.795 188.870 ;
      LAYER M5 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V4 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V3 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M3 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V2 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M2 ;
        RECT 20.165 188.300 20.775 189.000 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V1 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M1 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER M6 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V5 ;
        RECT 20.310 188.510 20.670 188.870 ;
      LAYER M5 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V4 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V3 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M3 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V2 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M2 ;
        RECT 10.080 188.300 10.280 189.000 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V1 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M1 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER M6 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V5 ;
        RECT 10.020 188.510 10.380 188.870 ;
      LAYER M5 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V4 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V3 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M3 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V2 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M2 ;
        RECT 37.945 188.300 38.145 189.000 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V1 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M1 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER M6 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V5 ;
        RECT 37.885 188.510 38.245 188.870 ;
      LAYER M5 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V4 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V3 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M3 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V2 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M2 ;
        RECT 12.010 188.300 12.210 189.000 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V1 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M1 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER M6 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V5 ;
        RECT 11.950 188.510 12.310 188.870 ;
      LAYER M5 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V4 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V3 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M3 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V2 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M2 ;
        RECT 8.270 188.300 8.470 189.000 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V1 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M1 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER M6 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V5 ;
        RECT 8.190 188.510 8.550 188.870 ;
      LAYER M5 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V4 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V3 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M3 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V2 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M2 ;
        RECT 13.680 188.300 13.880 189.000 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V1 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M1 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER M6 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V5 ;
        RECT 13.620 188.510 13.980 188.870 ;
      LAYER M5 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V4 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V3 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M3 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V2 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M2 ;
        RECT 36.230 188.300 36.430 189.000 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V1 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M1 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER M6 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V5 ;
        RECT 36.170 188.510 36.530 188.870 ;
      LAYER M5 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V4 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.345 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 86.665 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.585 72.380 0.700 77.200 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.375 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.830 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.000 187.475 0.700 187.775 ;
        RECT 0.000 171.540 0.700 171.805 ;
        RECT 0.000 171.540 0.335 184.975 ;
        RECT 0.000 184.725 0.700 184.975 ;
        RECT 0.590 163.110 0.700 169.020 ;
        RECT 0.000 162.140 0.700 162.440 ;
        RECT 0.000 162.140 0.335 170.040 ;
        RECT 0.000 169.795 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 79.900 ;
        RECT 0.000 79.600 0.335 84.480 ;
        RECT 0.000 81.030 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 186.355 39.340 187.775 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 40.000 187.775 ;
        RECT 39.300 187.475 40.000 187.775 ;
        RECT 39.300 171.540 40.000 171.805 ;
        RECT 39.300 171.540 39.340 180.590 ;
        RECT 39.300 171.540 39.330 181.440 ;
        RECT 39.665 171.540 40.000 184.975 ;
        RECT 39.300 184.725 40.000 184.975 ;
        RECT 39.300 162.140 40.000 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 162.140 39.320 165.910 ;
        RECT 39.300 167.375 39.325 170.040 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.665 162.140 40.000 170.040 ;
        RECT 39.300 169.795 40.000 170.040 ;
        RECT 39.300 85.980 40.000 86.720 ;
        RECT 39.300 153.910 40.000 154.360 ;
        RECT 39.310 153.910 40.000 154.370 ;
        RECT 39.320 153.910 40.000 154.380 ;
        RECT 39.300 156.960 40.000 157.560 ;
        RECT 39.310 156.950 40.000 157.570 ;
        RECT 39.320 156.940 40.000 157.580 ;
        RECT 39.320 160.140 40.000 160.610 ;
        RECT 39.310 160.150 40.000 160.610 ;
        RECT 39.330 85.980 40.000 160.610 ;
        RECT 39.300 160.160 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 74.300 ;
        RECT 39.300 0.000 40.000 74.300 ;
        RECT 0.585 0.000 0.700 76.635 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.800 0.700 78.100 ;
        RECT 39.630 0.000 40.000 78.100 ;
        RECT 39.300 77.800 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 86.665 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.585 75.065 0.700 77.200 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.000 0.000 0.360 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.830 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.100 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.100 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.335 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 92.335 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.940 ;
        RECT 0.000 0.000 0.365 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.935 39.330 181.400 ;
        RECT 39.665 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.430 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 92.335 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.900 187.775 ;
        RECT 39.300 187.475 39.900 187.775 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.630 0.000 40.000 75.080 ;
        RECT 39.635 0.000 40.000 78.100 ;
  END 
END PSBI4F

MACRO PSBI2F
  CLASS  PAD ;
  FOREIGN PSBI2F 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V3 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M3 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V2 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M2 ;
        RECT 6.495 188.300 6.695 189.000 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V1 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M1 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER M6 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V5 ;
        RECT 6.435 188.510 6.795 188.870 ;
      LAYER M5 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V4 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V3 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M3 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V2 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M2 ;
        RECT 20.165 188.300 20.775 189.000 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V1 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M1 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER M6 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V5 ;
        RECT 20.310 188.510 20.670 188.870 ;
      LAYER M5 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V4 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V3 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M3 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V2 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M2 ;
        RECT 10.080 188.300 10.280 189.000 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V1 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M1 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER M6 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V5 ;
        RECT 10.020 188.510 10.380 188.870 ;
      LAYER M5 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V4 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V3 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M3 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V2 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M2 ;
        RECT 37.945 188.300 38.145 189.000 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V1 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M1 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER M6 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V5 ;
        RECT 37.885 188.510 38.245 188.870 ;
      LAYER M5 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V4 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V3 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M3 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V2 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M2 ;
        RECT 12.010 188.300 12.210 189.000 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V1 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M1 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER M6 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V5 ;
        RECT 11.950 188.510 12.310 188.870 ;
      LAYER M5 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V4 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V3 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M3 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V2 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M2 ;
        RECT 8.270 188.300 8.470 189.000 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V1 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M1 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER M6 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V5 ;
        RECT 8.190 188.510 8.550 188.870 ;
      LAYER M5 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V4 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V3 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M3 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V2 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M2 ;
        RECT 13.680 188.300 13.880 189.000 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V1 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M1 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER M6 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V5 ;
        RECT 13.620 188.510 13.980 188.870 ;
      LAYER M5 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V4 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V3 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M3 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V2 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M2 ;
        RECT 36.230 188.300 36.430 189.000 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V1 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M1 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER M6 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V5 ;
        RECT 36.170 188.510 36.530 188.870 ;
      LAYER M5 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V4 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.345 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 86.665 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.585 72.380 0.700 77.200 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.375 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.830 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.000 187.475 0.700 187.775 ;
        RECT 0.000 171.540 0.700 171.805 ;
        RECT 0.000 171.540 0.335 184.975 ;
        RECT 0.000 184.725 0.700 184.975 ;
        RECT 0.590 163.110 0.700 169.020 ;
        RECT 0.000 162.140 0.700 162.440 ;
        RECT 0.000 162.140 0.335 170.040 ;
        RECT 0.000 169.795 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 79.900 ;
        RECT 0.000 79.600 0.335 84.480 ;
        RECT 0.000 81.030 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 186.355 39.340 187.775 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 40.000 187.775 ;
        RECT 39.300 187.475 40.000 187.775 ;
        RECT 39.300 171.540 40.000 171.805 ;
        RECT 39.300 171.540 39.340 180.590 ;
        RECT 39.300 171.540 39.330 181.440 ;
        RECT 39.665 171.540 40.000 184.975 ;
        RECT 39.300 184.725 40.000 184.975 ;
        RECT 39.300 162.140 40.000 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 162.140 39.320 165.910 ;
        RECT 39.300 167.375 39.325 170.040 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.665 162.140 40.000 170.040 ;
        RECT 39.300 169.795 40.000 170.040 ;
        RECT 39.300 85.980 40.000 86.720 ;
        RECT 39.300 153.910 40.000 154.360 ;
        RECT 39.310 153.910 40.000 154.370 ;
        RECT 39.320 153.910 40.000 154.380 ;
        RECT 39.300 156.960 40.000 157.560 ;
        RECT 39.310 156.950 40.000 157.570 ;
        RECT 39.320 156.940 40.000 157.580 ;
        RECT 39.320 160.140 40.000 160.610 ;
        RECT 39.310 160.150 40.000 160.610 ;
        RECT 39.330 85.980 40.000 160.610 ;
        RECT 39.300 160.160 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 74.300 ;
        RECT 39.300 0.000 40.000 74.300 ;
        RECT 0.585 0.000 0.700 76.635 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.800 0.700 78.100 ;
        RECT 39.630 0.000 40.000 78.100 ;
        RECT 39.300 77.800 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 86.665 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.585 75.065 0.700 77.200 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.000 0.000 0.360 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.830 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.100 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.100 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.335 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 92.335 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.940 ;
        RECT 0.000 0.000 0.365 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.935 39.330 181.400 ;
        RECT 39.665 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.430 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 92.335 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.900 187.775 ;
        RECT 39.300 187.475 39.900 187.775 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.630 0.000 40.000 75.080 ;
        RECT 39.635 0.000 40.000 78.100 ;
  END 
END PSBI2F

MACRO PSBI2S
  CLASS  PAD ;
  FOREIGN PSBI2S 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V3 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M3 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V2 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M2 ;
        RECT 6.495 188.300 6.695 189.000 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V1 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M1 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER M6 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V5 ;
        RECT 6.435 188.510 6.795 188.870 ;
      LAYER M5 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V4 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V3 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M3 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V2 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M2 ;
        RECT 20.165 188.300 20.775 189.000 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V1 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M1 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER M6 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V5 ;
        RECT 20.310 188.510 20.670 188.870 ;
      LAYER M5 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V4 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V3 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M3 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V2 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M2 ;
        RECT 10.080 188.300 10.280 189.000 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V1 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M1 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER M6 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V5 ;
        RECT 10.020 188.510 10.380 188.870 ;
      LAYER M5 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V4 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V3 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M3 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V2 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M2 ;
        RECT 37.945 188.300 38.145 189.000 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V1 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M1 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER M6 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V5 ;
        RECT 37.885 188.510 38.245 188.870 ;
      LAYER M5 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V4 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V3 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M3 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V2 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M2 ;
        RECT 12.010 188.300 12.210 189.000 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V1 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M1 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER M6 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V5 ;
        RECT 11.950 188.510 12.310 188.870 ;
      LAYER M5 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V4 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V3 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M3 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V2 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M2 ;
        RECT 8.270 188.300 8.470 189.000 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V1 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M1 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER M6 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V5 ;
        RECT 8.190 188.510 8.550 188.870 ;
      LAYER M5 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V4 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V3 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M3 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V2 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M2 ;
        RECT 13.680 188.300 13.880 189.000 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V1 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M1 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER M6 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V5 ;
        RECT 13.620 188.510 13.980 188.870 ;
      LAYER M5 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V4 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V3 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M3 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V2 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M2 ;
        RECT 36.230 188.300 36.430 189.000 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V1 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M1 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER M6 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V5 ;
        RECT 36.170 188.510 36.530 188.870 ;
      LAYER M5 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V4 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.345 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 86.665 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.585 72.380 0.700 77.200 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.375 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.830 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.000 187.475 0.700 187.775 ;
        RECT 0.000 171.540 0.700 171.805 ;
        RECT 0.000 171.540 0.335 184.975 ;
        RECT 0.000 184.725 0.700 184.975 ;
        RECT 0.590 165.170 0.700 169.020 ;
        RECT 0.000 162.140 0.700 162.440 ;
        RECT 0.000 162.140 0.335 170.040 ;
        RECT 0.000 169.795 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 79.900 ;
        RECT 0.000 79.600 0.335 84.480 ;
        RECT 0.000 81.030 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 186.355 39.340 187.775 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 40.000 187.775 ;
        RECT 39.300 187.475 40.000 187.775 ;
        RECT 39.300 171.540 40.000 171.805 ;
        RECT 39.300 171.540 39.340 180.590 ;
        RECT 39.300 171.540 39.330 181.440 ;
        RECT 39.665 171.540 40.000 184.975 ;
        RECT 39.300 184.725 40.000 184.975 ;
        RECT 39.300 162.140 40.000 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 162.140 39.320 165.910 ;
        RECT 39.300 167.375 39.325 170.040 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.665 162.140 40.000 170.040 ;
        RECT 39.300 169.795 40.000 170.040 ;
        RECT 39.300 85.980 40.000 86.720 ;
        RECT 39.300 153.910 40.000 154.360 ;
        RECT 39.310 153.910 40.000 154.370 ;
        RECT 39.320 153.910 40.000 154.380 ;
        RECT 39.300 156.960 40.000 157.560 ;
        RECT 39.310 156.950 40.000 157.570 ;
        RECT 39.320 156.940 40.000 157.580 ;
        RECT 39.320 160.140 40.000 160.610 ;
        RECT 39.310 160.150 40.000 160.610 ;
        RECT 39.330 85.980 40.000 160.610 ;
        RECT 39.300 160.160 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 74.300 ;
        RECT 39.300 0.000 40.000 74.300 ;
        RECT 0.585 0.000 0.700 76.635 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.800 0.700 78.100 ;
        RECT 39.630 0.000 40.000 78.100 ;
        RECT 39.300 77.800 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 86.665 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.585 75.065 0.700 77.200 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.000 0.000 0.360 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.830 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.100 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.100 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.335 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 92.335 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.940 ;
        RECT 0.000 0.000 0.365 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.935 39.330 181.400 ;
        RECT 39.665 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.430 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 92.335 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.900 187.775 ;
        RECT 39.300 187.475 39.900 187.775 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.630 0.000 40.000 75.080 ;
        RECT 39.635 0.000 40.000 78.100 ;
  END 
END PSBI2S

MACRO PSBI2N
  CLASS  PAD ;
  FOREIGN PSBI2N 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 189.000 ;
  SYMMETRY R90  ;
  SITE IOSite ;
  PIN P
    DIRECTION INOUT ;
    PORT
      LAYER M4 ;
        RECT 12.530 0.000 18.450 0.700 ;
      LAYER M3 ;
        RECT 12.530 0.000 18.450 0.700 ;
    END
  END P
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V3 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M3 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V2 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M2 ;
        RECT 6.495 188.300 6.695 189.000 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V1 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
      LAYER M1 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER M6 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V5 ;
        RECT 6.435 188.510 6.795 188.870 ;
      LAYER M5 ;
        RECT 6.115 188.380 7.115 189.000 ;
      LAYER V4 ;
        RECT 6.315 188.800 6.505 188.990 ;
        RECT 6.315 188.390 6.505 188.580 ;
        RECT 6.725 188.800 6.915 188.990 ;
        RECT 6.725 188.390 6.915 188.580 ;
    END
  END A
  PIN D
    DIRECTION OUTPUT ;
    PORT
      LAYER M4 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V3 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M3 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V2 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M2 ;
        RECT 20.165 188.300 20.775 189.000 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V1 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
      LAYER M1 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER M6 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V5 ;
        RECT 20.310 188.510 20.670 188.870 ;
      LAYER M5 ;
        RECT 19.990 188.380 20.990 189.000 ;
      LAYER V4 ;
        RECT 20.190 188.800 20.380 188.990 ;
        RECT 20.190 188.390 20.380 188.580 ;
        RECT 20.600 188.800 20.790 188.990 ;
        RECT 20.600 188.390 20.790 188.580 ;
    END
  END D
  PIN PD
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V3 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M3 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V2 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M2 ;
        RECT 10.080 188.300 10.280 189.000 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V1 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
      LAYER M1 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER M6 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V5 ;
        RECT 10.020 188.510 10.380 188.870 ;
      LAYER M5 ;
        RECT 9.700 188.380 10.700 189.000 ;
      LAYER V4 ;
        RECT 9.900 188.800 10.090 188.990 ;
        RECT 9.900 188.390 10.090 188.580 ;
        RECT 10.310 188.800 10.500 188.990 ;
        RECT 10.310 188.390 10.500 188.580 ;
    END
  END PD
  PIN SONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V3 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M3 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V2 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M2 ;
        RECT 37.945 188.300 38.145 189.000 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V1 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
      LAYER M1 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER M6 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V5 ;
        RECT 37.885 188.510 38.245 188.870 ;
      LAYER M5 ;
        RECT 37.565 188.380 38.565 189.000 ;
      LAYER V4 ;
        RECT 37.765 188.800 37.955 188.990 ;
        RECT 37.765 188.390 37.955 188.580 ;
        RECT 38.175 188.800 38.365 188.990 ;
        RECT 38.175 188.390 38.365 188.580 ;
    END
  END SONOF
  PIN PU
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V3 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M3 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V2 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M2 ;
        RECT 12.010 188.300 12.210 189.000 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V1 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
      LAYER M1 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER M6 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V5 ;
        RECT 11.950 188.510 12.310 188.870 ;
      LAYER M5 ;
        RECT 11.630 188.380 12.630 189.000 ;
      LAYER V4 ;
        RECT 11.830 188.800 12.020 188.990 ;
        RECT 11.830 188.390 12.020 188.580 ;
        RECT 12.240 188.800 12.430 188.990 ;
        RECT 12.240 188.390 12.430 188.580 ;
    END
  END PU
  PIN NEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V3 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M3 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V2 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M2 ;
        RECT 8.270 188.300 8.470 189.000 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V1 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
      LAYER M1 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER M6 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V5 ;
        RECT 8.190 188.510 8.550 188.870 ;
      LAYER M5 ;
        RECT 7.870 188.380 8.870 189.000 ;
      LAYER V4 ;
        RECT 8.070 188.800 8.260 188.990 ;
        RECT 8.070 188.390 8.260 188.580 ;
        RECT 8.480 188.800 8.670 188.990 ;
        RECT 8.480 188.390 8.670 188.580 ;
    END
  END NEN
  PIN PEN
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V3 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M3 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V2 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M2 ;
        RECT 13.680 188.300 13.880 189.000 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V1 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
      LAYER M1 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER M6 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V5 ;
        RECT 13.620 188.510 13.980 188.870 ;
      LAYER M5 ;
        RECT 13.300 188.380 14.300 189.000 ;
      LAYER V4 ;
        RECT 13.500 188.800 13.690 188.990 ;
        RECT 13.500 188.390 13.690 188.580 ;
        RECT 13.910 188.800 14.100 188.990 ;
        RECT 13.910 188.390 14.100 188.580 ;
    END
  END PEN
  PIN CONOF
    DIRECTION INPUT ;
    PORT
      LAYER M4 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V3 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M3 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V2 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M2 ;
        RECT 36.230 188.300 36.430 189.000 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V1 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
      LAYER M1 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER M6 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V5 ;
        RECT 36.170 188.510 36.530 188.870 ;
      LAYER M5 ;
        RECT 35.850 188.380 36.850 189.000 ;
      LAYER V4 ;
        RECT 36.050 188.800 36.240 188.990 ;
        RECT 36.050 188.390 36.240 188.580 ;
        RECT 36.460 188.800 36.650 188.990 ;
        RECT 36.460 188.390 36.650 188.580 ;
    END
  END CONOF
  OBS 
      LAYER M4 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.345 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 86.665 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 0.000 0.500 75.080 ;
        RECT 0.000 72.380 0.700 75.080 ;
        RECT 0.585 72.380 0.700 77.200 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.375 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.830 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.300 72.300 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M1 ;
        RECT 0.000 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.000 187.475 0.700 187.775 ;
        RECT 0.000 171.540 0.700 171.805 ;
        RECT 0.000 171.540 0.335 184.975 ;
        RECT 0.000 184.725 0.700 184.975 ;
        RECT 0.590 163.670 0.700 169.020 ;
        RECT 0.000 162.140 0.700 162.440 ;
        RECT 0.000 162.140 0.335 170.040 ;
        RECT 0.000 169.795 0.700 170.040 ;
        RECT 0.000 85.980 0.700 160.610 ;
        RECT 0.000 79.600 0.700 79.900 ;
        RECT 0.000 79.600 0.335 84.480 ;
        RECT 0.000 81.030 0.700 84.480 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 186.355 39.340 187.775 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 40.000 187.775 ;
        RECT 39.300 187.475 40.000 187.775 ;
        RECT 39.300 171.540 40.000 171.805 ;
        RECT 39.300 171.540 39.340 180.590 ;
        RECT 39.300 171.540 39.330 181.440 ;
        RECT 39.665 171.540 40.000 184.975 ;
        RECT 39.300 184.725 40.000 184.975 ;
        RECT 39.300 162.140 40.000 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 162.140 39.320 165.910 ;
        RECT 39.300 167.375 39.325 170.040 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.665 162.140 40.000 170.040 ;
        RECT 39.300 169.795 40.000 170.040 ;
        RECT 39.300 85.980 40.000 86.720 ;
        RECT 39.300 153.910 40.000 154.360 ;
        RECT 39.310 153.910 40.000 154.370 ;
        RECT 39.320 153.910 40.000 154.380 ;
        RECT 39.300 156.960 40.000 157.560 ;
        RECT 39.310 156.950 40.000 157.570 ;
        RECT 39.320 156.940 40.000 157.580 ;
        RECT 39.320 160.140 40.000 160.610 ;
        RECT 39.310 160.150 40.000 160.610 ;
        RECT 39.330 85.980 40.000 160.610 ;
        RECT 39.300 160.160 40.000 160.610 ;
        RECT 39.300 79.600 40.000 79.900 ;
        RECT 39.665 79.600 40.000 84.480 ;
        RECT 39.300 84.180 40.000 84.480 ;
        RECT 0.000 0.000 40.000 0.400 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 74.300 ;
        RECT 39.300 0.000 40.000 74.300 ;
        RECT 0.585 0.000 0.700 76.635 ;
        RECT 0.000 0.000 0.345 78.100 ;
        RECT 0.000 77.800 0.700 78.100 ;
        RECT 39.630 0.000 40.000 78.100 ;
        RECT 39.300 77.800 40.000 78.100 ;
      LAYER M3 ;
        RECT 0.130 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.130 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.330 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 86.665 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.585 75.065 0.700 77.200 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.000 0.000 0.360 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 3.510 0.000 9.430 0.700 ;
        RECT 21.550 0.000 27.470 0.700 ;
        RECT 30.570 0.000 36.490 0.700 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.855 39.330 181.400 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.870 187.775 ;
        RECT 39.300 187.475 39.870 187.775 ;
        RECT 39.670 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.350 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 85.080 39.870 87.830 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.500 0.000 40.000 75.080 ;
        RECT 39.625 0.000 40.000 78.100 ;
      LAYER M6 ;
        RECT 0.000 185.015 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.415 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 139.530 0.700 150.030 ;
        RECT 0.000 127.890 0.700 136.030 ;
        RECT 0.000 116.930 0.700 124.390 ;
        RECT 0.000 105.930 0.700 113.930 ;
        RECT 0.000 94.290 0.700 102.430 ;
        RECT 0.000 90.340 0.700 92.340 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.480 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 57.770 0.700 68.270 ;
        RECT 0.000 45.630 0.700 54.270 ;
        RECT 0.000 32.770 0.700 42.130 ;
        RECT 0.000 20.470 0.700 28.910 ;
        RECT 0.000 9.130 0.700 16.970 ;
        RECT 0.000 3.610 0.700 5.630 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.015 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.415 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 139.530 40.000 150.030 ;
        RECT 39.300 127.890 40.000 136.030 ;
        RECT 39.300 116.930 40.000 124.390 ;
        RECT 39.300 105.930 40.000 113.930 ;
        RECT 39.300 94.290 40.000 102.430 ;
        RECT 39.300 90.340 40.000 92.340 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.480 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 57.770 40.000 68.270 ;
        RECT 39.300 45.630 40.000 54.270 ;
        RECT 39.300 32.770 40.000 42.130 ;
        RECT 39.300 20.470 40.000 28.910 ;
        RECT 39.300 9.130 40.000 16.970 ;
        RECT 39.300 3.610 40.000 5.630 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M5 ;
        RECT 0.000 185.400 0.700 187.775 ;
        RECT 0.000 177.615 0.700 184.955 ;
        RECT 0.000 170.640 0.700 176.940 ;
        RECT 0.000 162.140 0.700 170.040 ;
        RECT 0.000 154.840 0.700 161.540 ;
        RECT 0.000 145.030 0.700 150.030 ;
        RECT 0.000 133.390 0.700 141.530 ;
        RECT 0.000 122.170 0.700 129.890 ;
        RECT 0.000 111.430 0.700 119.170 ;
        RECT 0.000 99.790 0.700 107.930 ;
        RECT 0.000 90.340 0.700 96.290 ;
        RECT 0.000 85.080 0.700 87.960 ;
        RECT 0.000 79.590 0.700 84.780 ;
        RECT 0.000 71.440 0.700 79.110 ;
        RECT 0.000 63.270 0.700 68.270 ;
        RECT 0.000 51.630 0.700 59.770 ;
        RECT 0.000 39.130 0.700 48.130 ;
        RECT 0.000 26.270 0.700 35.270 ;
        RECT 0.000 14.630 0.700 22.770 ;
        RECT 0.000 3.610 0.700 11.130 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 185.400 40.000 187.775 ;
        RECT 39.300 177.615 40.000 184.955 ;
        RECT 39.300 170.640 40.000 176.940 ;
        RECT 39.300 162.140 40.000 170.040 ;
        RECT 39.300 154.840 40.000 161.540 ;
        RECT 39.300 145.030 40.000 150.030 ;
        RECT 39.300 133.390 40.000 141.530 ;
        RECT 39.300 122.170 40.000 129.890 ;
        RECT 39.300 111.430 40.000 119.170 ;
        RECT 39.300 99.790 40.000 107.930 ;
        RECT 39.300 90.340 40.000 96.290 ;
        RECT 39.300 85.080 40.000 87.960 ;
        RECT 39.300 79.590 40.000 84.780 ;
        RECT 39.300 71.440 40.000 79.110 ;
        RECT 39.300 63.270 40.000 68.270 ;
        RECT 39.300 51.630 40.000 59.770 ;
        RECT 39.300 39.130 40.000 48.130 ;
        RECT 39.300 26.270 40.000 35.270 ;
        RECT 39.300 14.630 40.000 22.770 ;
        RECT 39.300 3.610 40.000 11.130 ;
        RECT 0.000 0.000 40.000 0.700 ;
        RECT 0.000 0.000 0.700 2.960 ;
        RECT 39.300 0.000 40.000 2.960 ;
      LAYER M2 ;
        RECT 0.100 185.345 0.330 187.775 ;
        RECT 0.655 186.435 0.700 187.775 ;
        RECT 0.100 187.475 0.700 187.775 ;
        RECT 0.130 178.335 0.335 184.955 ;
        RECT 0.130 184.655 0.700 184.955 ;
        RECT 0.130 171.540 0.700 171.840 ;
        RECT 0.130 171.540 0.330 177.660 ;
        RECT 0.130 162.140 0.700 162.440 ;
        RECT 0.130 162.140 0.330 170.040 ;
        RECT 0.130 169.740 0.700 170.040 ;
        RECT 0.130 154.840 0.700 160.610 ;
        RECT 0.130 86.045 0.700 92.335 ;
        RECT 0.130 79.590 0.700 79.890 ;
        RECT 0.130 79.590 0.330 84.480 ;
        RECT 0.130 84.180 0.700 84.480 ;
        RECT 0.000 0.000 1.500 0.700 ;
        RECT 0.000 0.000 0.700 1.820 ;
        RECT 0.000 72.380 0.700 74.300 ;
        RECT 0.585 72.380 0.700 76.940 ;
        RECT 0.000 0.000 0.365 78.100 ;
        RECT 0.000 77.770 0.700 78.100 ;
        RECT 1.100 1.100 38.900 187.900 ;
        RECT 39.300 178.935 39.330 181.400 ;
        RECT 39.665 178.335 39.870 184.955 ;
        RECT 39.300 184.655 39.870 184.955 ;
        RECT 39.300 171.540 39.870 171.840 ;
        RECT 39.300 171.540 39.340 177.430 ;
        RECT 39.670 171.540 39.870 177.660 ;
        RECT 39.300 162.140 39.870 162.440 ;
        RECT 39.300 162.140 39.360 165.715 ;
        RECT 39.300 167.425 39.360 170.040 ;
        RECT 39.670 162.140 39.870 170.040 ;
        RECT 39.300 169.740 39.870 170.040 ;
        RECT 39.300 154.840 39.870 160.610 ;
        RECT 39.300 86.045 39.870 92.335 ;
        RECT 39.670 79.590 39.870 84.480 ;
        RECT 39.300 186.435 39.350 187.775 ;
        RECT 39.670 185.345 39.900 187.775 ;
        RECT 39.300 187.475 39.900 187.775 ;
        RECT 38.500 0.000 40.000 0.700 ;
        RECT 39.300 0.000 40.000 1.905 ;
        RECT 39.300 72.300 40.000 74.300 ;
        RECT 39.630 0.000 40.000 75.080 ;
        RECT 39.635 0.000 40.000 78.100 ;
  END 
END PSBI2N

END LIBRARY
