module AND2CLKHD1XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2CLKHD2XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2CLKHD3XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2CLKHD4XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2HD1XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2HD1XSPGHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2HD2XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2HD2XSPGHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2HDLXHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2HDMXHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2HDUXHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND3HD1XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module AND3HD2XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module AND3HDLXHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module AND3HDMXHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module AND4HD1XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AND4HD2XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AND4HDLXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AND4HDMXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module ANTFIXHD (Z);
    output Z;

endmodule
module AOI211HD1XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI211HD2XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI211HDLXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI211HDMXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI21B2HD1XHT (Z, AN, BN, C);
    output Z;
    input AN;
    input BN;
    input C;

endmodule
module AOI21B2HD2XHT (Z, AN, BN, C);
    output Z;
    input AN;
    input BN;
    input C;

endmodule
module AOI21B2HDLXHT (Z, AN, BN, C);
    output Z;
    input AN;
    input BN;
    input C;

endmodule
module AOI21B2HDMXHT (Z, AN, BN, C);
    output Z;
    input AN;
    input BN;
    input C;

endmodule
module AOI21HD1XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module AOI21HD2XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module AOI21HDLXHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module AOI21HDMXHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module AOI21HDUXHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module AOI221HD1XHT (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module AOI221HD2XHT (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module AOI221HDLXHT (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module AOI221HDMXHT (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module AOI222HD1XHT (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module AOI222HD2XHT (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module AOI222HDLXHT (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module AOI222HDMXHT (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module AOI22B2HD1XHT (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module AOI22B2HD2XHT (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module AOI22B2HDLXHT (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module AOI22B2HDMXHT (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module AOI22HD1XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI22HD2XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI22HDLXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI22HDMXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI22HDUXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI31HD1XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI31HD2XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI31HDLXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI31HDMXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI32HD1XHT (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module AOI32HD2XHT (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module AOI32HDLXHT (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module AOI32HDMXHT (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module AOI33HD1XHT (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module AOI33HD2XHT (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module AOI33HDLXHT (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module AOI33HDMXHT (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module BUFCLKHD10XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD12XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD14XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD16XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD1XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD20XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD2XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD30XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD3XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD40XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD4XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD5XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD6XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD7XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD80XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD8XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHDLXHT (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHDMXHT (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHDUXHT (Z, A);
    output Z;
    input A;

endmodule
module BUFHD12XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFHD16XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFHD1XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFHD20XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFHD2XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFHD3XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFHD4XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFHD5XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFHD6XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFHD7XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFHD8XHT (Z, A);
    output Z;
    input A;

endmodule
module BUFHD8XSPGHT (Z, A);
    output Z;
    input A;

endmodule
module BUFHDLXHT (Z, A);
    output Z;
    input A;

endmodule
module BUFHDMXHT (Z, A);
    output Z;
    input A;

endmodule
module BUFHDUXHT (Z, A);
    output Z;
    input A;

endmodule
module BUFTSHD12XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD16XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD1XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD20XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD2XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD3XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD4XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD5XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD6XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD7XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD8XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHDLXHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHDMXHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHDUXHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module DEL1HD1XHT (Z, A);
    output Z;
    input A;

endmodule
module DEL1HDMXHT (Z, A);
    output Z;
    input A;

endmodule
module DEL1HDMXSPGHT (Z, A);
    output Z;
    input A;

endmodule
module DEL2HD1XHT (Z, A);
    output Z;
    input A;

endmodule
module DEL2HDMXHT (Z, A);
    output Z;
    input A;

endmodule
module DEL2HDMXSPGHT (Z, A);
    output Z;
    input A;

endmodule
module DEL3HD1XHT (Z, A);
    output Z;
    input A;

endmodule
module DEL3HDMXHT (Z, A);
    output Z;
    input A;

endmodule
module DEL4HD1XHT (Z, A);
    output Z;
    input A;

endmodule
module DEL4HDMXHT (Z, A);
    output Z;
    input A;

endmodule
module DEL4HDMXSPGHT (Z, A);
    output Z;
    input A;

endmodule
module FAHD1XHT (CO, S, A, B, CI);
    output CO;
    output S;
    input A;
    input B;
    input CI;

endmodule
module FAHD2XHT (CO, S, A, B, CI);
    output CO;
    output S;
    input A;
    input B;
    input CI;

endmodule
module FAHDLXHT (CO, S, A, B, CI);
    output CO;
    output S;
    input A;
    input B;
    input CI;

endmodule
module FAHDMXHT (CO, S, A, B, CI);
    output CO;
    output S;
    input A;
    input B;
    input CI;

endmodule
module FAHDUXHT (CO, S, A, B, CI);
    output CO;
    output S;
    input A;
    input B;
    input CI;

endmodule
module FAHHD1XHT (CO, S, A, B, CI);
    output CO;
    output S;
    input A;
    input B;
    input CI;

endmodule
module FAHHD2XHT (CO, S, A, B, CI);
    output CO;
    output S;
    input A;
    input B;
    input CI;

endmodule
module FAHHDLXHT (CO, S, A, B, CI);
    output CO;
    output S;
    input A;
    input B;
    input CI;

endmodule
module FAHHDMXHT (CO, S, A, B, CI);
    output CO;
    output S;
    input A;
    input B;
    input CI;

endmodule
module FFDCRHD1XHT (Q, QN, CK, D, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;

endmodule
module FFDCRHD2XHT (Q, QN, CK, D, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;

endmodule
module FFDCRHDLXHT (Q, QN, CK, D, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;

endmodule
module FFDCRHDMXHT (Q, QN, CK, D, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;

endmodule
module FFDHD1XHT (Q, QN, CK, D);
    output Q;
    output QN;
    input CK;
    input D;

endmodule
module FFDHD1XSPGHT (Q, QN, CK, D);
    output Q;
    output QN;
    input CK;
    input D;

endmodule
module FFDHD2XHT (Q, QN, CK, D);
    output Q;
    output QN;
    input CK;
    input D;

endmodule
module FFDHDLXHT (Q, QN, CK, D);
    output Q;
    output QN;
    input CK;
    input D;

endmodule
module FFDHDMXHT (Q, QN, CK, D);
    output Q;
    output QN;
    input CK;
    input D;

endmodule
module FFDHQHD1XHT (Q, CK, D);
    output Q;
    input CK;
    input D;

endmodule
module FFDHQHD2XHT (Q, CK, D);
    output Q;
    input CK;
    input D;

endmodule
module FFDHQHD3XHT (Q, CK, D);
    output Q;
    input CK;
    input D;

endmodule
module FFDHQHDMXHT (Q, CK, D);
    output Q;
    input CK;
    input D;

endmodule
module FFDNHD1XHT (Q, QN, CKN, D);
    output Q;
    output QN;
    input CKN;
    input D;

endmodule
module FFDNHD2XHT (Q, QN, CKN, D);
    output Q;
    output QN;
    input CKN;
    input D;

endmodule
module FFDNHDLXHT (Q, QN, CKN, D);
    output Q;
    output QN;
    input CKN;
    input D;

endmodule
module FFDNHDMXHT (Q, QN, CKN, D);
    output Q;
    output QN;
    input CKN;
    input D;

endmodule
module FFDNRHD1XHT (Q, QN, CKN, D, RN);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;

endmodule
module FFDNRHD2XHT (Q, QN, CKN, D, RN);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;

endmodule
module FFDNRHDLXHT (Q, QN, CKN, D, RN);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;

endmodule
module FFDNRHDMXHT (Q, QN, CKN, D, RN);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;

endmodule
module FFDNSHD1XHT (Q, QN, CKN, D, SN);
    output Q;
    output QN;
    input CKN;
    input D;
    input SN;

endmodule
module FFDNSHD2XHT (Q, QN, CKN, D, SN);
    output Q;
    output QN;
    input CKN;
    input D;
    input SN;

endmodule
module FFDNSHDLXHT (Q, QN, CKN, D, SN);
    output Q;
    output QN;
    input CKN;
    input D;
    input SN;

endmodule
module FFDNSHDMXHT (Q, QN, CKN, D, SN);
    output Q;
    output QN;
    input CKN;
    input D;
    input SN;

endmodule
module FFDNSRHD1XHT (Q, QN, CKN, D, RN, SN);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input SN;

endmodule
module FFDNSRHD2XHT (Q, QN, CKN, D, RN, SN);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input SN;

endmodule
module FFDNSRHDLXHT (Q, QN, CKN, D, RN, SN);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input SN;

endmodule
module FFDNSRHDMXHT (Q, QN, CKN, D, RN, SN);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input SN;

endmodule
module FFDQHD1XHT (Q, CK, D);
    output Q;
    input CK;
    input D;

endmodule
module FFDQHD2XHT (Q, CK, D);
    output Q;
    input CK;
    input D;

endmodule
module FFDQHDLXHT (Q, CK, D);
    output Q;
    input CK;
    input D;

endmodule
module FFDQHDMXHT (Q, CK, D);
    output Q;
    input CK;
    input D;

endmodule
module FFDQRHD1XHT (Q, CK, D, RN);
    output Q;
    input CK;
    input D;
    input RN;

endmodule
module FFDQRHD2XHT (Q, CK, D, RN);
    output Q;
    input CK;
    input D;
    input RN;

endmodule
module FFDQRHDLXHT (Q, CK, D, RN);
    output Q;
    input CK;
    input D;
    input RN;

endmodule
module FFDQRHDMXHT (Q, CK, D, RN);
    output Q;
    input CK;
    input D;
    input RN;

endmodule
module FFDQSHD1XHT (Q, CK, D, SN);
    output Q;
    input CK;
    input D;
    input SN;

endmodule
module FFDQSHD2XHT (Q, CK, D, SN);
    output Q;
    input CK;
    input D;
    input SN;

endmodule
module FFDQSHDLXHT (Q, CK, D, SN);
    output Q;
    input CK;
    input D;
    input SN;

endmodule
module FFDQSHDMXHT (Q, CK, D, SN);
    output Q;
    input CK;
    input D;
    input SN;

endmodule
module FFDQSRHD1XHT (Q, CK, D, RN, SN);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDQSRHD2XHT (Q, CK, D, RN, SN);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDQSRHDLXHT (Q, CK, D, RN, SN);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDQSRHDMXHT (Q, CK, D, RN, SN);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDRHD1XHT (Q, QN, CK, D, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;

endmodule
module FFDRHD2XHT (Q, QN, CK, D, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;

endmodule
module FFDRHDLXHT (Q, QN, CK, D, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;

endmodule
module FFDRHDMXHT (Q, QN, CK, D, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;

endmodule
module FFDRHQHD1XHT (Q, CK, D, RN);
    output Q;
    input CK;
    input D;
    input RN;

endmodule
module FFDRHQHD2XHT (Q, CK, D, RN);
    output Q;
    input CK;
    input D;
    input RN;

endmodule
module FFDRHQHD3XHT (Q, CK, D, RN);
    output Q;
    input CK;
    input D;
    input RN;

endmodule
module FFDRHQHDMXHT (Q, CK, D, RN);
    output Q;
    input CK;
    input D;
    input RN;

endmodule
module FFDSHD1XHT (Q, QN, CK, D, SN);
    output Q;
    output QN;
    input CK;
    input D;
    input SN;

endmodule
module FFDSHD2XHT (Q, QN, CK, D, SN);
    output Q;
    output QN;
    input CK;
    input D;
    input SN;

endmodule
module FFDSHDLXHT (Q, QN, CK, D, SN);
    output Q;
    output QN;
    input CK;
    input D;
    input SN;

endmodule
module FFDSHDMXHT (Q, QN, CK, D, SN);
    output Q;
    output QN;
    input CK;
    input D;
    input SN;

endmodule
module FFDSHQHD1XHT (Q, CK, D, SN);
    output Q;
    input CK;
    input D;
    input SN;

endmodule
module FFDSHQHD2XHT (Q, CK, D, SN);
    output Q;
    input CK;
    input D;
    input SN;

endmodule
module FFDSHQHD3XHT (Q, CK, D, SN);
    output Q;
    input CK;
    input D;
    input SN;

endmodule
module FFDSHQHDMXHT (Q, CK, D, SN);
    output Q;
    input CK;
    input D;
    input SN;

endmodule
module FFDSRHD1XHT (Q, QN, CK, D, RN, SN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDSRHD2XHT (Q, QN, CK, D, RN, SN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDSRHDLXHT (Q, QN, CK, D, RN, SN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDSRHDMXHT (Q, QN, CK, D, RN, SN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDSRHQHD1XHT (Q, CK, D, RN, SN);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDSRHQHD2XHT (Q, CK, D, RN, SN);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDSRHQHD3XHT (Q, CK, D, RN, SN);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDSRHQHDMXHT (Q, CK, D, RN, SN);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFEDCRHD1XHT (Q, QN, CK, D, E, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input RN;

endmodule
module FFEDCRHD2XHT (Q, QN, CK, D, E, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input RN;

endmodule
module FFEDCRHDLXHT (Q, QN, CK, D, E, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input RN;

endmodule
module FFEDCRHDMXHT (Q, QN, CK, D, E, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input RN;

endmodule
module FFEDHD1XHT (Q, QN, CK, D, E);
    output Q;
    output QN;
    input CK;
    input D;
    input E;

endmodule
module FFEDHD2XHT (Q, QN, CK, D, E);
    output Q;
    output QN;
    input CK;
    input D;
    input E;

endmodule
module FFEDHDLXHT (Q, QN, CK, D, E);
    output Q;
    output QN;
    input CK;
    input D;
    input E;

endmodule
module FFEDHDMXHT (Q, QN, CK, D, E);
    output Q;
    output QN;
    input CK;
    input D;
    input E;

endmodule
module FFEDHQHD1XHT (Q, CK, D, E);
    output Q;
    input CK;
    input D;
    input E;

endmodule
module FFEDHQHD2XHT (Q, CK, D, E);
    output Q;
    input CK;
    input D;
    input E;

endmodule
module FFEDHQHD3XHT (Q, CK, D, E);
    output Q;
    input CK;
    input D;
    input E;

endmodule
module FFEDHQHDMXHT (Q, CK, D, E);
    output Q;
    input CK;
    input D;
    input E;

endmodule
module FFEDQHD1XHT (Q, CK, D, E);
    output Q;
    input CK;
    input D;
    input E;

endmodule
module FFEDQHD2XHT (Q, CK, D, E);
    output Q;
    input CK;
    input D;
    input E;

endmodule
module FFEDQHDLXHT (Q, CK, D, E);
    output Q;
    input CK;
    input D;
    input E;

endmodule
module FFEDQHDMXHT (Q, CK, D, E);
    output Q;
    input CK;
    input D;
    input E;

endmodule
module FFSDCRHD1XHT (Q, QN, CK, D, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDCRHD2XHT (Q, QN, CK, D, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDCRHDLXHT (Q, QN, CK, D, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDCRHDMXHT (Q, QN, CK, D, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDHD1XHT (Q, QN, CK, D, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDHD1XSPGHT (Q, QN, CK, D, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDHD2XHT (Q, QN, CK, D, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDHDLXHT (Q, QN, CK, D, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDHDMXHT (Q, QN, CK, D, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDHQHD1XHT (Q, CK, D, TE, TI);
    output Q;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDHQHD2XHT (Q, CK, D, TE, TI);
    output Q;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDHQHD3XHT (Q, CK, D, TE, TI);
    output Q;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDHQHDMXHT (Q, CK, D, TE, TI);
    output Q;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDNHD1XHT (Q, QN, CKN, D, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input TE;
    input TI;

endmodule
module FFSDNHD2XHT (Q, QN, CKN, D, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input TE;
    input TI;

endmodule
module FFSDNHDLXHT (Q, QN, CKN, D, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input TE;
    input TI;

endmodule
module FFSDNHDMXHT (Q, QN, CKN, D, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input TE;
    input TI;

endmodule
module FFSDNRHD1XHT (Q, QN, CKN, D, RN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDNRHD2XHT (Q, QN, CKN, D, RN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDNRHDLXHT (Q, QN, CKN, D, RN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDNRHDMXHT (Q, QN, CKN, D, RN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDNSHD1XHT (Q, QN, CKN, D, SN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDNSHD2XHT (Q, QN, CKN, D, SN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDNSHDLXHT (Q, QN, CKN, D, SN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDNSHDMXHT (Q, QN, CKN, D, SN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDNSRHD1XHT (Q, QN, CKN, D, RN, SN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDNSRHD2XHT (Q, QN, CKN, D, RN, SN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDNSRHDLXHT (Q, QN, CKN, D, RN, SN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDNSRHDMXHT (Q, QN, CKN, D, RN, SN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDQHD1XHT (Q, CK, D, TE, TI);
    output Q;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDQHD2XHT (Q, CK, D, TE, TI);
    output Q;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDQHDLXHT (Q, CK, D, TE, TI);
    output Q;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDQHDMXHT (Q, CK, D, TE, TI);
    output Q;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDQRHD1XHT (Q, CK, D, RN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDQRHD2XHT (Q, CK, D, RN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDQRHDLXHT (Q, CK, D, RN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDQRHDMXHT (Q, CK, D, RN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDQSHD1XHT (Q, CK, D, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDQSHD2XHT (Q, CK, D, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDQSHDLXHT (Q, CK, D, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDQSHDMXHT (Q, CK, D, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDQSRHD1XHT (Q, CK, D, RN, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDQSRHD2XHT (Q, CK, D, RN, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDQSRHDLXHT (Q, CK, D, RN, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDQSRHDMXHT (Q, CK, D, RN, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDRHD1XHT (Q, QN, CK, D, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDRHD2XHT (Q, QN, CK, D, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDRHDLXHT (Q, QN, CK, D, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDRHDMXHT (Q, QN, CK, D, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDRHQHD1XHT (Q, CK, D, RN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDRHQHD2XHT (Q, CK, D, RN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDRHQHD3XHT (Q, CK, D, RN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDRHQHDMXHT (Q, CK, D, RN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDSHD1XHT (Q, QN, CK, D, SN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSHD2XHT (Q, QN, CK, D, SN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSHDLXHT (Q, QN, CK, D, SN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSHDMXHT (Q, QN, CK, D, SN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSHQHD1XHT (Q, CK, D, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSHQHD2XHT (Q, CK, D, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSHQHD3XHT (Q, CK, D, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSHQHDMXHT (Q, CK, D, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSRHD1XHT (Q, QN, CK, D, RN, SN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSRHD2XHT (Q, QN, CK, D, RN, SN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSRHDLXHT (Q, QN, CK, D, RN, SN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSRHDMXHT (Q, QN, CK, D, RN, SN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSRHQHD1XHT (Q, CK, D, RN, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSRHQHD2XHT (Q, CK, D, RN, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSRHQHD3XHT (Q, CK, D, RN, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSRHQHDMXHT (Q, CK, D, RN, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSEDCRHD1XHT (Q, QN, CK, D, E, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input RN;
    input TE;
    input TI;

endmodule
module FFSEDCRHD2XHT (Q, QN, CK, D, E, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input RN;
    input TE;
    input TI;

endmodule
module FFSEDCRHDLXHT (Q, QN, CK, D, E, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input RN;
    input TE;
    input TI;

endmodule
module FFSEDCRHDMXHT (Q, QN, CK, D, E, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input RN;
    input TE;
    input TI;

endmodule
module FFSEDHD1XHT (Q, QN, CK, D, E, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDHD2XHT (Q, QN, CK, D, E, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDHDLXHT (Q, QN, CK, D, E, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDHDMXHT (Q, QN, CK, D, E, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDHQHD1XHT (Q, CK, D, E, TE, TI);
    output Q;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDHQHD2XHT (Q, CK, D, E, TE, TI);
    output Q;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDHQHD3XHT (Q, CK, D, E, TE, TI);
    output Q;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDHQHDMXHT (Q, CK, D, E, TE, TI);
    output Q;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDQHD1XHT (Q, CK, D, E, TE, TI);
    output Q;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDQHD2XHT (Q, CK, D, E, TE, TI);
    output Q;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDQHDLXHT (Q, CK, D, E, TE, TI);
    output Q;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDQHDMXHT (Q, CK, D, E, TE, TI);
    output Q;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FILLER16HD ;

endmodule
module FILLER1HD ;

endmodule
module FILLER2HD ;

endmodule
module FILLER32HD ;

endmodule
module FILLER3HD ;

endmodule
module FILLER4HD ;

endmodule
module FILLER64HD ;

endmodule
module FILLER6HD ;

endmodule
module FILLER8HD ;

endmodule
module FILLERC16HD ;

endmodule
module FILLERC1HD ;

endmodule
module FILLERC2HD ;

endmodule
module FILLERC32HD ;

endmodule
module FILLERC3HD ;

endmodule
module FILLERC4HD ;

endmodule
module FILLERC64HD ;

endmodule
module FILLERC6HD ;

endmodule
module FILLERC8HD ;

endmodule
module HAHD1XHT (CO, S, A, B);
    output CO;
    output S;
    input A;
    input B;

endmodule
module HAHD2XHT (CO, S, A, B);
    output CO;
    output S;
    input A;
    input B;

endmodule
module HAHDLXHT (CO, S, A, B);
    output CO;
    output S;
    input A;
    input B;

endmodule
module HAHDMXHT (CO, S, A, B);
    output CO;
    output S;
    input A;
    input B;

endmodule
module HOLDHDHT (Z);
    inout Z;

endmodule
module INVCLKHD10XHT (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD12XHT (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD14XHT (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD16XHT (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD1XHT (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD20XHT (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD2XHT (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD30XHT (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD3XHT (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD40XHT (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD4XHT (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD5XHT (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD6XHT (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD7XHT (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD80XHT (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD8XHT (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHDLXHT (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHDMXHT (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHDUXHT (Z, A);
    output Z;
    input A;

endmodule
module INVHD12XHT (Z, A);
    output Z;
    input A;

endmodule
module INVHD16XHT (Z, A);
    output Z;
    input A;

endmodule
module INVHD1XHT (Z, A);
    output Z;
    input A;

endmodule
module INVHD1XSPGHT (Z, A);
    output Z;
    input A;

endmodule
module INVHD20XHT (Z, A);
    output Z;
    input A;

endmodule
module INVHD2XHT (Z, A);
    output Z;
    input A;

endmodule
module INVHD3XHT (Z, A);
    output Z;
    input A;

endmodule
module INVHD4XHT (Z, A);
    output Z;
    input A;

endmodule
module INVHD5XHT (Z, A);
    output Z;
    input A;

endmodule
module INVHD6XHT (Z, A);
    output Z;
    input A;

endmodule
module INVHD7XHT (Z, A);
    output Z;
    input A;

endmodule
module INVHD8XHT (Z, A);
    output Z;
    input A;

endmodule
module INVHDLXHT (Z, A);
    output Z;
    input A;

endmodule
module INVHDMXHT (Z, A);
    output Z;
    input A;

endmodule
module INVHDPXHT (Z, A);
    output Z;
    input A;

endmodule
module INVHDUXHT (Z, A);
    output Z;
    input A;

endmodule
module INVODHD8XHT (Z0, Z1, Z2, Z3, Z4, Z5, Z6, Z7, A);
    output Z0;
    output Z1;
    output Z2;
    output Z3;
    output Z4;
    output Z5;
    output Z6;
    output Z7;
    input A;

endmodule
module INVTSHD12XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD16XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD1XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD20XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD2XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD3XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD4XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD5XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD6XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD7XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD8XHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHDLXHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHDMXHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHDUXHT (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module LATHD1XHT (Q, QN, D, G);
    output Q;
    output QN;
    input D;
    input G;

endmodule
module LATHD1XSPGHT (Q, QN, D, G);
    output Q;
    output QN;
    input D;
    input G;

endmodule
module LATHD2XHT (Q, QN, D, G);
    output Q;
    output QN;
    input D;
    input G;

endmodule
module LATHDLXHT (Q, QN, D, G);
    output Q;
    output QN;
    input D;
    input G;

endmodule
module LATHDMXHT (Q, QN, D, G);
    output Q;
    output QN;
    input D;
    input G;

endmodule
module LATNHD1XHT (Q, QN, D, GN);
    output Q;
    output QN;
    input D;
    input GN;

endmodule
module LATNHD2XHT (Q, QN, D, GN);
    output Q;
    output QN;
    input D;
    input GN;

endmodule
module LATNHDLXHT (Q, QN, D, GN);
    output Q;
    output QN;
    input D;
    input GN;

endmodule
module LATNHDMXHT (Q, QN, D, GN);
    output Q;
    output QN;
    input D;
    input GN;

endmodule
module LATNRHD1XHT (Q, QN, D, GN, RN);
    output Q;
    output QN;
    input D;
    input GN;
    input RN;

endmodule
module LATNRHD2XHT (Q, QN, D, GN, RN);
    output Q;
    output QN;
    input D;
    input GN;
    input RN;

endmodule
module LATNRHDLXHT (Q, QN, D, GN, RN);
    output Q;
    output QN;
    input D;
    input GN;
    input RN;

endmodule
module LATNRHDMXHT (Q, QN, D, GN, RN);
    output Q;
    output QN;
    input D;
    input GN;
    input RN;

endmodule
module LATNSHD1XHT (Q, QN, D, GN, SN);
    output Q;
    output QN;
    input D;
    input GN;
    input SN;

endmodule
module LATNSHD2XHT (Q, QN, D, GN, SN);
    output Q;
    output QN;
    input D;
    input GN;
    input SN;

endmodule
module LATNSHDLXHT (Q, QN, D, GN, SN);
    output Q;
    output QN;
    input D;
    input GN;
    input SN;

endmodule
module LATNSHDMXHT (Q, QN, D, GN, SN);
    output Q;
    output QN;
    input D;
    input GN;
    input SN;

endmodule
module LATNSRHD1XHT (Q, QN, D, GN, RN, SN);
    output Q;
    output QN;
    input D;
    input GN;
    input RN;
    input SN;

endmodule
module LATNSRHD2XHT (Q, QN, D, GN, RN, SN);
    output Q;
    output QN;
    input D;
    input GN;
    input RN;
    input SN;

endmodule
module LATNSRHDLXHT (Q, QN, D, GN, RN, SN);
    output Q;
    output QN;
    input D;
    input GN;
    input RN;
    input SN;

endmodule
module LATNSRHDMXHT (Q, QN, D, GN, RN, SN);
    output Q;
    output QN;
    input D;
    input GN;
    input RN;
    input SN;

endmodule
module LATRHD1XHT (Q, QN, D, G, RN);
    output Q;
    output QN;
    input D;
    input G;
    input RN;

endmodule
module LATRHD2XHT (Q, QN, D, G, RN);
    output Q;
    output QN;
    input D;
    input G;
    input RN;

endmodule
module LATRHDLXHT (Q, QN, D, G, RN);
    output Q;
    output QN;
    input D;
    input G;
    input RN;

endmodule
module LATRHDMXHT (Q, QN, D, G, RN);
    output Q;
    output QN;
    input D;
    input G;
    input RN;

endmodule
module LATSHD1XHT (Q, QN, D, G, SN);
    output Q;
    output QN;
    input D;
    input G;
    input SN;

endmodule
module LATSHD2XHT (Q, QN, D, G, SN);
    output Q;
    output QN;
    input D;
    input G;
    input SN;

endmodule
module LATSHDLXHT (Q, QN, D, G, SN);
    output Q;
    output QN;
    input D;
    input G;
    input SN;

endmodule
module LATSHDMXHT (Q, QN, D, G, SN);
    output Q;
    output QN;
    input D;
    input G;
    input SN;

endmodule
module LATSRHD1XHT (Q, QN, D, G, RN, SN);
    output Q;
    output QN;
    input D;
    input G;
    input RN;
    input SN;

endmodule
module LATSRHD2XHT (Q, QN, D, G, RN, SN);
    output Q;
    output QN;
    input D;
    input G;
    input RN;
    input SN;

endmodule
module LATSRHDLXHT (Q, QN, D, G, RN, SN);
    output Q;
    output QN;
    input D;
    input G;
    input RN;
    input SN;

endmodule
module LATSRHDMXHT (Q, QN, D, G, RN, SN);
    output Q;
    output QN;
    input D;
    input G;
    input RN;
    input SN;

endmodule
module LATTSHD1XHT (Q, D, E, G);
    output Q;
    input D;
    input E;
    input G;

endmodule
module LATTSHD2XHT (Q, D, E, G);
    output Q;
    input D;
    input E;
    input G;

endmodule
module LATTSHDLXHT (Q, D, E, G);
    output Q;
    input D;
    input E;
    input G;

endmodule
module LATTSHDMXHT (Q, D, E, G);
    output Q;
    input D;
    input E;
    input G;

endmodule
module MUX2CLKHD1XHT (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2CLKHD2XHT (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2CLKHD3XHT (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2CLKHD4XHT (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2HD1XHT (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2HD1XSPGHT (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2HD2XHT (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2HD3XHT (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2HDLXHT (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2HDMXHT (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2HDUXHT (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX4HD1XHT (Z, A, B, C, D, S0, S1);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input S0;
    input S1;

endmodule
module MUX4HD2XHT (Z, A, B, C, D, S0, S1);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input S0;
    input S1;

endmodule
module MUX4HDLXHT (Z, A, B, C, D, S0, S1);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input S0;
    input S1;

endmodule
module MUX4HDMXHT (Z, A, B, C, D, S0, S1);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input S0;
    input S1;

endmodule
module MUXI2HD1XHT (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUXI2HD2XHT (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUXI2HD3XHT (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUXI2HDLXHT (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUXI2HDMXHT (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUXI4HD1XHT (Z, A, B, C, D, S0, S1);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input S0;
    input S1;

endmodule
module MUXI4HD2XHT (Z, A, B, C, D, S0, S1);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input S0;
    input S1;

endmodule
module MUXI4HDLXHT (Z, A, B, C, D, S0, S1);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input S0;
    input S1;

endmodule
module MUXI4HDMXHT (Z, A, B, C, D, S0, S1);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input S0;
    input S1;

endmodule
module NAND2B1HD1XHT (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NAND2B1HD2XHT (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NAND2B1HDLXHT (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NAND2B1HDMXHT (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NAND2B1HDUXHT (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NAND2HD1XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NAND2HD1XSPGHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NAND2HD2XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NAND2HD2XSPGHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NAND2HD3XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NAND2HDLXHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NAND2HDMXHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NAND2HDUXHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NAND2ODHDHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NAND3B1HD1XHT (Z, AN, B, C);
    output Z;
    input AN;
    input B;
    input C;

endmodule
module NAND3B1HD2XHT (Z, AN, B, C);
    output Z;
    input AN;
    input B;
    input C;

endmodule
module NAND3B1HDLXHT (Z, AN, B, C);
    output Z;
    input AN;
    input B;
    input C;

endmodule
module NAND3B1HDMXHT (Z, AN, B, C);
    output Z;
    input AN;
    input B;
    input C;

endmodule
module NAND3HD1XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NAND3HD2XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NAND3HD3XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NAND3HDLXHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NAND3HDMXHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NAND3ODHDHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NAND4B1HD1XHT (Z, AN, B, C, D);
    output Z;
    input AN;
    input B;
    input C;
    input D;

endmodule
module NAND4B1HD2XHT (Z, AN, B, C, D);
    output Z;
    input AN;
    input B;
    input C;
    input D;

endmodule
module NAND4B1HDLXHT (Z, AN, B, C, D);
    output Z;
    input AN;
    input B;
    input C;
    input D;

endmodule
module NAND4B1HDMXHT (Z, AN, B, C, D);
    output Z;
    input AN;
    input B;
    input C;
    input D;

endmodule
module NAND4B2HD1XHT (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module NAND4B2HD2XHT (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module NAND4B2HDLXHT (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module NAND4B2HDMXHT (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module NAND4HD1XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module NAND4HD2XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module NAND4HD3XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module NAND4HDLXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module NAND4HDMXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module NOR2B1HD1XHT (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NOR2B1HD2XHT (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NOR2B1HDLXHT (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NOR2B1HDMXHT (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NOR2B1HDUXHT (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NOR2HD1XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NOR2HD1XSPGHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NOR2HD2XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NOR2HD2XSPGHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NOR2HD3XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NOR2HDLXHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NOR2HDMXHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NOR2HDUXHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NOR3B1HD1XHT (Z, AN, B, C);
    output Z;
    input AN;
    input B;
    input C;

endmodule
module NOR3B1HD2XHT (Z, AN, B, C);
    output Z;
    input AN;
    input B;
    input C;

endmodule
module NOR3B1HDLXHT (Z, AN, B, C);
    output Z;
    input AN;
    input B;
    input C;

endmodule
module NOR3B1HDMXHT (Z, AN, B, C);
    output Z;
    input AN;
    input B;
    input C;

endmodule
module NOR3HD1XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NOR3HD2XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NOR3HD3XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NOR3HDLXHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NOR3HDMXHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NOR4B1HD1XHT (Z, AN, B, C, D);
    output Z;
    input AN;
    input B;
    input C;
    input D;

endmodule
module NOR4B1HD2XHT (Z, AN, B, C, D);
    output Z;
    input AN;
    input B;
    input C;
    input D;

endmodule
module NOR4B1HDLXHT (Z, AN, B, C, D);
    output Z;
    input AN;
    input B;
    input C;
    input D;

endmodule
module NOR4B1HDMXHT (Z, AN, B, C, D);
    output Z;
    input AN;
    input B;
    input C;
    input D;

endmodule
module NOR4B2HD1XHT (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module NOR4B2HD2XHT (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module NOR4B2HDLXHT (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module NOR4B2HDMXHT (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module NOR4HD1XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module NOR4HD2XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module NOR4HD3XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module NOR4HDLXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module NOR4HDMXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI211HD1XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI211HD2XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI211HDLXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI211HDMXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI21B2HD1XHT (Z, AN, BN, C);
    output Z;
    input AN;
    input BN;
    input C;

endmodule
module OAI21B2HD2XHT (Z, AN, BN, C);
    output Z;
    input AN;
    input BN;
    input C;

endmodule
module OAI21B2HDLXHT (Z, AN, BN, C);
    output Z;
    input AN;
    input BN;
    input C;

endmodule
module OAI21B2HDMXHT (Z, AN, BN, C);
    output Z;
    input AN;
    input BN;
    input C;

endmodule
module OAI21HD1XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module OAI21HD2XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module OAI21HDLXHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module OAI21HDMXHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module OAI21HDUXHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module OAI221HD1XHT (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module OAI221HD2XHT (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module OAI221HDLXHT (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module OAI221HDMXHT (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module OAI222HD1XHT (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module OAI222HD2XHT (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module OAI222HDLXHT (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module OAI222HDMXHT (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module OAI22B2HD1XHT (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module OAI22B2HD2XHT (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module OAI22B2HDLXHT (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module OAI22B2HDMXHT (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module OAI22HD1XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI22HD2XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI22HDLXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI22HDMXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI22HDUXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI31HD1XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI31HD2XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI31HDLXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI31HDMXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI32HD1XHT (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module OAI32HD2XHT (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module OAI32HDLXHT (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module OAI32HDMXHT (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module OAI33HD1XHT (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module OAI33HD2XHT (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module OAI33HDLXHT (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module OAI33HDMXHT (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module OR2HD1XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module OR2HD1XSPGHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module OR2HD2XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module OR2HD2XSPGHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module OR2HDLXHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module OR2HDMXHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module OR2HDUXHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module OR2ODHDHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module OR3HD1XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module OR3HD2XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module OR3HDLXHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module OR3HDMXHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module OR4HD1XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OR4HD2XHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OR4HDLXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OR4HDMXHT (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module PULLDHDHT (Z, EN);
    output Z;
    input EN;

endmodule
module PULLUHDHT (Z, E);
    output Z;
    input E;

endmodule
module RSLATHD1XHT (Q, QN, R, S);
    output Q;
    output QN;
    input R;
    input S;

endmodule
module RSLATHD2XHT (Q, QN, R, S);
    output Q;
    output QN;
    input R;
    input S;

endmodule
module RSLATHDLXHT (Q, QN, R, S);
    output Q;
    output QN;
    input R;
    input S;

endmodule
module RSLATHDMXHT (Q, QN, R, S);
    output Q;
    output QN;
    input R;
    input S;

endmodule
module RSLATNHD1XHT (Q, QN, RN, SN);
    output Q;
    output QN;
    input RN;
    input SN;

endmodule
module RSLATNHD2XHT (Q, QN, RN, SN);
    output Q;
    output QN;
    input RN;
    input SN;

endmodule
module RSLATNHDLXHT (Q, QN, RN, SN);
    output Q;
    output QN;
    input RN;
    input SN;

endmodule
module RSLATNHDMXHT (Q, QN, RN, SN);
    output Q;
    output QN;
    input RN;
    input SN;

endmodule
module TIEHHDHT (Z);
    output Z;

endmodule
module TIELHDHT (Z);
    output Z;

endmodule
module XNOR2HD1XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XNOR2HD2XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XNOR2HD3XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XNOR2HDLXHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XNOR2HDMXHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XNOR3HD1XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module XNOR3HD2XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module XNOR3HD3XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module XNOR3HDLXHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module XNOR3HDMXHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module XOR2CLKHD1XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XOR2CLKHD2XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XOR2CLKHD3XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XOR2CLKHD4XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XOR2HD1XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XOR2HD2XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XOR2HD3XHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XOR2HDLXHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XOR2HDMXHT (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XOR3HD1XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module XOR3HD2XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module XOR3HD3XHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module XOR3HDLXHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module XOR3HDMXHT (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
