module PLBIAR (AI, P);
    inout AI;
    inout P;

endmodule
module PLBIA (P);
    inout P;

endmodule
module PLBI16F (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PLBI16N (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PLBI16S (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PLBI24F (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PLBI24N (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PLBI24S (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PLBI2F (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PLBI2N (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PLBI2S (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PLBI4F (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PLBI4N (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PLBI4S (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PLBI8F (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PLBI8N (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PLBI8S (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PLOSCR14M (CK, XTALOUT, EI, EO, XTALIN);
    output CK;
    output XTALOUT;
    input EI;
    input EO;
    input XTALIN;

endmodule
module PLOSC14M (CK, XTALOUT, EI, EO, XTALIN);
    output CK;
    output XTALOUT;
    input EI;
    input EO;
    input XTALIN;

endmodule
module PLVDDC (vdd);
    inout vdd;

endmodule
module PLVDDH (VDDH);
    inout VDDH;

endmodule
module PLVDDO (VDDO);
    inout VDDO;

endmodule
module PLVSSC (gnd);
    inout gnd;

endmodule
module PLVSSH (VSSH);
    inout VSSH;

endmodule
module PLVSSO (VSSO);
    inout VSSO;

endmodule
module PSBIAR (AI, P);
    inout AI;
    inout P;

endmodule
module PSBIA (P);
    inout P;

endmodule
module PSBI16F (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PSBI16N (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PSBI16S (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PSBI24F (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PSBI24N (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PSBI24S (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PSBI2F (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PSBI2N (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PSBI2S (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PSBI4F (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PSBI4N (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PSBI4S (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PSBI8F (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PSBI8N (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PSBI8S (D, P, A, CONOF, NEN, PD, PEN, PU, SONOF);
    output D;
    inout P;
    input A;
    input CONOF;
    input NEN;
    input PD;
    input PEN;
    input PU;
    input SONOF;

endmodule
module PSOSCR14M (CK, XTALOUT, EI, EO, XTALIN);
    output CK;
    output XTALOUT;
    input EI;
    input EO;
    input XTALIN;

endmodule
module PSOSC14M (CK, XTALOUT, EI, EO, XTALIN);
    output CK;
    output XTALOUT;
    input EI;
    input EO;
    input XTALIN;

endmodule
module PSVDDC (vdd);
    inout vdd;

endmodule
module PSVDDH (VDDH);
    inout VDDH;

endmodule
module PSVDDO (VDDO);
    inout VDDO;

endmodule
module PSVSSC (gnd);
    inout gnd;

endmodule
module PSVSSH (VSSH);
    inout VSSH;

endmodule
module PSVSSO (VSSO);
    inout VSSO;

endmodule
