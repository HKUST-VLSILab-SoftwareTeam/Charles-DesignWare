module AND2CLKHD1X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2CLKHD2X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2CLKHD3X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2CLKHD4X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2HD1X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2HD1XSPG (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2HD2X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2HD2XSPG (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2HDLX (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2HDMX (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND2HDUX (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module AND3HD1X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module AND3HD2X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module AND3HDLX (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module AND3HDMX (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module AND4HD1X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AND4HD2X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AND4HDLX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AND4HDMX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module ANTFIXHD (Z);
    output Z;

endmodule
module AOI211HD1X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI211HD2X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI211HDLX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI211HDMX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI21B2HD1X (Z, AN, BN, C);
    output Z;
    input AN;
    input BN;
    input C;

endmodule
module AOI21B2HD2X (Z, AN, BN, C);
    output Z;
    input AN;
    input BN;
    input C;

endmodule
module AOI21B2HDLX (Z, AN, BN, C);
    output Z;
    input AN;
    input BN;
    input C;

endmodule
module AOI21B2HDMX (Z, AN, BN, C);
    output Z;
    input AN;
    input BN;
    input C;

endmodule
module AOI21HD1X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module AOI21HD2X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module AOI21HDLX (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module AOI21HDMX (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module AOI21HDUX (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module AOI221HD1X (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module AOI221HD2X (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module AOI221HDLX (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module AOI221HDMX (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module AOI222HD1X (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module AOI222HD2X (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module AOI222HDLX (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module AOI222HDMX (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module AOI22B2HD1X (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module AOI22B2HD2X (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module AOI22B2HDLX (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module AOI22B2HDMX (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module AOI22HD1X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI22HD2X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI22HDLX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI22HDMX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI22HDUX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI31HD1X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI31HD2X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI31HDLX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI31HDMX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module AOI32HD1X (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module AOI32HD2X (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module AOI32HDLX (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module AOI32HDMX (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module AOI33HD1X (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module AOI33HD2X (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module AOI33HDLX (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module AOI33HDMX (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module BUFCLKHD10X (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD12X (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD14X (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD16X (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD1X (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD20X (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD2X (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD30X (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD3X (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD40X (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD4X (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD5X (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD6X (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD7X (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD80X (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHD8X (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHDLX (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHDMX (Z, A);
    output Z;
    input A;

endmodule
module BUFCLKHDUX (Z, A);
    output Z;
    input A;

endmodule
module BUFHD12X (Z, A);
    output Z;
    input A;

endmodule
module BUFHD16X (Z, A);
    output Z;
    input A;

endmodule
module BUFHD1X (Z, A);
    output Z;
    input A;

endmodule
module BUFHD20X (Z, A);
    output Z;
    input A;

endmodule
module BUFHD2X (Z, A);
    output Z;
    input A;

endmodule
module BUFHD3X (Z, A);
    output Z;
    input A;

endmodule
module BUFHD4X (Z, A);
    output Z;
    input A;

endmodule
module BUFHD5X (Z, A);
    output Z;
    input A;

endmodule
module BUFHD6X (Z, A);
    output Z;
    input A;

endmodule
module BUFHD7X (Z, A);
    output Z;
    input A;

endmodule
module BUFHD8X (Z, A);
    output Z;
    input A;

endmodule
module BUFHD8XSPG (Z, A);
    output Z;
    input A;

endmodule
module BUFHDLX (Z, A);
    output Z;
    input A;

endmodule
module BUFHDMX (Z, A);
    output Z;
    input A;

endmodule
module BUFHDUX (Z, A);
    output Z;
    input A;

endmodule
module BUFTSHD12X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD16X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD1X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD20X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD2X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD3X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD4X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD5X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD6X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD7X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHD8X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHDLX (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHDMX (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module BUFTSHDUX (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module DEL1HD1X (Z, A);
    output Z;
    input A;

endmodule
module DEL1HDMX (Z, A);
    output Z;
    input A;

endmodule
module DEL1HDMXSPG (Z, A);
    output Z;
    input A;

endmodule
module DEL2HD1X (Z, A);
    output Z;
    input A;

endmodule
module DEL2HDMX (Z, A);
    output Z;
    input A;

endmodule
module DEL2HDMXSPG (Z, A);
    output Z;
    input A;

endmodule
module DEL3HD1X (Z, A);
    output Z;
    input A;

endmodule
module DEL3HDMX (Z, A);
    output Z;
    input A;

endmodule
module DEL4HD1X (Z, A);
    output Z;
    input A;

endmodule
module DEL4HDMX (Z, A);
    output Z;
    input A;

endmodule
module DEL4HDMXSPG (Z, A);
    output Z;
    input A;

endmodule
module FAHD1X (CO, S, A, B, CI);
    output CO;
    output S;
    input A;
    input B;
    input CI;

endmodule
module FAHD2X (CO, S, A, B, CI);
    output CO;
    output S;
    input A;
    input B;
    input CI;

endmodule
module FAHDLX (CO, S, A, B, CI);
    output CO;
    output S;
    input A;
    input B;
    input CI;

endmodule
module FAHDMX (CO, S, A, B, CI);
    output CO;
    output S;
    input A;
    input B;
    input CI;

endmodule
module FAHDUX (CO, S, A, B, CI);
    output CO;
    output S;
    input A;
    input B;
    input CI;

endmodule
module FAHHD1X (CO, S, A, B, CI);
    output CO;
    output S;
    input A;
    input B;
    input CI;

endmodule
module FAHHD2X (CO, S, A, B, CI);
    output CO;
    output S;
    input A;
    input B;
    input CI;

endmodule
module FAHHDLX (CO, S, A, B, CI);
    output CO;
    output S;
    input A;
    input B;
    input CI;

endmodule
module FAHHDMX (CO, S, A, B, CI);
    output CO;
    output S;
    input A;
    input B;
    input CI;

endmodule
module FFDCRHD1X (Q, QN, CK, D, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;

endmodule
module FFDCRHD2X (Q, QN, CK, D, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;

endmodule
module FFDCRHDLX (Q, QN, CK, D, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;

endmodule
module FFDCRHDMX (Q, QN, CK, D, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;

endmodule
module FFDHD1X (Q, QN, CK, D);
    output Q;
    output QN;
    input CK;
    input D;

endmodule
module FFDHD1XSPG (Q, QN, CK, D);
    output Q;
    output QN;
    input CK;
    input D;

endmodule
module FFDHD2X (Q, QN, CK, D);
    output Q;
    output QN;
    input CK;
    input D;

endmodule
module FFDHDLX (Q, QN, CK, D);
    output Q;
    output QN;
    input CK;
    input D;

endmodule
module FFDHDMX (Q, QN, CK, D);
    output Q;
    output QN;
    input CK;
    input D;

endmodule
module FFDHQHD1X (Q, CK, D);
    output Q;
    input CK;
    input D;

endmodule
module FFDHQHD2X (Q, CK, D);
    output Q;
    input CK;
    input D;

endmodule
module FFDHQHD3X (Q, CK, D);
    output Q;
    input CK;
    input D;

endmodule
module FFDHQHDMX (Q, CK, D);
    output Q;
    input CK;
    input D;

endmodule
module FFDNHD1X (Q, QN, CKN, D);
    output Q;
    output QN;
    input CKN;
    input D;

endmodule
module FFDNHD2X (Q, QN, CKN, D);
    output Q;
    output QN;
    input CKN;
    input D;

endmodule
module FFDNHDLX (Q, QN, CKN, D);
    output Q;
    output QN;
    input CKN;
    input D;

endmodule
module FFDNHDMX (Q, QN, CKN, D);
    output Q;
    output QN;
    input CKN;
    input D;

endmodule
module FFDNRHD1X (Q, QN, CKN, D, RN);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;

endmodule
module FFDNRHD2X (Q, QN, CKN, D, RN);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;

endmodule
module FFDNRHDLX (Q, QN, CKN, D, RN);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;

endmodule
module FFDNRHDMX (Q, QN, CKN, D, RN);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;

endmodule
module FFDNSHD1X (Q, QN, CKN, D, SN);
    output Q;
    output QN;
    input CKN;
    input D;
    input SN;

endmodule
module FFDNSHD2X (Q, QN, CKN, D, SN);
    output Q;
    output QN;
    input CKN;
    input D;
    input SN;

endmodule
module FFDNSHDLX (Q, QN, CKN, D, SN);
    output Q;
    output QN;
    input CKN;
    input D;
    input SN;

endmodule
module FFDNSHDMX (Q, QN, CKN, D, SN);
    output Q;
    output QN;
    input CKN;
    input D;
    input SN;

endmodule
module FFDNSRHD1X (Q, QN, CKN, D, RN, SN);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input SN;

endmodule
module FFDNSRHD2X (Q, QN, CKN, D, RN, SN);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input SN;

endmodule
module FFDNSRHDLX (Q, QN, CKN, D, RN, SN);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input SN;

endmodule
module FFDNSRHDMX (Q, QN, CKN, D, RN, SN);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input SN;

endmodule
module FFDQHD1X (Q, CK, D);
    output Q;
    input CK;
    input D;

endmodule
module FFDQHD2X (Q, CK, D);
    output Q;
    input CK;
    input D;

endmodule
module FFDQHDLX (Q, CK, D);
    output Q;
    input CK;
    input D;

endmodule
module FFDQHDMX (Q, CK, D);
    output Q;
    input CK;
    input D;

endmodule
module FFDQRHD1X (Q, CK, D, RN);
    output Q;
    input CK;
    input D;
    input RN;

endmodule
module FFDQRHD2X (Q, CK, D, RN);
    output Q;
    input CK;
    input D;
    input RN;

endmodule
module FFDQRHDLX (Q, CK, D, RN);
    output Q;
    input CK;
    input D;
    input RN;

endmodule
module FFDQRHDMX (Q, CK, D, RN);
    output Q;
    input CK;
    input D;
    input RN;

endmodule
module FFDQSHD1X (Q, CK, D, SN);
    output Q;
    input CK;
    input D;
    input SN;

endmodule
module FFDQSHD2X (Q, CK, D, SN);
    output Q;
    input CK;
    input D;
    input SN;

endmodule
module FFDQSHDLX (Q, CK, D, SN);
    output Q;
    input CK;
    input D;
    input SN;

endmodule
module FFDQSHDMX (Q, CK, D, SN);
    output Q;
    input CK;
    input D;
    input SN;

endmodule
module FFDQSRHD1X (Q, CK, D, RN, SN);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDQSRHD2X (Q, CK, D, RN, SN);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDQSRHDLX (Q, CK, D, RN, SN);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDQSRHDMX (Q, CK, D, RN, SN);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDRHD1X (Q, QN, CK, D, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;

endmodule
module FFDRHD2X (Q, QN, CK, D, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;

endmodule
module FFDRHDLX (Q, QN, CK, D, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;

endmodule
module FFDRHDMX (Q, QN, CK, D, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;

endmodule
module FFDRHQHD1X (Q, CK, D, RN);
    output Q;
    input CK;
    input D;
    input RN;

endmodule
module FFDRHQHD2X (Q, CK, D, RN);
    output Q;
    input CK;
    input D;
    input RN;

endmodule
module FFDRHQHD3X (Q, CK, D, RN);
    output Q;
    input CK;
    input D;
    input RN;

endmodule
module FFDRHQHDMX (Q, CK, D, RN);
    output Q;
    input CK;
    input D;
    input RN;

endmodule
module FFDSHD1X (Q, QN, CK, D, SN);
    output Q;
    output QN;
    input CK;
    input D;
    input SN;

endmodule
module FFDSHD2X (Q, QN, CK, D, SN);
    output Q;
    output QN;
    input CK;
    input D;
    input SN;

endmodule
module FFDSHDLX (Q, QN, CK, D, SN);
    output Q;
    output QN;
    input CK;
    input D;
    input SN;

endmodule
module FFDSHDMX (Q, QN, CK, D, SN);
    output Q;
    output QN;
    input CK;
    input D;
    input SN;

endmodule
module FFDSHQHD1X (Q, CK, D, SN);
    output Q;
    input CK;
    input D;
    input SN;

endmodule
module FFDSHQHD2X (Q, CK, D, SN);
    output Q;
    input CK;
    input D;
    input SN;

endmodule
module FFDSHQHD3X (Q, CK, D, SN);
    output Q;
    input CK;
    input D;
    input SN;

endmodule
module FFDSHQHDMX (Q, CK, D, SN);
    output Q;
    input CK;
    input D;
    input SN;

endmodule
module FFDSRHD1X (Q, QN, CK, D, RN, SN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDSRHD2X (Q, QN, CK, D, RN, SN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDSRHDLX (Q, QN, CK, D, RN, SN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDSRHDMX (Q, QN, CK, D, RN, SN);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDSRHQHD1X (Q, CK, D, RN, SN);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDSRHQHD2X (Q, CK, D, RN, SN);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDSRHQHD3X (Q, CK, D, RN, SN);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFDSRHQHDMX (Q, CK, D, RN, SN);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;

endmodule
module FFEDCRHD1X (Q, QN, CK, D, E, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input RN;

endmodule
module FFEDCRHD2X (Q, QN, CK, D, E, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input RN;

endmodule
module FFEDCRHDLX (Q, QN, CK, D, E, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input RN;

endmodule
module FFEDCRHDMX (Q, QN, CK, D, E, RN);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input RN;

endmodule
module FFEDHD1X (Q, QN, CK, D, E);
    output Q;
    output QN;
    input CK;
    input D;
    input E;

endmodule
module FFEDHD2X (Q, QN, CK, D, E);
    output Q;
    output QN;
    input CK;
    input D;
    input E;

endmodule
module FFEDHDLX (Q, QN, CK, D, E);
    output Q;
    output QN;
    input CK;
    input D;
    input E;

endmodule
module FFEDHDMX (Q, QN, CK, D, E);
    output Q;
    output QN;
    input CK;
    input D;
    input E;

endmodule
module FFEDHQHD1X (Q, CK, D, E);
    output Q;
    input CK;
    input D;
    input E;

endmodule
module FFEDHQHD2X (Q, CK, D, E);
    output Q;
    input CK;
    input D;
    input E;

endmodule
module FFEDHQHD3X (Q, CK, D, E);
    output Q;
    input CK;
    input D;
    input E;

endmodule
module FFEDHQHDMX (Q, CK, D, E);
    output Q;
    input CK;
    input D;
    input E;

endmodule
module FFEDQHD1X (Q, CK, D, E);
    output Q;
    input CK;
    input D;
    input E;

endmodule
module FFEDQHD2X (Q, CK, D, E);
    output Q;
    input CK;
    input D;
    input E;

endmodule
module FFEDQHDLX (Q, CK, D, E);
    output Q;
    input CK;
    input D;
    input E;

endmodule
module FFEDQHDMX (Q, CK, D, E);
    output Q;
    input CK;
    input D;
    input E;

endmodule
module FFSDCRHD1X (Q, QN, CK, D, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDCRHD2X (Q, QN, CK, D, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDCRHDLX (Q, QN, CK, D, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDCRHDMX (Q, QN, CK, D, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDHD1X (Q, QN, CK, D, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDHD1XSPG (Q, QN, CK, D, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDHD2X (Q, QN, CK, D, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDHDLX (Q, QN, CK, D, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDHDMX (Q, QN, CK, D, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDHQHD1X (Q, CK, D, TE, TI);
    output Q;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDHQHD2X (Q, CK, D, TE, TI);
    output Q;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDHQHD3X (Q, CK, D, TE, TI);
    output Q;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDHQHDMX (Q, CK, D, TE, TI);
    output Q;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDNHD1X (Q, QN, CKN, D, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input TE;
    input TI;

endmodule
module FFSDNHD2X (Q, QN, CKN, D, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input TE;
    input TI;

endmodule
module FFSDNHDLX (Q, QN, CKN, D, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input TE;
    input TI;

endmodule
module FFSDNHDMX (Q, QN, CKN, D, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input TE;
    input TI;

endmodule
module FFSDNRHD1X (Q, QN, CKN, D, RN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDNRHD2X (Q, QN, CKN, D, RN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDNRHDLX (Q, QN, CKN, D, RN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDNRHDMX (Q, QN, CKN, D, RN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDNSHD1X (Q, QN, CKN, D, SN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDNSHD2X (Q, QN, CKN, D, SN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDNSHDLX (Q, QN, CKN, D, SN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDNSHDMX (Q, QN, CKN, D, SN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDNSRHD1X (Q, QN, CKN, D, RN, SN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDNSRHD2X (Q, QN, CKN, D, RN, SN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDNSRHDLX (Q, QN, CKN, D, RN, SN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDNSRHDMX (Q, QN, CKN, D, RN, SN, TE, TI);
    output Q;
    output QN;
    input CKN;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDQHD1X (Q, CK, D, TE, TI);
    output Q;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDQHD2X (Q, CK, D, TE, TI);
    output Q;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDQHDLX (Q, CK, D, TE, TI);
    output Q;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDQHDMX (Q, CK, D, TE, TI);
    output Q;
    input CK;
    input D;
    input TE;
    input TI;

endmodule
module FFSDQRHD1X (Q, CK, D, RN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDQRHD2X (Q, CK, D, RN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDQRHDLX (Q, CK, D, RN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDQRHDMX (Q, CK, D, RN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDQSHD1X (Q, CK, D, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDQSHD2X (Q, CK, D, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDQSHDLX (Q, CK, D, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDQSHDMX (Q, CK, D, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDQSRHD1X (Q, CK, D, RN, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDQSRHD2X (Q, CK, D, RN, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDQSRHDLX (Q, CK, D, RN, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDQSRHDMX (Q, CK, D, RN, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDRHD1X (Q, QN, CK, D, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDRHD2X (Q, QN, CK, D, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDRHDLX (Q, QN, CK, D, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDRHDMX (Q, QN, CK, D, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDRHQHD1X (Q, CK, D, RN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDRHQHD2X (Q, CK, D, RN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDRHQHD3X (Q, CK, D, RN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDRHQHDMX (Q, CK, D, RN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input TE;
    input TI;

endmodule
module FFSDSHD1X (Q, QN, CK, D, SN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSHD2X (Q, QN, CK, D, SN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSHDLX (Q, QN, CK, D, SN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSHDMX (Q, QN, CK, D, SN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSHQHD1X (Q, CK, D, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSHQHD2X (Q, CK, D, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSHQHD3X (Q, CK, D, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSHQHDMX (Q, CK, D, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSRHD1X (Q, QN, CK, D, RN, SN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSRHD2X (Q, QN, CK, D, RN, SN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSRHDLX (Q, QN, CK, D, RN, SN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSRHDMX (Q, QN, CK, D, RN, SN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSRHQHD1X (Q, CK, D, RN, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSRHQHD2X (Q, CK, D, RN, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSRHQHD3X (Q, CK, D, RN, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSDSRHQHDMX (Q, CK, D, RN, SN, TE, TI);
    output Q;
    input CK;
    input D;
    input RN;
    input SN;
    input TE;
    input TI;

endmodule
module FFSEDCRHD1X (Q, QN, CK, D, E, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input RN;
    input TE;
    input TI;

endmodule
module FFSEDCRHD2X (Q, QN, CK, D, E, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input RN;
    input TE;
    input TI;

endmodule
module FFSEDCRHDLX (Q, QN, CK, D, E, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input RN;
    input TE;
    input TI;

endmodule
module FFSEDCRHDMX (Q, QN, CK, D, E, RN, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input RN;
    input TE;
    input TI;

endmodule
module FFSEDHD1X (Q, QN, CK, D, E, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDHD2X (Q, QN, CK, D, E, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDHDLX (Q, QN, CK, D, E, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDHDMX (Q, QN, CK, D, E, TE, TI);
    output Q;
    output QN;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDHQHD1X (Q, CK, D, E, TE, TI);
    output Q;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDHQHD2X (Q, CK, D, E, TE, TI);
    output Q;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDHQHD3X (Q, CK, D, E, TE, TI);
    output Q;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDHQHDMX (Q, CK, D, E, TE, TI);
    output Q;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDQHD1X (Q, CK, D, E, TE, TI);
    output Q;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDQHD2X (Q, CK, D, E, TE, TI);
    output Q;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDQHDLX (Q, CK, D, E, TE, TI);
    output Q;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FFSEDQHDMX (Q, CK, D, E, TE, TI);
    output Q;
    input CK;
    input D;
    input E;
    input TE;
    input TI;

endmodule
module FILLER16HD ;

endmodule
module FILLER1HD ;

endmodule
module FILLER2HD ;

endmodule
module FILLER32HD ;

endmodule
module FILLER3HD ;

endmodule
module FILLER4HD ;

endmodule
module FILLER64HD ;

endmodule
module FILLER6HD ;

endmodule
module FILLER8HD ;

endmodule
module FILLERC16HD ;

endmodule
module FILLERC1HD ;

endmodule
module FILLERC2HD ;

endmodule
module FILLERC32HD ;

endmodule
module FILLERC3HD ;

endmodule
module FILLERC4HD ;

endmodule
module FILLERC64HD ;

endmodule
module FILLERC6HD ;

endmodule
module FILLERC8HD ;

endmodule
module HAHD1X (CO, S, A, B);
    output CO;
    output S;
    input A;
    input B;

endmodule
module HAHD2X (CO, S, A, B);
    output CO;
    output S;
    input A;
    input B;

endmodule
module HAHDLX (CO, S, A, B);
    output CO;
    output S;
    input A;
    input B;

endmodule
module HAHDMX (CO, S, A, B);
    output CO;
    output S;
    input A;
    input B;

endmodule
module HOLDHD (Z);
    inout Z;

endmodule
module INVCLKHD10X (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD12X (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD14X (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD16X (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD1X (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD20X (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD2X (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD30X (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD3X (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD40X (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD4X (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD5X (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD6X (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD7X (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD80X (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHD8X (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHDLX (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHDMX (Z, A);
    output Z;
    input A;

endmodule
module INVCLKHDUX (Z, A);
    output Z;
    input A;

endmodule
module INVHD12X (Z, A);
    output Z;
    input A;

endmodule
module INVHD16X (Z, A);
    output Z;
    input A;

endmodule
module INVHD1X (Z, A);
    output Z;
    input A;

endmodule
module INVHD1XSPG (Z, A);
    output Z;
    input A;

endmodule
module INVHD20X (Z, A);
    output Z;
    input A;

endmodule
module INVHD2X (Z, A);
    output Z;
    input A;

endmodule
module INVHD3X (Z, A);
    output Z;
    input A;

endmodule
module INVHD4X (Z, A);
    output Z;
    input A;

endmodule
module INVHD5X (Z, A);
    output Z;
    input A;

endmodule
module INVHD6X (Z, A);
    output Z;
    input A;

endmodule
module INVHD7X (Z, A);
    output Z;
    input A;

endmodule
module INVHD8X (Z, A);
    output Z;
    input A;

endmodule
module INVHDLX (Z, A);
    output Z;
    input A;

endmodule
module INVHDMX (Z, A);
    output Z;
    input A;

endmodule
module INVHDPX (Z, A);
    output Z;
    input A;

endmodule
module INVHDUX (Z, A);
    output Z;
    input A;

endmodule
module INVODHD8X (Z0, Z1, Z2, Z3, Z4, Z5, Z6, Z7, A);
    output Z0;
    output Z1;
    output Z2;
    output Z3;
    output Z4;
    output Z5;
    output Z6;
    output Z7;
    input A;

endmodule
module INVTSHD12X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD16X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD1X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD20X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD2X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD3X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD4X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD5X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD6X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD7X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHD8X (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHDLX (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHDMX (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module INVTSHDUX (Z, A, E);
    output Z;
    input A;
    input E;

endmodule
module LATHD1X (Q, QN, D, G);
    output Q;
    output QN;
    input D;
    input G;

endmodule
module LATHD1XSPG (Q, QN, D, G);
    output Q;
    output QN;
    input D;
    input G;

endmodule
module LATHD2X (Q, QN, D, G);
    output Q;
    output QN;
    input D;
    input G;

endmodule
module LATHDLX (Q, QN, D, G);
    output Q;
    output QN;
    input D;
    input G;

endmodule
module LATHDMX (Q, QN, D, G);
    output Q;
    output QN;
    input D;
    input G;

endmodule
module LATNHD1X (Q, QN, D, GN);
    output Q;
    output QN;
    input D;
    input GN;

endmodule
module LATNHD2X (Q, QN, D, GN);
    output Q;
    output QN;
    input D;
    input GN;

endmodule
module LATNHDLX (Q, QN, D, GN);
    output Q;
    output QN;
    input D;
    input GN;

endmodule
module LATNHDMX (Q, QN, D, GN);
    output Q;
    output QN;
    input D;
    input GN;

endmodule
module LATNRHD1X (Q, QN, D, GN, RN);
    output Q;
    output QN;
    input D;
    input GN;
    input RN;

endmodule
module LATNRHD2X (Q, QN, D, GN, RN);
    output Q;
    output QN;
    input D;
    input GN;
    input RN;

endmodule
module LATNRHDLX (Q, QN, D, GN, RN);
    output Q;
    output QN;
    input D;
    input GN;
    input RN;

endmodule
module LATNRHDMX (Q, QN, D, GN, RN);
    output Q;
    output QN;
    input D;
    input GN;
    input RN;

endmodule
module LATNSHD1X (Q, QN, D, GN, SN);
    output Q;
    output QN;
    input D;
    input GN;
    input SN;

endmodule
module LATNSHD2X (Q, QN, D, GN, SN);
    output Q;
    output QN;
    input D;
    input GN;
    input SN;

endmodule
module LATNSHDLX (Q, QN, D, GN, SN);
    output Q;
    output QN;
    input D;
    input GN;
    input SN;

endmodule
module LATNSHDMX (Q, QN, D, GN, SN);
    output Q;
    output QN;
    input D;
    input GN;
    input SN;

endmodule
module LATNSRHD1X (Q, QN, D, GN, RN, SN);
    output Q;
    output QN;
    input D;
    input GN;
    input RN;
    input SN;

endmodule
module LATNSRHD2X (Q, QN, D, GN, RN, SN);
    output Q;
    output QN;
    input D;
    input GN;
    input RN;
    input SN;

endmodule
module LATNSRHDLX (Q, QN, D, GN, RN, SN);
    output Q;
    output QN;
    input D;
    input GN;
    input RN;
    input SN;

endmodule
module LATNSRHDMX (Q, QN, D, GN, RN, SN);
    output Q;
    output QN;
    input D;
    input GN;
    input RN;
    input SN;

endmodule
module LATRHD1X (Q, QN, D, G, RN);
    output Q;
    output QN;
    input D;
    input G;
    input RN;

endmodule
module LATRHD2X (Q, QN, D, G, RN);
    output Q;
    output QN;
    input D;
    input G;
    input RN;

endmodule
module LATRHDLX (Q, QN, D, G, RN);
    output Q;
    output QN;
    input D;
    input G;
    input RN;

endmodule
module LATRHDMX (Q, QN, D, G, RN);
    output Q;
    output QN;
    input D;
    input G;
    input RN;

endmodule
module LATSHD1X (Q, QN, D, G, SN);
    output Q;
    output QN;
    input D;
    input G;
    input SN;

endmodule
module LATSHD2X (Q, QN, D, G, SN);
    output Q;
    output QN;
    input D;
    input G;
    input SN;

endmodule
module LATSHDLX (Q, QN, D, G, SN);
    output Q;
    output QN;
    input D;
    input G;
    input SN;

endmodule
module LATSHDMX (Q, QN, D, G, SN);
    output Q;
    output QN;
    input D;
    input G;
    input SN;

endmodule
module LATSRHD1X (Q, QN, D, G, RN, SN);
    output Q;
    output QN;
    input D;
    input G;
    input RN;
    input SN;

endmodule
module LATSRHD2X (Q, QN, D, G, RN, SN);
    output Q;
    output QN;
    input D;
    input G;
    input RN;
    input SN;

endmodule
module LATSRHDLX (Q, QN, D, G, RN, SN);
    output Q;
    output QN;
    input D;
    input G;
    input RN;
    input SN;

endmodule
module LATSRHDMX (Q, QN, D, G, RN, SN);
    output Q;
    output QN;
    input D;
    input G;
    input RN;
    input SN;

endmodule
module LATTSHD1X (Q, D, E, G);
    output Q;
    input D;
    input E;
    input G;

endmodule
module LATTSHD2X (Q, D, E, G);
    output Q;
    input D;
    input E;
    input G;

endmodule
module LATTSHDLX (Q, D, E, G);
    output Q;
    input D;
    input E;
    input G;

endmodule
module LATTSHDMX (Q, D, E, G);
    output Q;
    input D;
    input E;
    input G;

endmodule
module MUX2CLKHD1X (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2CLKHD2X (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2CLKHD3X (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2CLKHD4X (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2HD1X (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2HD1XSPG (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2HD2X (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2HD3X (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2HDLX (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2HDMX (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX2HDUX (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUX4HD1X (Z, A, B, C, D, S0, S1);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input S0;
    input S1;

endmodule
module MUX4HD2X (Z, A, B, C, D, S0, S1);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input S0;
    input S1;

endmodule
module MUX4HDLX (Z, A, B, C, D, S0, S1);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input S0;
    input S1;

endmodule
module MUX4HDMX (Z, A, B, C, D, S0, S1);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input S0;
    input S1;

endmodule
module MUXI2HD1X (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUXI2HD2X (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUXI2HD3X (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUXI2HDLX (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUXI2HDMX (Z, A, B, S0);
    output Z;
    input A;
    input B;
    input S0;

endmodule
module MUXI4HD1X (Z, A, B, C, D, S0, S1);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input S0;
    input S1;

endmodule
module MUXI4HD2X (Z, A, B, C, D, S0, S1);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input S0;
    input S1;

endmodule
module MUXI4HDLX (Z, A, B, C, D, S0, S1);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input S0;
    input S1;

endmodule
module MUXI4HDMX (Z, A, B, C, D, S0, S1);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input S0;
    input S1;

endmodule
module NAND2B1HD1X (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NAND2B1HD2X (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NAND2B1HDLX (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NAND2B1HDMX (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NAND2B1HDUX (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NAND2HD1X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NAND2HD1XSPG (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NAND2HD2X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NAND2HD2XSPG (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NAND2HD3X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NAND2HDLX (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NAND2HDMX (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NAND2HDUX (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NAND2ODHD (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NAND3B1HD1X (Z, AN, B, C);
    output Z;
    input AN;
    input B;
    input C;

endmodule
module NAND3B1HD2X (Z, AN, B, C);
    output Z;
    input AN;
    input B;
    input C;

endmodule
module NAND3B1HDLX (Z, AN, B, C);
    output Z;
    input AN;
    input B;
    input C;

endmodule
module NAND3B1HDMX (Z, AN, B, C);
    output Z;
    input AN;
    input B;
    input C;

endmodule
module NAND3HD1X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NAND3HD2X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NAND3HD3X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NAND3HDLX (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NAND3HDMX (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NAND3ODHD (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NAND4B1HD1X (Z, AN, B, C, D);
    output Z;
    input AN;
    input B;
    input C;
    input D;

endmodule
module NAND4B1HD2X (Z, AN, B, C, D);
    output Z;
    input AN;
    input B;
    input C;
    input D;

endmodule
module NAND4B1HDLX (Z, AN, B, C, D);
    output Z;
    input AN;
    input B;
    input C;
    input D;

endmodule
module NAND4B1HDMX (Z, AN, B, C, D);
    output Z;
    input AN;
    input B;
    input C;
    input D;

endmodule
module NAND4B2HD1X (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module NAND4B2HD2X (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module NAND4B2HDLX (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module NAND4B2HDMX (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module NAND4HD1X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module NAND4HD2X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module NAND4HD3X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module NAND4HDLX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module NAND4HDMX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module NOR2B1HD1X (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NOR2B1HD2X (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NOR2B1HDLX (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NOR2B1HDMX (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NOR2B1HDUX (Z, AN, B);
    output Z;
    input AN;
    input B;

endmodule
module NOR2HD1X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NOR2HD1XSPG (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NOR2HD2X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NOR2HD2XSPG (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NOR2HD3X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NOR2HDLX (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NOR2HDMX (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NOR2HDUX (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module NOR3B1HD1X (Z, AN, B, C);
    output Z;
    input AN;
    input B;
    input C;

endmodule
module NOR3B1HD2X (Z, AN, B, C);
    output Z;
    input AN;
    input B;
    input C;

endmodule
module NOR3B1HDLX (Z, AN, B, C);
    output Z;
    input AN;
    input B;
    input C;

endmodule
module NOR3B1HDMX (Z, AN, B, C);
    output Z;
    input AN;
    input B;
    input C;

endmodule
module NOR3HD1X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NOR3HD2X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NOR3HD3X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NOR3HDLX (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NOR3HDMX (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module NOR4B1HD1X (Z, AN, B, C, D);
    output Z;
    input AN;
    input B;
    input C;
    input D;

endmodule
module NOR4B1HD2X (Z, AN, B, C, D);
    output Z;
    input AN;
    input B;
    input C;
    input D;

endmodule
module NOR4B1HDLX (Z, AN, B, C, D);
    output Z;
    input AN;
    input B;
    input C;
    input D;

endmodule
module NOR4B1HDMX (Z, AN, B, C, D);
    output Z;
    input AN;
    input B;
    input C;
    input D;

endmodule
module NOR4B2HD1X (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module NOR4B2HD2X (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module NOR4B2HDLX (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module NOR4B2HDMX (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module NOR4HD1X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module NOR4HD2X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module NOR4HD3X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module NOR4HDLX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module NOR4HDMX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI211HD1X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI211HD2X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI211HDLX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI211HDMX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI21B2HD1X (Z, AN, BN, C);
    output Z;
    input AN;
    input BN;
    input C;

endmodule
module OAI21B2HD2X (Z, AN, BN, C);
    output Z;
    input AN;
    input BN;
    input C;

endmodule
module OAI21B2HDLX (Z, AN, BN, C);
    output Z;
    input AN;
    input BN;
    input C;

endmodule
module OAI21B2HDMX (Z, AN, BN, C);
    output Z;
    input AN;
    input BN;
    input C;

endmodule
module OAI21HD1X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module OAI21HD2X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module OAI21HDLX (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module OAI21HDMX (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module OAI21HDUX (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module OAI221HD1X (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module OAI221HD2X (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module OAI221HDLX (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module OAI221HDMX (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module OAI222HD1X (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module OAI222HD2X (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module OAI222HDLX (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module OAI222HDMX (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module OAI22B2HD1X (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module OAI22B2HD2X (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module OAI22B2HDLX (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module OAI22B2HDMX (Z, AN, BN, C, D);
    output Z;
    input AN;
    input BN;
    input C;
    input D;

endmodule
module OAI22HD1X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI22HD2X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI22HDLX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI22HDMX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI22HDUX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI31HD1X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI31HD2X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI31HDLX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI31HDMX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OAI32HD1X (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module OAI32HD2X (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module OAI32HDLX (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module OAI32HDMX (Z, A, B, C, D, E);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;

endmodule
module OAI33HD1X (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module OAI33HD2X (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module OAI33HDLX (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module OAI33HDMX (Z, A, B, C, D, E, F);
    output Z;
    input A;
    input B;
    input C;
    input D;
    input E;
    input F;

endmodule
module OR2HD1X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module OR2HD1XSPG (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module OR2HD2X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module OR2HD2XSPG (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module OR2HDLX (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module OR2HDMX (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module OR2HDUX (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module OR2ODHD (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module OR3HD1X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module OR3HD2X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module OR3HDLX (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module OR3HDMX (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module OR4HD1X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OR4HD2X (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OR4HDLX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module OR4HDMX (Z, A, B, C, D);
    output Z;
    input A;
    input B;
    input C;
    input D;

endmodule
module PULLDHD (Z, EN);
    output Z;
    input EN;

endmodule
module PULLUHD (Z, E);
    output Z;
    input E;

endmodule
module RSLATHD1X (Q, QN, R, S);
    output Q;
    output QN;
    input R;
    input S;

endmodule
module RSLATHD2X (Q, QN, R, S);
    output Q;
    output QN;
    input R;
    input S;

endmodule
module RSLATHDLX (Q, QN, R, S);
    output Q;
    output QN;
    input R;
    input S;

endmodule
module RSLATHDMX (Q, QN, R, S);
    output Q;
    output QN;
    input R;
    input S;

endmodule
module RSLATNHD1X (Q, QN, RN, SN);
    output Q;
    output QN;
    input RN;
    input SN;

endmodule
module RSLATNHD2X (Q, QN, RN, SN);
    output Q;
    output QN;
    input RN;
    input SN;

endmodule
module RSLATNHDLX (Q, QN, RN, SN);
    output Q;
    output QN;
    input RN;
    input SN;

endmodule
module RSLATNHDMX (Q, QN, RN, SN);
    output Q;
    output QN;
    input RN;
    input SN;

endmodule
module TIEHHD (Z);
    output Z;

endmodule
module TIELHD (Z);
    output Z;

endmodule
module XNOR2HD1X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XNOR2HD2X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XNOR2HD3X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XNOR2HDLX (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XNOR2HDMX (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XNOR3HD1X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module XNOR3HD2X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module XNOR3HD3X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module XNOR3HDLX (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module XNOR3HDMX (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module XOR2CLKHD1X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XOR2CLKHD2X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XOR2CLKHD3X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XOR2CLKHD4X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XOR2HD1X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XOR2HD2X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XOR2HD3X (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XOR2HDLX (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XOR2HDMX (Z, A, B);
    output Z;
    input A;
    input B;

endmodule
module XOR3HD1X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module XOR3HD2X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module XOR3HD3X (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module XOR3HDLX (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
module XOR3HDMX (Z, A, B, C);
    output Z;
    input A;
    input B;
    input C;

endmodule
