MACRO PSBI16F
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 6.5676 LAYER M2 ;
    AntennaDiffArea 6.5676 LAYER M3 ;
    AntennaDiffArea 6.5676 LAYER M4 ;
    AntennaDiffArea 6.5676 LAYER M5 ;
    AntennaDiffArea 6.5676 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 2417.89 LAYER M3 ;
    AntennaDiffArea 2417.89 LAYER M4 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PSBI16F
MACRO PSBI16N
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 6.5676 LAYER M2 ;
    AntennaDiffArea 6.5676 LAYER M3 ;
    AntennaDiffArea 6.5676 LAYER M4 ;
    AntennaDiffArea 6.5676 LAYER M5 ;
    AntennaDiffArea 6.5676 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 2417.89 LAYER M3 ;
    AntennaDiffArea 2417.89 LAYER M4 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PSBI16N
MACRO PSBI16S
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 6.5676 LAYER M2 ;
    AntennaDiffArea 6.5676 LAYER M3 ;
    AntennaDiffArea 6.5676 LAYER M4 ;
    AntennaDiffArea 6.5676 LAYER M5 ;
    AntennaDiffArea 6.5676 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 2417.89 LAYER M3 ;
    AntennaDiffArea 2417.89 LAYER M4 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PSBI16S
MACRO PSBI24F
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 6.5676 LAYER M2 ;
    AntennaDiffArea 6.5676 LAYER M3 ;
    AntennaDiffArea 6.5676 LAYER M4 ;
    AntennaDiffArea 6.5676 LAYER M5 ;
    AntennaDiffArea 6.5676 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 2417.89 LAYER M3 ;
    AntennaDiffArea 2417.89 LAYER M4 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PSBI24F
MACRO PSBI24N
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 6.5676 LAYER M2 ;
    AntennaDiffArea 6.5676 LAYER M3 ;
    AntennaDiffArea 6.5676 LAYER M4 ;
    AntennaDiffArea 6.5676 LAYER M5 ;
    AntennaDiffArea 6.5676 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 2417.89 LAYER M3 ;
    AntennaDiffArea 2417.89 LAYER M4 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PSBI24N
MACRO PSBI24S
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 6.5676 LAYER M2 ;
    AntennaDiffArea 6.5676 LAYER M3 ;
    AntennaDiffArea 6.5676 LAYER M4 ;
    AntennaDiffArea 6.5676 LAYER M5 ;
    AntennaDiffArea 6.5676 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 2417.89 LAYER M3 ;
    AntennaDiffArea 2417.89 LAYER M4 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PSBI24S
MACRO PSBI2F
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 6.5676 LAYER M2 ;
    AntennaDiffArea 6.5676 LAYER M3 ;
    AntennaDiffArea 6.5676 LAYER M4 ;
    AntennaDiffArea 6.5676 LAYER M5 ;
    AntennaDiffArea 6.5676 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 2417.89 LAYER M3 ;
    AntennaDiffArea 2417.89 LAYER M4 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PSBI2F
MACRO PSBI2N
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 6.5676 LAYER M2 ;
    AntennaDiffArea 6.5676 LAYER M3 ;
    AntennaDiffArea 6.5676 LAYER M4 ;
    AntennaDiffArea 6.5676 LAYER M5 ;
    AntennaDiffArea 6.5676 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 2417.89 LAYER M3 ;
    AntennaDiffArea 2417.89 LAYER M4 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PSBI2N
MACRO PSBI2S
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 6.5676 LAYER M2 ;
    AntennaDiffArea 6.5676 LAYER M3 ;
    AntennaDiffArea 6.5676 LAYER M4 ;
    AntennaDiffArea 6.5676 LAYER M5 ;
    AntennaDiffArea 6.5676 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 2417.89 LAYER M3 ;
    AntennaDiffArea 2417.89 LAYER M4 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PSBI2S
MACRO PSBI4F
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 6.5676 LAYER M2 ;
    AntennaDiffArea 6.5676 LAYER M3 ;
    AntennaDiffArea 6.5676 LAYER M4 ;
    AntennaDiffArea 6.5676 LAYER M5 ;
    AntennaDiffArea 6.5676 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 2417.89 LAYER M3 ;
    AntennaDiffArea 2417.89 LAYER M4 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PSBI4F
MACRO PSBI4N
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 6.5676 LAYER M2 ;
    AntennaDiffArea 6.5676 LAYER M3 ;
    AntennaDiffArea 6.5676 LAYER M4 ;
    AntennaDiffArea 6.5676 LAYER M5 ;
    AntennaDiffArea 6.5676 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 2417.89 LAYER M3 ;
    AntennaDiffArea 2417.89 LAYER M4 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PSBI4N
MACRO PSBI4S
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 6.5676 LAYER M2 ;
    AntennaDiffArea 6.5676 LAYER M3 ;
    AntennaDiffArea 6.5676 LAYER M4 ;
    AntennaDiffArea 6.5676 LAYER M5 ;
    AntennaDiffArea 6.5676 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 2417.89 LAYER M3 ;
    AntennaDiffArea 2417.89 LAYER M4 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PSBI4S
MACRO PSBI8F
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 6.5676 LAYER M2 ;
    AntennaDiffArea 6.5676 LAYER M3 ;
    AntennaDiffArea 6.5676 LAYER M4 ;
    AntennaDiffArea 6.5676 LAYER M5 ;
    AntennaDiffArea 6.5676 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 2417.89 LAYER M3 ;
    AntennaDiffArea 2417.89 LAYER M4 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PSBI8F
MACRO PSBI8N
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 6.5676 LAYER M2 ;
    AntennaDiffArea 6.5676 LAYER M3 ;
    AntennaDiffArea 6.5676 LAYER M4 ;
    AntennaDiffArea 6.5676 LAYER M5 ;
    AntennaDiffArea 6.5676 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 2417.89 LAYER M3 ;
    AntennaDiffArea 2417.89 LAYER M4 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PSBI8N
MACRO PSBI8S
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN A
    AntennaGateArea 10.2288 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END A
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN CONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END CONOF
  PIN D
    AntennaDiffArea 6.5676 LAYER M2 ;
    AntennaDiffArea 6.5676 LAYER M3 ;
    AntennaDiffArea 6.5676 LAYER M4 ;
    AntennaDiffArea 6.5676 LAYER M5 ;
    AntennaDiffArea 6.5676 LAYER M6 ;
  END D
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN NEN
    AntennaGateArea 2.2648 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END NEN
  PIN P
    AntennaDiffArea 2417.89 LAYER M3 ;
    AntennaDiffArea 2417.89 LAYER M4 ;
  END P
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PD
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PD
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PEN
    AntennaGateArea 4.5296 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PEN
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN PU
    AntennaGateArea 1.8212 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END PU
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
  PIN SONOF
    AntennaGateArea 4.085 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END SONOF
END PSBI8S
MACRO PSBIA
  PIN P
    AntennaDiffArea 3113.2 LAYER M3 ;
    AntennaDiffArea 3113.2 LAYER M4 ;
    AntennaDiffArea 3113.2 LAYER M5 ;
    AntennaDiffArea 3113.2 LAYER M6 ;
  END P
END PSBIA
MACRO PSBIAR
  PIN AI
    AntennaDiffArea 3113.2 LAYER M3 ;
    AntennaDiffArea 3113.2 LAYER M4 ;
    AntennaDiffArea 3113.2 LAYER M5 ;
    AntennaDiffArea 3113.2 LAYER M6 ;
  END AI
END PSBIAR
MACRO PSOSC14M
  PIN CK
    AntennaDiffArea 23.89 LAYER M2 ;
    AntennaDiffArea 23.89 LAYER M3 ;
    AntennaDiffArea 23.89 LAYER M4 ;
    AntennaDiffArea 23.89 LAYER M5 ;
    AntennaDiffArea 23.89 LAYER M6 ;
  END CK
  PIN EI
    AntennaGateArea 3.14 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END EI
  PIN EI
    AntennaGateArea 3.14 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END EI
  PIN EO
    AntennaGateArea 3.14 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END EO
  PIN EO
    AntennaGateArea 3.14 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END EO
  PIN XTALIN
    AntennaGateArea 61.2 ;
    AntennaDiffArea 3125.4 LAYER M3 ;
    AntennaDiffArea 3125.4 LAYER M4 ;
  END XTALIN
  PIN XTALIN
    AntennaGateArea 61.2 ;
    AntennaDiffArea 3125.4 LAYER M3 ;
    AntennaDiffArea 3125.4 LAYER M4 ;
  END XTALIN
  PIN XTALOUT
    AntennaDiffArea 3158.97 LAYER M3 ;
    AntennaDiffArea 3158.97 LAYER M4 ;
  END XTALOUT
END PSOSC14M
MACRO PSOSCR14M
  PIN CK
    AntennaDiffArea 24.73 LAYER M2 ;
    AntennaDiffArea 24.73 LAYER M3 ;
    AntennaDiffArea 24.73 LAYER M4 ;
    AntennaDiffArea 24.73 LAYER M5 ;
    AntennaDiffArea 24.73 LAYER M6 ;
  END CK
  PIN EI
    AntennaGateArea 3.5062 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END EI
  PIN EI
    AntennaGateArea 3.5062 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END EI
  PIN EO
    AntennaGateArea 3.5062 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END EO
  PIN EO
    AntennaGateArea 3.5062 ;
    AntennaDiffArea 0.25 LAYER M2 ;
    AntennaDiffArea 0.25 LAYER M3 ;
    AntennaDiffArea 0.25 LAYER M4 ;
    AntennaDiffArea 0.25 LAYER M5 ;
    AntennaDiffArea 0.25 LAYER M6 ;
  END EO
  PIN XTALIN
    AntennaGateArea 1971.24 ;
    AntennaDiffArea 3126.44 LAYER M3 ;
    AntennaDiffArea 3126.44 LAYER M4 ;
  END XTALIN
  PIN XTALIN
    AntennaGateArea 1971.24 ;
    AntennaDiffArea 3126.44 LAYER M3 ;
    AntennaDiffArea 3126.44 LAYER M4 ;
  END XTALIN
  PIN XTALOUT
    AntennaGateArea 1800 ;
    AntennaDiffArea 3186.71 LAYER M3 ;
    AntennaDiffArea 3186.71 LAYER M4 ;
  END XTALOUT
  PIN XTALOUT
    AntennaGateArea 1800 ;
    AntennaDiffArea 3186.71 LAYER M3 ;
    AntennaDiffArea 3186.71 LAYER M4 ;
  END XTALOUT
END PSOSCR14M
END LIBRARY
