VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS

LAYER M1
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		0.41  ;
  WIDTH         0.16 ;
  SPACING       0.18 ;
  SPACING 0.18 LENGTHTHRESHOLD  1.0 ;
  SPACING 0.20 RANGE 0.4 10.005 USELENGTHTHRESHOLD ;
  SPACING 0.6 RANGE 10 1000 USELENGTHTHRESHOLD ;
  SPACING 0.6 RANGE 10 1000 INFLUENCE 1 ;
  RESISTANCE	RPERSQ 0.1038 ;
  CAPACITANCE	CPERSQDIST 0.000195 ;
  EDGECAPACITANCE 8.79e-05 ;
  HEIGHT 1.17 ;
  THICKNESS 0.26 ;
END M1

LAYER V1
  TYPE	CUT ;
  SPACING	0.22 ;
END V1

LAYER M2
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		0.41  ;
  WIDTH		0.2 ;
  SPACING 0.21 ;
  SPACING 0.21 LENGTHTHRESHOLD  1.0 ;
  SPACING 0.22 RANGE 0.5 10.005 USELENGTHTHRESHOLD ;
  SPACING 0.6 RANGE 10 1000 USELENGTHTHRESHOLD ;
  SPACING 0.6 RANGE 10 1000 INFLUENCE 1 ;
  RESISTANCE	RPERSQ 0.0591 ;
  CAPACITANCE	CPERSQDIST 0.0001385 ;
  EDGECAPACITANCE 0.0001121 ;
  HEIGHT 1.93 ;
  THICKNESS 0.385 ;
END M2

LAYER V2
  TYPE	CUT ;
  SPACING	0.22 ;
END V2

LAYER M3
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		0.41  ;
  WIDTH         0.2 ;
  SPACING 0.21 ;
  SPACING 0.21 LENGTHTHRESHOLD  1.0 ;
  SPACING 0.22 RANGE 0.5 10.005 USELENGTHTHRESHOLD ;
  SPACING 0.6 RANGE 10 1000 USELENGTHTHRESHOLD ;
  SPACING 0.6 RANGE 10 1000 INFLUENCE 1 ;
  RESISTANCE	RPERSQ 0.0591 ;
  CAPACITANCE	CPERSQDIST 0.000123 ;
  EDGECAPACITANCE 0.0001226 ;
  HEIGHT 2.69 ;
  THICKNESS 0.385 ;
END M3

LAYER V3
  TYPE	CUT ;
  SPACING	0.22 ;
END V3

LAYER M4
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		0.41  ;
  WIDTH         0.2 ;
  SPACING 0.21 ;
  SPACING 0.21 LENGTHTHRESHOLD  1.0 ;
  SPACING 0.22 RANGE 0.5 10.005 USELENGTHTHRESHOLD ;
  SPACING 0.6 RANGE 10 1000 USELENGTHTHRESHOLD ;
  SPACING 0.6 RANGE 10 1000 INFLUENCE 1 ;
  RESISTANCE	RPERSQ 0.0591 ;
  CAPACITANCE	CPERSQDIST 0.0001165 ;
  EDGECAPACITANCE 0.0001222 ;
  HEIGHT 3.45 ;
  THICKNESS 0.385 ;
END M4

LAYER V4
  TYPE	CUT ;
  SPACING	0.22 ;
END V4

LAYER M5
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		0.41  ;
  WIDTH         0.2 ;
  SPACING 0.21 ;
  SPACING 0.21 LENGTHTHRESHOLD  1.0 ;
  SPACING 0.22 RANGE 0.5 10.005 USELENGTHTHRESHOLD ;
  SPACING 0.6 RANGE 10 1000 USELENGTHTHRESHOLD ;
  SPACING 0.6 RANGE 10 1000 INFLUENCE 1 ;
  RESISTANCE	RPERSQ 0.0591 ;
  CAPACITANCE	CPERSQDIST 0.0001262 ;
  EDGECAPACITANCE 0.000123 ;
  HEIGHT 4.21 ;
  THICKNESS 0.385 ;
END M5

LAYER V5
  TYPE	CUT ;
  SPACING	0.22 ;
END V5

LAYER M6
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		0.41  ;
  WIDTH         0.2 ;
  SPACING 0.21 ;
  SPACING 0.21 LENGTHTHRESHOLD  1.0 ;
  SPACING 0.22 RANGE 0.5 10.005 USELENGTHTHRESHOLD ;
  SPACING 0.6 RANGE 10 1000 USELENGTHTHRESHOLD ;
  SPACING 0.6 RANGE 10 1000 INFLUENCE 1 ;
  RESISTANCE	RPERSQ 0.0591 ;
  CAPACITANCE	CPERSQDIST 0.0001151 ;
  EDGECAPACITANCE 0.0001221 ;
  HEIGHT 4.97 ;
  THICKNESS 0.385 ;
END M6

LAYER V6
  TYPE	CUT ;
  SPACING	0.22 ;
END V6

LAYER M7
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		0.5  ;
  WIDTH         0.2 ;
  SPACING 0.21 ;
  SPACING 0.21 LENGTHTHRESHOLD  1.0 ;
  SPACING 0.22 RANGE 0.5 10.005 USELENGTHTHRESHOLD ;
  SPACING 0.6 RANGE 10 1000 USELENGTHTHRESHOLD ;
  SPACING 0.6 RANGE 10 1000 INFLUENCE 1 ;
  RESISTANCE	RPERSQ 0.0591 ;
  CAPACITANCE	CPERSQDIST 9.79e-05 ;
  EDGECAPACITANCE 9.36e-05 ;
  HEIGHT 5.73 ;
  THICKNESS 0.385 ;
END M7

LAYER V7
  TYPE	CUT ;
  SPACING	0.35 ;
END V7

LAYER M8
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		1  ;
  WIDTH		0.44 ;
  SPACING	0.46 ;
  SPACING 0.60 RANGE 10.005 100000.0 ;
  SPACING 0.6 RANGE 0.2 10
  RANGE 10.005  1000 ;
  RESISTANCE	RPERSQ 0.019 ;
  CAPACITANCE	CPERSQDIST 3.72e-05 ;
  EDGECAPACITANCE 0.0001131 ;
  HEIGHT 7.33 ;
  THICKNESS 0.9 ;
END M8

SPACING
  SAMENET M1  M1	0.18 ;
  SAMENET M2  M2	0.21  STACK ;
  SAMENET M3  M3	0.21  STACK ;
  SAMENET M4  M4	0.21  STACK ;
  SAMENET M5  M5	0.21  STACK ;
  SAMENET M6  M6        0.21  STACK ;
  SAMENET M7  M7        0.21  STACK ;
  SAMENET M8  M8        0.46 ;
  SAMENET V1  V1	0.22 ;
  SAMENET V2  V2	0.22 ;
  SAMENET V3  V3	0.22 ;
  SAMENET V4  V4	0.22 ;
  SAMENET V5  V5        0.22 ;
  SAMENET V6  V6        0.22 ;
  SAMENET V7  V7        0.35 ;
  SAMENET V1  V2	0.00  STACK ;
  SAMENET V2  V3	0.00  STACK ;
  SAMENET V3  V4	0.00  STACK ;
  SAMENET V4  V5        0.00  STACK ;
  SAMENET V5  V6        0.00  STACK ;
  SAMENET V6  V7        0.00  STACK ;
  SAMENET M1  V1	0.00 ;
  SAMENET M2  V1	0.00 ;
  SAMENET M2  V2	0.00 ;
  SAMENET M3  V2	0.00 ;
  SAMENET M3  V3	0.00 ;
  SAMENET M4  V3	0.00 ;
  SAMENET M4  V4	0.00 ;
  SAMENET M5  V4	0.00 ;
  SAMENET M5  V5	0.00 ;
  SAMENET M6  V5	0.00 ;
  SAMENET M6  V6	0.00 ;
  SAMENET M7  V6	0.00 ;
  SAMENET M7  V7	0.00 ;
  SAMENET M8  V7	0.00 ;
END SPACING

VIA V12_H DEFAULT
  LAYER M1 ;
    RECT -0.165 -0.105 0.165 0.105 ;
  LAYER V1 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER M2 ;
    RECT -0.100 -0.165 0.100 0.165 ;
  RESISTANCE 6.00 ;
END V12_H

VIA V12_V DEFAULT
  LAYER M1 ;
    RECT -0.105 -0.165 0.105 0.165 ;
  LAYER V1 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER M2 ;
    RECT -0.100 -0.165 0.100 0.165 ;
  RESISTANCE 6.00 ;
END V12_V

VIA V23 DEFAULT
  LAYER M2 ;
    RECT -0.100 -0.165 0.100 0.165 ;
  LAYER V2 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER M3 ;
    RECT -0.165 -0.100 0.165 0.100 ;
  RESISTANCE 6.00 ;
END V23

VIA V34 DEFAULT
  LAYER M3 ;
    RECT -0.165 -0.100 0.165 0.100 ;
  LAYER V3 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER M4 ;
    RECT -0.100 -0.165 0.100 0.165 ;
  RESISTANCE 6.00 ;
END V34

VIA V45 DEFAULT
  LAYER M4 ;
    RECT -0.100 -0.165 0.100 0.165 ;
  LAYER V4 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER M5 ;
    RECT -0.165 -0.100 0.165 0.100 ;
  RESISTANCE 6.00 ;
END V45

VIA V56 DEFAULT
  LAYER M5 ;
    RECT -0.165 -0.100 0.165 0.100 ;
  LAYER V5 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER M6 ;
    RECT -0.100 -0.165 0.100 0.165 ;
  RESISTANCE 6.00 ;
END V56

VIA V23S_NORTH DEFAULT
  TOPOFSTACKONLY
  LAYER M2 ;
    RECT -0.100 -0.165 0.100 0.555 ;
  LAYER V2 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER M3 ;
    RECT -0.165 -0.100 0.165 0.100 ;
  RESISTANCE 6.00 ;
END V23S_NORTH

VIA V23S_SOUTH DEFAULT
  TOPOFSTACKONLY
  LAYER M2 ;
    RECT -0.100 -0.555 0.100 0.165 ;
  LAYER V2 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER M3 ;
    RECT -0.165 -0.100 0.165 0.100 ;
  RESISTANCE 6.00 ;
END V23S_SOUTH

VIA V34S_EAST DEFAULT
  TOPOFSTACKONLY
  LAYER M3 ;
    RECT -0.165 -0.100 0.555 0.100 ;
  LAYER V3 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER M4 ;
    RECT -0.100 -0.165 0.100 0.165 ;
  RESISTANCE 6.00 ;
END V34S_EAST

VIA V34S_WEST DEFAULT
  TOPOFSTACKONLY
  LAYER M3 ;
    RECT -0.555 -0.100 0.165 0.100 ;
  LAYER V3 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER M4 ;
    RECT -0.100 -0.165 0.100 0.165 ;
  RESISTANCE 6.00 ;
END V34S_WEST

VIA V45S_NORTH DEFAULT
  TOPOFSTACKONLY
  LAYER M4 ;
    RECT -0.100 -0.165 0.100 0.555 ;
  LAYER V4 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER M5 ;
    RECT -0.165 -0.100 0.165 0.100 ;
  RESISTANCE 6.00 ;
END V45S_NORTH

VIA V45S_SOUTH DEFAULT
  TOPOFSTACKONLY
  LAYER M4 ;
    RECT -0.100 -0.555 0.100 0.165 ;
  LAYER V4 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER M5 ;
    RECT -0.165 -0.100 0.165 0.100 ;
  RESISTANCE 6.00 ;
END V45S_SOUTH

VIA V56S_EAST DEFAULT
  TOPOFSTACKONLY
  LAYER M5 ;
    RECT -0.165 -0.100 0.555 0.100 ;
  LAYER V5 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER M6 ;
    RECT -0.100 -0.165 0.100 0.165 ;
  RESISTANCE 6.00 ;
END V56S_EAST

VIA V56S_WEST DEFAULT
  TOPOFSTACKONLY
  LAYER M5 ;
    RECT -0.555 -0.100 0.165 0.100 ;
  LAYER V5 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER M6 ;
    RECT -0.100 -0.165 0.100 0.165 ;
  RESISTANCE 6.00 ;
END V56S_WEST

VIA V67S_NORTH DEFAULT
  TOPOFSTACKONLY
  LAYER M6 ;
    RECT -0.100 -0.165 0.100 0.555 ;
  LAYER V6 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER M7 ;
    RECT -0.165 -0.100 0.165 0.100 ;
  RESISTANCE 6.00 ;
END V67S_NORTH

VIA V67S_SOUTH DEFAULT
  TOPOFSTACKONLY
  LAYER M6 ;
    RECT -0.100 -0.555 0.100 0.165 ;
  LAYER V6 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER M7 ;
    RECT -0.165 -0.100 0.165 0.100 ;
  RESISTANCE 6.00 ;
END V67S_SOUTH

VIA V78S DEFAULT
  TOPOFSTACKONLY
  LAYER M7 ;
    RECT -0.360 -0.190 0.360 0.190 ;
  LAYER V7 ;
    RECT -0.180 -0.180 0.180 0.180 ;
  LAYER M8 ;
    RECT -0.270 -0.510 0.270 0.510 ;
  RESISTANCE 6.00 ;
END V78S

VIA V67 DEFAULT
  LAYER M6 ;
    RECT -0.100 -0.165 0.100 0.165 ;
  LAYER V6 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER M7 ;
    RECT -0.165 -0.100 0.165 0.100 ;
  RESISTANCE 6.00 ;
END V67

VIA V78 DEFAULT
  LAYER M7 ;
    RECT -0.250 -0.190 0.250 0.190 ;
  LAYER V7 ;
    RECT -0.180 -0.180 0.180 0.180 ;
  LAYER M8 ;
    RECT -0.270 -0.290 0.270 0.290 ;
  RESISTANCE 6.00 ;
END V78

VIARULE VIAGEN12 GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.07 ;
    METALOVERHANG 0 ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.07 ;
    METALOVERHANG 0 ;
  LAYER V1 ;
    RECT -0.095 -0.095 0.095 0.095 ;
    SPACING 0.48 BY 0.48 ;
END VIAGEN12

VIARULE VIAGEN23 GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.07 ;
    METALOVERHANG 0 ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.07 ;
    METALOVERHANG 0 ;
  LAYER V2 ;
    RECT -0.095 -0.095 0.095 0.095 ;
    SPACING 0.48 BY 0.48 ;
END VIAGEN23

VIARULE VIAGEN34 GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.07 ;
    METALOVERHANG 0 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.07 ;
    METALOVERHANG 0 ;
  LAYER V3 ;
    RECT -0.095 -0.095 0.095 0.095 ;
    SPACING 0.48 BY 0.48 ;
END VIAGEN34

VIARULE TURNM1 GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
  LAYER M1 ;
    DIRECTION VERTICAL ;
END TURNM1

VIARULE TURNM2 GENERATE
  LAYER M2 ;
    DIRECTION HORIZONTAL ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
END TURNM2

VIARULE TURNM3 GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
  LAYER M3 ;
    DIRECTION VERTICAL ;
END TURNM3

VIARULE TURNM4 GENERATE
  LAYER M4 ;
    DIRECTION HORIZONTAL ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
END TURNM4

VIARULE VIAGEN45 GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.07 ;
    METALOVERHANG 0 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.07 ;
    METALOVERHANG 0 ;
  LAYER V4 ;
    RECT -0.095 -0.095 0.095 0.095 ;
    SPACING 0.48 BY 0.48 ;
END VIAGEN45

VIARULE TURNM5 GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
  LAYER M5 ;
    DIRECTION VERTICAL ;
END TURNM5

VIARULE VIAGEN56 GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.07 ;
    METALOVERHANG 0 ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.07 ;
    METALOVERHANG 0 ;
  LAYER V5 ;
    RECT -0.095 -0.095 0.095 0.095 ;
    SPACING 0.48 BY 0.48 ;
END VIAGEN56

VIARULE TURNM6 GENERATE
  LAYER M6 ;
    DIRECTION HORIZONTAL ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
END TURNM6

VIARULE VIAGEN67 GENERATE
  LAYER M7 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.07 ;
    METALOVERHANG 0 ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.07 ;
    METALOVERHANG 0 ;
  LAYER V6 ;
    RECT -0.095 -0.095 0.095 0.095 ;
    SPACING 0.48 BY 0.48 ;
END VIAGEN67

VIARULE TURNM7 GENERATE
  LAYER M7 ;
    DIRECTION HORIZONTAL ;
  LAYER M7 ;
    DIRECTION VERTICAL ;
END TURNM7

VIARULE VIAGEN78 GENERATE
  LAYER M7 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.07 ;
    METALOVERHANG 0 ;
  LAYER M8 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.11 ;
    METALOVERHANG 0 ;
  LAYER V7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.9 BY 0.9 ;
END VIAGEN78

VIARULE TURNM8 GENERATE
  LAYER M8 ;
    DIRECTION HORIZONTAL ;
  LAYER M8 ;
    DIRECTION VERTICAL ;
END TURNM8

SITE  CoreSite
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	0.410 BY 3.690 ;
END  CoreSite

MACRO XOR2CLKHD2XHT
  CLASS  CORE ;
  FOREIGN XOR2CLKHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.510 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.895 1.530 3.240 1.955 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.670 0.585 2.015 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 -0.300 0.860 0.810 ;
        RECT 3.100 -0.300 3.270 0.780 ;
        RECT 4.105 -0.300 4.405 1.060 ;
        RECT 0.000 -0.300 4.510 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.645 2.510 3.820 3.150 ;
        RECT 3.585 1.060 3.885 1.420 ;
        RECT 3.585 1.250 4.410 1.420 ;
        RECT 4.200 1.250 4.410 2.680 ;
        RECT 3.645 2.510 4.410 2.680 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.545 0.925 3.990 ;
        RECT 3.035 3.075 3.335 3.990 ;
        RECT 4.170 2.910 4.340 3.990 ;
        RECT 0.000 3.390 4.510 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 1.480 ;
        RECT 0.870 1.310 1.040 2.365 ;
        RECT 0.105 2.195 1.040 2.365 ;
        RECT 1.180 0.575 1.400 1.480 ;
        RECT 0.170 1.310 1.400 1.480 ;
        RECT 1.180 0.575 2.300 0.745 ;
        RECT 2.130 0.575 2.300 2.395 ;
        RECT 2.480 1.060 2.650 2.335 ;
        RECT 2.480 1.060 2.810 1.360 ;
        RECT 2.480 2.165 2.875 2.335 ;
        RECT 1.580 1.060 1.750 2.780 ;
        RECT 3.240 2.135 3.465 2.780 ;
        RECT 1.580 2.610 3.465 2.780 ;
        RECT 3.465 1.600 3.645 2.315 ;
        RECT 3.240 2.135 3.645 2.315 ;
        RECT 3.465 1.600 3.985 1.900 ;
  END 
END XOR2CLKHD2XHT

MACRO RSLATNHD1XHT
  CLASS  CORE ;
  FOREIGN RSLATNHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.875 1.125 3.045 2.430 ;
        RECT 2.875 1.125 3.175 1.295 ;
        RECT 2.875 2.110 3.300 2.430 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.090 1.235 2.260 2.280 ;
        RECT 2.325 1.125 2.625 1.615 ;
        RECT 2.090 1.235 2.625 1.615 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.485 2.900 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 1.805 -0.300 2.105 1.055 ;
        RECT 3.435 -0.300 3.735 0.595 ;
        RECT 4.590 -0.300 4.785 1.295 ;
        RECT 4.405 1.125 4.785 1.295 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.380 2.010 4.820 2.430 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.100 0.860 3.990 ;
        RECT 2.545 2.975 2.845 3.990 ;
        RECT 4.470 2.610 4.640 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.605 1.030 1.775 ;
        RECT 0.860 1.540 1.030 1.840 ;
        RECT 1.200 0.480 1.500 0.650 ;
        RECT 1.145 1.125 1.500 1.295 ;
        RECT 1.330 0.480 1.500 2.215 ;
        RECT 1.330 2.045 1.815 2.215 ;
        RECT 3.400 1.570 3.630 1.880 ;
        RECT 1.335 2.625 1.635 2.875 ;
        RECT 3.410 1.570 3.630 1.890 ;
        RECT 3.420 1.570 3.630 1.900 ;
        RECT 3.430 1.570 3.630 1.910 ;
        RECT 3.440 1.570 3.630 1.920 ;
        RECT 3.450 1.570 3.630 1.930 ;
        RECT 3.460 1.125 3.630 1.939 ;
        RECT 3.470 1.875 3.650 1.949 ;
        RECT 3.290 1.570 3.630 1.870 ;
        RECT 3.400 1.865 3.640 1.880 ;
        RECT 3.480 1.875 3.650 2.795 ;
        RECT 1.335 2.625 3.815 2.795 ;
        RECT 3.460 1.125 4.185 1.295 ;
        RECT 2.605 0.480 2.905 0.945 ;
        RECT 4.175 0.640 4.410 0.945 ;
        RECT 2.605 0.775 4.410 0.945 ;
        RECT 3.810 1.475 3.980 1.775 ;
        RECT 4.985 1.060 5.170 1.660 ;
        RECT 3.810 1.475 5.170 1.660 ;
        RECT 5.000 1.060 5.170 2.910 ;
        RECT 4.950 2.610 5.170 2.910 ;
  END 
END RSLATNHD1XHT

MACRO PULLDHDHT
  CLASS  CORE ;
  FOREIGN PULLDHDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.860 ;
    END
  END EN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.295 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.235 0.860 1.540 1.295 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.745 2.100 0.915 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.175 1.755 ;
  END 
END PULLDHDHT

MACRO OR3HDMXHT
  CLASS  CORE ;
  FOREIGN OR3HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.850 2.710 1.400 3.180 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.585 0.720 2.020 ;
        RECT 0.510 1.585 1.070 1.755 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.260 0.330 1.820 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.555 -0.300 0.855 1.295 ;
        RECT 1.505 -0.300 1.805 0.715 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.120 1.060 2.360 1.360 ;
        RECT 2.170 1.060 2.360 2.430 ;
        RECT 2.065 2.080 2.360 2.430 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.600 2.310 1.770 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.060 0.505 1.230 1.295 ;
        RECT 1.060 1.125 1.420 1.295 ;
        RECT 1.250 1.125 1.420 2.370 ;
        RECT 0.105 2.200 1.420 2.370 ;
        RECT 1.250 1.610 1.990 1.910 ;
  END 
END OR3HDMXHT

MACRO OAI22B2HD2XHT
  CLASS  CORE ;
  FOREIGN OAI22B2HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.245 1.280 1.730 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.530 1.245 1.950 1.730 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.500 1.330 2.855 1.730 ;
        RECT 2.500 1.560 3.550 1.730 ;
    END
  END D
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.570 0.390 2.015 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.150 -0.300 1.450 1.055 ;
        RECT 2.230 -0.300 2.530 0.715 ;
        RECT 3.270 -0.300 3.570 0.715 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.750 2.635 3.050 3.145 ;
        RECT 3.790 2.285 4.090 3.145 ;
        RECT 2.750 2.975 4.090 3.145 ;
        RECT 4.310 1.125 5.065 1.295 ;
        RECT 3.790 2.285 5.065 2.455 ;
        RECT 4.895 1.125 5.065 2.620 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.195 2.280 0.365 3.990 ;
        RECT 1.200 2.295 1.500 3.990 ;
        RECT 2.240 2.635 2.540 3.990 ;
        RECT 4.310 2.635 4.610 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.720 2.260 2.020 3.145 ;
        RECT 1.720 2.260 3.570 2.430 ;
        RECT 3.270 2.260 3.570 2.770 ;
        RECT 0.130 1.050 0.740 1.220 ;
        RECT 0.570 1.050 0.740 2.080 ;
        RECT 0.715 1.910 0.885 2.280 ;
        RECT 4.015 1.605 4.185 2.080 ;
        RECT 0.570 1.910 4.185 2.080 ;
        RECT 4.015 1.605 4.705 1.775 ;
        RECT 4.535 1.540 4.705 1.840 ;
        RECT 1.710 0.545 2.010 1.065 ;
        RECT 2.750 0.545 3.050 1.065 ;
        RECT 3.790 0.545 4.090 1.065 ;
        RECT 1.710 0.895 4.090 1.065 ;
        RECT 3.790 0.545 5.065 0.715 ;
        RECT 4.895 0.545 5.065 0.845 ;
  END 
END OAI22B2HD2XHT

MACRO OAI222HDMXHT
  CLASS  CORE ;
  FOREIGN OAI222HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.635 0.310 2.015 ;
        RECT 0.100 1.635 0.585 1.870 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.765 1.635 1.000 2.360 ;
        RECT 0.445 2.150 1.000 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.865 1.650 2.430 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.215 1.635 1.655 1.950 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.655 1.480 3.180 1.780 ;
        RECT 2.970 1.480 3.180 2.420 ;
    END
  END E
  PIN F
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.720 1.680 4.000 2.830 ;
    END
  END F
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.585 -0.300 0.885 0.555 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.210 2.130 1.380 3.180 ;
        RECT 0.860 2.970 1.380 3.180 ;
        RECT 1.210 2.130 2.790 2.300 ;
        RECT 2.620 2.130 2.790 2.775 ;
        RECT 3.175 1.125 3.530 1.295 ;
        RECT 3.360 1.125 3.530 2.775 ;
        RECT 2.620 2.605 3.530 2.775 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.540 0.405 3.990 ;
        RECT 2.140 2.540 2.440 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 1.455 ;
        RECT 1.200 1.060 1.370 1.455 ;
        RECT 2.270 1.060 2.440 1.455 ;
        RECT 0.170 1.285 2.440 1.455 ;
        RECT 1.900 0.640 2.070 1.105 ;
        RECT 1.685 0.935 2.070 1.105 ;
        RECT 1.900 0.640 3.930 0.810 ;
        RECT 3.760 0.640 3.930 1.170 ;
  END 
END OAI222HDMXHT

MACRO OAI221HD2XHT
  CLASS  CORE ;
  FOREIGN OAI221HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.740 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.640 0.310 2.015 ;
        RECT 0.100 1.640 0.585 1.810 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.850 2.665 1.200 3.180 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.875 1.630 2.430 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.215 1.575 1.610 1.950 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.800 1.265 3.180 1.820 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.045 ;
        RECT 4.340 -0.300 4.510 1.060 ;
        RECT 5.315 -0.300 5.615 1.055 ;
        RECT 0.000 -0.300 5.740 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.860 0.720 5.030 2.960 ;
        RECT 4.860 1.235 5.230 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 2.215 2.480 2.855 3.990 ;
        RECT 4.275 2.295 4.575 3.990 ;
        RECT 5.315 2.295 5.615 3.990 ;
        RECT 0.000 3.390 5.740 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.900 0.340 1.395 ;
        RECT 1.210 0.900 1.380 1.395 ;
        RECT 2.280 0.900 2.450 1.395 ;
        RECT 0.170 1.225 2.450 1.395 ;
        RECT 1.910 0.550 2.080 1.045 ;
        RECT 1.695 0.875 2.080 1.045 ;
        RECT 1.910 0.550 2.895 0.720 ;
        RECT 2.725 0.550 2.895 1.045 ;
        RECT 2.725 0.875 3.025 1.045 ;
        RECT 1.210 2.130 1.380 2.430 ;
        RECT 3.310 0.810 3.530 1.110 ;
        RECT 3.105 2.045 3.530 2.300 ;
        RECT 3.360 0.810 3.530 2.300 ;
        RECT 1.210 2.130 3.530 2.300 ;
        RECT 3.360 1.590 4.235 1.760 ;
        RECT 3.790 1.945 3.960 2.280 ;
        RECT 3.820 0.900 3.990 1.410 ;
        RECT 3.820 1.240 4.680 1.410 ;
        RECT 4.510 1.240 4.680 2.115 ;
        RECT 3.790 1.945 4.680 2.115 ;
  END 
END OAI221HD2XHT

MACRO OAI211HD2XHT
  CLASS  CORE ;
  FOREIGN OAI211HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.575 0.310 2.015 ;
        RECT 0.100 1.575 0.520 1.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.830 1.575 1.000 2.360 ;
        RECT 0.445 2.150 1.000 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.215 1.575 1.605 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.135 1.265 2.395 1.865 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.045 ;
        RECT 3.275 -0.300 3.575 1.055 ;
        RECT 4.315 -0.300 4.615 1.055 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.860 0.720 4.030 2.960 ;
        RECT 3.860 1.235 4.410 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.540 0.405 3.990 ;
        RECT 1.695 2.540 1.995 3.990 ;
        RECT 3.275 2.295 3.575 3.990 ;
        RECT 4.315 2.295 4.615 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.900 0.340 1.395 ;
        RECT 1.210 0.900 1.380 1.395 ;
        RECT 0.170 1.225 1.380 1.395 ;
        RECT 1.210 2.130 1.380 2.525 ;
        RECT 1.785 0.895 1.955 2.300 ;
        RECT 1.210 2.130 2.450 2.300 ;
        RECT 2.280 2.130 2.450 2.775 ;
        RECT 1.785 0.895 2.745 1.065 ;
        RECT 2.575 0.895 2.745 1.755 ;
        RECT 2.575 1.585 3.205 1.755 ;
        RECT 2.725 0.545 3.095 0.715 ;
        RECT 2.790 1.935 2.960 2.315 ;
        RECT 2.925 0.545 3.095 1.405 ;
        RECT 2.925 1.235 3.650 1.405 ;
        RECT 3.480 1.235 3.650 2.105 ;
        RECT 2.790 1.935 3.650 2.105 ;
  END 
END OAI211HD2XHT

MACRO NOR4B2HDLXHT
  CLASS  CORE ;
  FOREIGN NOR4B2HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.205 0.740 1.615 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.960 1.500 3.130 2.430 ;
        RECT 2.960 2.080 3.185 2.430 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.310 1.360 3.655 1.950 ;
    END
  END D
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.030 1.205 1.540 1.615 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.025 ;
        RECT 1.575 -0.300 1.875 0.545 ;
        RECT 2.595 -0.300 2.895 0.435 ;
        RECT 3.695 -0.300 3.995 0.685 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.125 0.865 4.005 1.035 ;
        RECT 3.835 0.865 4.005 2.840 ;
        RECT 3.645 2.155 4.005 2.840 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.165 0.925 3.990 ;
        RECT 1.655 2.495 1.955 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.090 0.855 0.260 1.965 ;
        RECT 0.170 1.795 0.340 2.280 ;
        RECT 0.090 0.855 0.405 1.025 ;
        RECT 1.835 1.585 2.005 1.965 ;
        RECT 0.090 1.795 2.005 1.965 ;
        RECT 1.835 1.585 2.135 1.755 ;
        RECT 1.145 0.855 1.920 1.025 ;
        RECT 1.750 0.855 1.920 1.405 ;
        RECT 1.750 1.235 2.635 1.405 ;
        RECT 2.465 1.235 2.635 2.315 ;
        RECT 1.145 2.145 2.635 2.315 ;
  END 
END NOR4B2HDLXHT

MACRO NOR4B1HD1XHT
  CLASS  CORE ;
  FOREIGN NOR4B1HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.380 1.565 1.680 2.360 ;
        RECT 1.260 2.150 1.680 2.360 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.215 0.850 1.620 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.990 1.565 2.225 2.770 ;
        RECT 1.670 2.560 2.225 2.770 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.470 1.565 2.640 3.180 ;
        RECT 2.470 2.970 2.840 3.180 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.035 ;
        RECT 1.665 -0.300 1.965 1.035 ;
        RECT 2.705 -0.300 3.005 1.035 ;
        RECT 3.885 -0.300 4.185 0.715 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.470 0.720 4.640 2.960 ;
        RECT 4.470 1.670 4.820 2.020 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.155 0.955 3.990 ;
        RECT 3.885 2.295 4.185 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.090 1.800 0.340 1.975 ;
        RECT 0.090 0.865 0.260 1.975 ;
        RECT 0.170 1.800 0.340 2.280 ;
        RECT 0.090 0.865 0.405 1.035 ;
        RECT 1.030 1.590 1.200 1.970 ;
        RECT 0.090 1.800 1.200 1.970 ;
        RECT 1.210 0.800 1.380 1.385 ;
        RECT 2.250 0.800 2.420 1.385 ;
        RECT 1.210 1.215 2.990 1.385 ;
        RECT 2.820 1.215 2.990 2.620 ;
        RECT 2.820 1.530 3.720 1.730 ;
        RECT 3.400 1.945 3.570 2.280 ;
        RECT 3.335 1.125 4.290 1.295 ;
        RECT 4.120 1.125 4.290 2.115 ;
        RECT 3.400 1.945 4.290 2.115 ;
  END 
END NOR4B1HD1XHT

MACRO NOR2HD2XSPGHT
  CLASS  CORE ;
  FOREIGN NOR2HD2XSPGHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 0.345 0.300 0.885 3.075 ;
      LAYER V7 ;
        RECT 0.435 0.845 0.795 1.205 ;
      LAYER M7 ;
        RECT 0.345 0.835 1.160 1.215 ;
      LAYER V6 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M4 ;
        RECT 0.925 0.835 1.125 1.620 ;
      LAYER V3 ;
        RECT 0.930 1.340 1.120 1.530 ;
      LAYER M3 ;
        RECT 0.405 1.335 1.210 1.535 ;
      LAYER V2 ;
        RECT 0.520 1.340 0.710 1.530 ;
      LAYER M2 ;
        RECT 0.515 1.220 0.715 2.030 ;
      LAYER V1 ;
        RECT 0.520 1.750 0.710 1.940 ;
      LAYER M1 ;
        RECT 0.430 1.540 1.385 1.950 ;
        RECT 1.215 1.540 1.385 3.170 ;
        RECT 2.130 2.130 2.300 3.170 ;
        RECT 1.215 3.000 2.300 3.170 ;
        RECT 2.830 1.610 3.000 2.300 ;
        RECT 2.130 2.130 3.000 2.300 ;
      LAYER M6 ;
        RECT 0.515 0.300 0.715 2.160 ;
      LAYER V5 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M5 ;
        RECT 0.345 0.925 1.240 1.125 ;
      LAYER V4 ;
        RECT 0.930 0.930 1.120 1.120 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 2.805 0.300 3.345 3.075 ;
      LAYER V7 ;
        RECT 2.895 0.845 3.255 1.205 ;
      LAYER M7 ;
        RECT 2.565 0.835 3.345 1.215 ;
      LAYER V6 ;
        RECT 2.980 0.930 3.170 1.120 ;
      LAYER M4 ;
        RECT 2.565 0.835 2.765 1.700 ;
      LAYER V3 ;
        RECT 2.570 1.340 2.760 1.530 ;
      LAYER M3 ;
        RECT 1.895 1.335 2.850 1.535 ;
      LAYER V2 ;
        RECT 2.160 1.340 2.350 1.530 ;
      LAYER M2 ;
        RECT 2.155 1.200 2.355 2.050 ;
      LAYER V1 ;
        RECT 2.160 1.750 2.350 1.940 ;
      LAYER M1 ;
        RECT 1.915 1.540 2.430 1.950 ;
      LAYER M6 ;
        RECT 2.975 0.300 3.175 2.160 ;
      LAYER V5 ;
        RECT 2.980 0.930 3.170 1.120 ;
      LAYER M5 ;
        RECT 2.565 0.835 3.345 1.215 ;
      LAYER V4 ;
        RECT 2.570 0.930 2.760 1.120 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 -0.300 0.895 1.035 ;
        RECT 1.710 -0.300 2.010 0.875 ;
        RECT 2.835 -0.300 3.135 0.435 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 1.575 0.300 2.115 3.075 ;
      LAYER V7 ;
        RECT 1.665 0.845 2.025 1.205 ;
      LAYER M7 ;
        RECT 1.575 0.835 2.355 1.215 ;
      LAYER V6 ;
        RECT 1.750 0.930 1.940 1.120 ;
      LAYER M4 ;
        RECT 2.155 0.835 2.355 2.450 ;
      LAYER V3 ;
        RECT 2.160 2.160 2.350 2.350 ;
      LAYER M3 ;
        RECT 1.495 2.155 2.450 2.355 ;
      LAYER V2 ;
        RECT 1.750 2.160 1.940 2.350 ;
      LAYER M2 ;
        RECT 1.745 2.050 1.945 2.820 ;
      LAYER V1 ;
        RECT 1.750 2.405 1.940 2.595 ;
      LAYER M1 ;
        RECT 1.210 0.890 1.380 1.360 ;
        RECT 1.565 1.190 1.735 2.820 ;
        RECT 1.565 2.180 1.950 2.820 ;
        RECT 2.340 0.890 2.510 1.360 ;
        RECT 1.210 1.190 2.510 1.360 ;
      LAYER M6 ;
        RECT 1.745 0.300 1.945 2.160 ;
      LAYER V5 ;
        RECT 1.750 0.930 1.940 1.120 ;
      LAYER M5 ;
        RECT 1.575 0.835 2.355 1.215 ;
      LAYER V4 ;
        RECT 2.160 0.930 2.350 1.120 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.800 2.230 1.035 3.990 ;
        RECT 2.600 2.635 2.900 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
END NOR2HD2XSPGHT

MACRO NOR2B1HD1XHT
  CLASS  CORE ;
  FOREIGN NOR2B1HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.305 1.565 1.570 2.030 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.500 0.520 2.015 ;
    END
  END AN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.570 -0.300 0.870 0.745 ;
        RECT 1.640 -0.300 1.940 0.955 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.185 0.720 1.355 1.385 ;
        RECT 1.185 1.215 1.950 1.385 ;
        RECT 1.780 1.215 1.950 3.210 ;
        RECT 1.705 2.230 1.950 3.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.675 2.635 0.975 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 1.005 1.295 ;
        RECT 0.835 1.125 1.005 2.365 ;
        RECT 0.105 2.195 1.005 2.365 ;
        RECT 0.835 1.540 1.090 1.840 ;
  END 
END NOR2B1HD1XHT

MACRO NAND4B1HDMXHT
  CLASS  CORE ;
  FOREIGN NAND4B1HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.235 2.560 1.475 2.980 ;
        RECT 1.235 2.560 1.610 2.770 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.510 2.905 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.670 1.330 2.020 1.750 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.245 1.590 2.770 1.760 ;
        RECT 2.560 1.590 2.770 2.020 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.745 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.275 0.920 1.455 2.215 ;
        RECT 1.085 2.045 2.365 2.215 ;
        RECT 1.275 0.920 2.660 1.130 ;
        RECT 2.490 0.720 2.660 1.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.740 2.860 0.910 3.990 ;
        RECT 1.735 2.925 2.035 3.990 ;
        RECT 2.585 2.375 2.885 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.085 1.755 ;
  END 
END NAND4B1HDMXHT

MACRO NAND3B1HD2XHT
  CLASS  CORE ;
  FOREIGN NAND3B1HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.510 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 1.170 1.560 1.820 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.510 2.905 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 0.855 1.955 1.820 ;
        RECT 1.740 1.520 2.040 1.820 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 3.055 -0.300 3.355 1.055 ;
        RECT 4.095 -0.300 4.395 1.055 ;
        RECT 0.000 -0.300 4.510 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.640 0.720 3.810 2.965 ;
        RECT 3.640 1.740 4.090 1.950 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 1.980 0.860 3.990 ;
        RECT 1.635 2.625 1.935 3.990 ;
        RECT 3.055 2.295 3.355 3.990 ;
        RECT 4.095 2.295 4.395 3.990 ;
        RECT 0.000 3.390 4.510 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.100 1.755 ;
        RECT 1.120 2.045 1.290 2.845 ;
        RECT 2.150 1.060 2.425 1.360 ;
        RECT 2.255 1.060 2.425 2.215 ;
        RECT 1.120 2.045 2.425 2.215 ;
        RECT 2.255 1.585 2.985 1.755 ;
        RECT 2.475 0.620 2.815 0.790 ;
        RECT 2.645 0.620 2.815 1.405 ;
        RECT 2.705 1.935 2.875 2.735 ;
        RECT 2.505 2.565 2.875 2.735 ;
        RECT 2.645 1.235 3.385 1.405 ;
        RECT 3.215 1.235 3.385 2.105 ;
        RECT 2.705 1.935 3.385 2.105 ;
        RECT 3.215 1.520 3.430 1.820 ;
  END 
END NAND3B1HD2XHT

MACRO NAND2B1HD1XHT
  CLASS  CORE ;
  FOREIGN NAND2B1HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.305 1.260 1.560 1.820 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.495 0.315 2.835 ;
        RECT 0.100 2.495 0.585 2.705 ;
    END
  END AN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.645 -0.300 0.945 0.715 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.605 0.935 1.950 1.055 ;
        RECT 1.150 2.000 1.320 2.980 ;
        RECT 1.740 0.480 1.905 2.170 ;
        RECT 1.605 0.480 1.905 1.055 ;
        RECT 1.740 0.935 1.950 2.170 ;
        RECT 1.150 2.000 1.950 2.170 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 2.905 0.835 3.990 ;
        RECT 1.605 2.465 1.905 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.125 1.755 ;
  END 
END NAND2B1HD1XHT

MACRO MUX2CLKHD1XHT
  CLASS  CORE ;
  FOREIGN MUX2CLKHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.265 1.180 2.020 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.675 2.360 2.430 ;
        RECT 2.150 1.675 2.555 1.910 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.065 ;
        RECT 2.500 -0.300 2.670 1.130 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.900 0.895 3.370 1.130 ;
        RECT 3.170 0.895 3.370 2.960 ;
        RECT 3.050 1.980 3.370 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.555 0.955 3.990 ;
        RECT 2.465 2.635 2.765 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.260 0.720 1.950 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.090 0.895 0.260 2.370 ;
        RECT 0.090 0.895 0.405 1.065 ;
        RECT 0.090 2.175 0.405 2.370 ;
        RECT 1.430 1.330 1.600 2.370 ;
        RECT 0.090 2.200 1.600 2.370 ;
        RECT 1.545 0.895 1.950 1.065 ;
        RECT 1.780 0.895 1.950 2.725 ;
        RECT 1.545 2.555 1.950 2.725 ;
        RECT 1.780 1.325 2.970 1.495 ;
        RECT 2.735 1.325 2.970 1.670 ;
  END 
END MUX2CLKHD1XHT

MACRO INVHDMXHT
  CLASS  CORE ;
  FOREIGN INVHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.230 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.310 2.015 ;
        RECT 0.100 1.520 0.600 1.820 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.195 -0.300 0.495 1.145 ;
        RECT 0.000 -0.300 1.230 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.780 1.060 0.950 2.280 ;
        RECT 0.780 1.265 1.130 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.195 2.375 0.495 3.990 ;
        RECT 0.000 3.390 1.230 3.990 ;
    END
  END VDD
END INVHDMXHT

MACRO INVHD8XHT
  CLASS  CORE ;
  FOREIGN INVHD8XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.425 1.610 0.800 1.950 ;
        RECT 0.425 1.610 2.565 1.780 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.225 -0.300 0.525 1.055 ;
        RECT 1.265 -0.300 1.565 0.715 ;
        RECT 2.305 -0.300 2.605 0.715 ;
        RECT 3.345 -0.300 3.645 0.715 ;
        RECT 4.385 -0.300 4.685 1.055 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.745 0.785 1.045 1.360 ;
        RECT 0.745 2.140 1.050 3.055 ;
        RECT 1.785 0.785 2.085 1.360 ;
        RECT 1.785 2.140 2.085 3.055 ;
        RECT 0.745 0.940 4.165 1.360 ;
        RECT 2.855 0.785 3.125 3.055 ;
        RECT 2.825 0.785 3.125 1.360 ;
        RECT 2.855 0.940 3.130 3.055 ;
        RECT 2.825 2.140 3.130 3.055 ;
        RECT 2.855 0.940 4.165 2.410 ;
        RECT 0.745 2.140 4.165 2.410 ;
        RECT 3.865 0.785 4.165 3.055 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.225 2.295 0.525 3.990 ;
        RECT 1.265 2.635 1.565 3.990 ;
        RECT 2.305 2.635 2.605 3.990 ;
        RECT 3.345 2.635 3.645 3.990 ;
        RECT 4.385 2.295 4.685 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
END INVHD8XHT

MACRO INVHD1XSPGHT
  CLASS  CORE ;
  FOREIGN INVHD1XSPGHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 0.345 0.425 0.885 3.070 ;
      LAYER V7 ;
        RECT 0.435 0.845 0.795 1.205 ;
      LAYER M7 ;
        RECT 0.195 0.835 0.965 1.215 ;
      LAYER V6 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M4 ;
        RECT 0.515 0.825 0.715 1.620 ;
      LAYER V3 ;
        RECT 0.520 1.340 0.710 1.530 ;
      LAYER M3 ;
        RECT 0.105 1.250 0.720 1.620 ;
      LAYER V2 ;
        RECT 0.110 1.340 0.300 1.530 ;
      LAYER M2 ;
        RECT 0.105 1.240 0.305 2.015 ;
      LAYER V1 ;
        RECT 0.110 1.750 0.300 1.940 ;
      LAYER M1 ;
        RECT 0.100 1.520 0.310 2.015 ;
        RECT 0.100 1.520 1.200 1.820 ;
      LAYER M6 ;
        RECT 0.515 0.425 0.715 1.855 ;
      LAYER V5 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M5 ;
        RECT 0.195 0.925 0.965 1.125 ;
      LAYER V4 ;
        RECT 0.520 0.930 0.710 1.120 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.805 -0.300 1.105 1.120 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 1.575 0.325 2.115 3.065 ;
      LAYER V7 ;
        RECT 1.665 0.435 2.025 0.795 ;
      LAYER M7 ;
        RECT 1.390 0.425 2.115 0.805 ;
      LAYER V6 ;
        RECT 1.750 0.520 1.940 0.710 ;
      LAYER M4 ;
        RECT 1.745 0.430 1.945 1.210 ;
      LAYER V3 ;
        RECT 1.750 0.930 1.940 1.120 ;
      LAYER M3 ;
        RECT 1.310 0.840 2.105 1.210 ;
      LAYER V2 ;
        RECT 1.750 0.930 1.940 1.120 ;
      LAYER M2 ;
        RECT 1.745 0.840 1.945 1.670 ;
      LAYER V1 ;
        RECT 1.750 1.340 1.940 1.530 ;
      LAYER M1 ;
        RECT 1.385 0.720 1.575 2.960 ;
        RECT 1.385 1.265 1.950 1.605 ;
      LAYER M6 ;
        RECT 1.745 0.325 1.945 1.855 ;
      LAYER V5 ;
        RECT 1.750 0.520 1.940 0.710 ;
      LAYER M5 ;
        RECT 1.390 0.515 2.115 0.715 ;
      LAYER V4 ;
        RECT 1.750 0.520 1.940 0.710 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.805 2.230 1.105 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
END INVHD1XSPGHT

MACRO INVCLKHD5XHT
  CLASS  CORE ;
  FOREIGN INVCLKHD5XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.445 1.645 0.790 1.950 ;
        RECT 0.445 1.645 1.425 1.815 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.180 ;
        RECT 1.145 -0.300 1.445 1.115 ;
        RECT 2.185 -0.300 2.485 1.115 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.625 1.060 0.925 1.465 ;
        RECT 0.625 2.130 0.925 3.120 ;
        RECT 1.665 1.060 1.965 1.465 ;
        RECT 0.625 1.295 3.005 1.465 ;
        RECT 1.765 1.060 1.965 3.120 ;
        RECT 1.665 2.130 1.965 3.120 ;
        RECT 1.765 1.295 3.005 2.365 ;
        RECT 0.625 2.130 3.005 2.365 ;
        RECT 2.705 1.060 3.005 3.120 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.140 0.405 3.990 ;
        RECT 1.145 2.545 1.445 3.990 ;
        RECT 2.185 2.545 2.485 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
END INVCLKHD5XHT

MACRO INVCLKHD3XHT
  CLASS  CORE ;
  FOREIGN INVCLKHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.430 1.585 0.820 1.950 ;
        RECT 0.430 1.585 1.595 1.760 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.275 -0.300 0.575 0.960 ;
        RECT 1.315 -0.300 1.615 0.960 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.795 1.010 1.095 1.385 ;
        RECT 0.795 2.190 1.095 3.105 ;
        RECT 0.795 1.205 2.135 1.385 ;
        RECT 0.795 2.190 2.135 2.410 ;
        RECT 1.835 1.010 2.135 1.385 ;
        RECT 0.795 1.255 2.360 1.385 ;
        RECT 1.840 1.010 2.135 2.895 ;
        RECT 1.835 2.190 2.135 2.895 ;
        RECT 1.840 1.255 2.360 1.610 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.275 2.295 0.575 3.990 ;
        RECT 1.315 2.635 1.615 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
END INVCLKHD3XHT

MACRO INVCLKHD12XHT
  CLASS  CORE ;
  FOREIGN INVCLKHD12XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.740 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.210 1.675 0.800 1.955 ;
        RECT 0.210 1.675 3.195 1.845 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.020 ;
        RECT 1.145 -0.300 1.445 1.020 ;
        RECT 2.185 -0.300 2.485 1.020 ;
        RECT 3.225 -0.300 3.525 1.020 ;
        RECT 4.265 -0.300 4.565 1.020 ;
        RECT 5.305 -0.300 5.605 1.020 ;
        RECT 0.000 -0.300 5.740 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.625 1.060 0.925 1.495 ;
        RECT 0.625 2.145 0.925 2.995 ;
        RECT 1.665 1.060 1.965 1.495 ;
        RECT 1.665 2.145 1.965 2.995 ;
        RECT 2.705 1.060 3.005 1.495 ;
        RECT 2.705 2.145 3.005 2.995 ;
        RECT 0.625 1.205 5.515 1.495 ;
        RECT 3.745 1.060 4.045 2.895 ;
        RECT 4.785 1.060 5.085 2.895 ;
        RECT 3.690 1.205 5.515 2.410 ;
        RECT 0.625 2.145 5.515 2.410 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 1.145 2.635 1.445 3.990 ;
        RECT 2.185 2.635 2.485 3.990 ;
        RECT 3.225 2.635 3.525 3.990 ;
        RECT 4.265 2.635 4.565 3.990 ;
        RECT 5.305 2.635 5.605 3.990 ;
        RECT 0.000 3.390 5.740 3.990 ;
    END
  END VDD
END INVCLKHD12XHT

MACRO FILLERC2HDHT
  CLASS  CORE ;
  FOREIGN FILLERC2HDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.820 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 -0.300 0.820 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 3.390 0.820 3.990 ;
    END
  END VDD
END FILLERC2HDHT

MACRO FILLER64HDHT
  CLASS  CORE ;
  FOREIGN FILLER64HDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.240 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 -0.300 26.240 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 3.390 26.240 3.990 ;
    END
  END VDD
END FILLER64HDHT

MACRO FILLER32HDHT
  CLASS  CORE ;
  FOREIGN FILLER32HDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.120 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 -0.300 13.120 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 3.390 13.120 3.990 ;
    END
  END VDD
END FILLER32HDHT

MACRO FFSEDHQHDMXHT
  CLASS  CORE ;
  FOREIGN FFSEDHQHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.990 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 15.650 0.720 15.895 2.455 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 1.325 1.220 1.920 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.625 0.620 2.010 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.905 1.545 3.205 2.020 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.775 -0.300 1.075 0.775 ;
        RECT 2.560 -0.300 2.880 0.570 ;
        RECT 3.640 -0.300 3.960 0.570 ;
        RECT 5.410 -0.300 5.710 0.570 ;
        RECT 7.040 -0.300 7.340 0.520 ;
        RECT 7.975 -0.300 8.275 0.520 ;
        RECT 9.370 -0.300 9.540 0.820 ;
        RECT 11.175 -0.300 11.475 0.525 ;
        RECT 12.185 -0.300 12.505 0.565 ;
        RECT 14.095 -0.300 14.395 0.695 ;
        RECT 15.020 -0.300 15.320 0.620 ;
        RECT 0.000 -0.300 15.990 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 6.485 1.525 6.935 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.805 1.465 6.130 2.010 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.775 2.640 1.085 3.990 ;
        RECT 2.655 2.910 2.955 3.990 ;
        RECT 3.520 2.910 3.820 3.990 ;
        RECT 5.460 2.890 5.760 3.990 ;
        RECT 7.070 2.890 7.710 3.990 ;
        RECT 9.340 2.535 9.510 3.990 ;
        RECT 11.390 3.160 12.370 3.990 ;
        RECT 14.105 2.830 14.405 3.990 ;
        RECT 15.035 2.865 15.335 3.990 ;
        RECT 0.000 3.390 15.990 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.270 0.975 0.440 1.345 ;
        RECT 0.270 0.975 1.600 1.145 ;
        RECT 1.430 0.975 1.600 2.375 ;
        RECT 0.205 2.205 1.600 2.375 ;
        RECT 1.430 1.705 1.700 2.005 ;
        RECT 1.780 1.045 2.050 1.345 ;
        RECT 1.880 1.045 2.050 2.730 ;
        RECT 1.780 2.375 2.050 2.730 ;
        RECT 3.805 1.775 3.975 2.730 ;
        RECT 1.780 2.550 3.975 2.730 ;
        RECT 3.430 1.110 3.600 2.370 ;
        RECT 3.130 2.200 3.600 2.370 ;
        RECT 3.130 1.110 4.290 1.280 ;
        RECT 4.120 1.110 4.290 1.650 ;
        RECT 4.165 1.480 4.335 3.190 ;
        RECT 4.120 1.480 4.520 1.650 ;
        RECT 4.165 3.020 5.020 3.190 ;
        RECT 5.245 1.110 5.415 2.360 ;
        RECT 5.245 1.110 6.280 1.280 ;
        RECT 5.245 2.190 6.280 2.360 ;
        RECT 6.490 1.125 7.285 1.295 ;
        RECT 7.115 1.125 7.285 2.360 ;
        RECT 6.490 2.190 7.285 2.360 ;
        RECT 7.115 1.525 7.415 1.825 ;
        RECT 7.595 1.125 7.765 2.215 ;
        RECT 7.530 1.125 7.830 1.295 ;
        RECT 7.570 2.045 8.540 2.215 ;
        RECT 8.370 2.045 8.540 2.630 ;
        RECT 8.370 2.460 9.000 2.630 ;
        RECT 4.515 1.890 4.685 2.710 ;
        RECT 4.470 1.110 4.870 1.280 ;
        RECT 4.700 1.110 4.870 2.070 ;
        RECT 4.515 1.890 4.870 2.070 ;
        RECT 4.515 2.540 8.185 2.710 ;
        RECT 8.015 2.540 8.185 3.080 ;
        RECT 8.015 2.910 9.140 3.080 ;
        RECT 8.970 2.910 9.140 3.210 ;
        RECT 10.410 0.955 10.580 2.280 ;
        RECT 10.345 0.955 10.645 1.125 ;
        RECT 10.410 1.675 11.845 1.845 ;
        RECT 11.755 1.125 12.055 1.495 ;
        RECT 11.065 1.325 12.615 1.495 ;
        RECT 12.445 1.325 12.615 2.215 ;
        RECT 11.725 2.045 12.615 2.215 ;
        RECT 8.565 1.125 8.890 1.295 ;
        RECT 8.720 1.125 8.890 2.260 ;
        RECT 8.720 2.090 9.860 2.260 ;
        RECT 9.690 2.090 9.860 2.980 ;
        RECT 9.690 2.810 13.195 2.980 ;
        RECT 12.895 2.810 13.195 3.195 ;
        RECT 9.090 1.455 10.210 1.625 ;
        RECT 10.040 1.455 10.210 2.630 ;
        RECT 12.795 1.310 12.965 2.630 ;
        RECT 12.795 1.310 13.195 1.480 ;
        RECT 10.040 2.460 13.650 2.630 ;
        RECT 13.480 2.460 13.650 2.945 ;
        RECT 2.460 0.750 2.630 1.825 ;
        RECT 2.460 0.750 7.870 0.930 ;
        RECT 2.460 0.750 8.950 0.920 ;
        RECT 9.855 0.605 10.025 1.200 ;
        RECT 9.310 1.030 10.025 1.200 ;
        RECT 9.855 0.605 10.860 0.775 ;
        RECT 11.155 0.765 12.805 0.945 ;
        RECT 13.065 0.575 13.630 0.760 ;
        RECT 14.005 0.935 14.135 1.480 ;
        RECT 14.005 0.935 15.025 1.110 ;
        RECT 14.855 0.935 15.025 2.215 ;
        RECT 14.645 2.045 15.025 2.215 ;
        RECT 13.835 0.715 13.845 1.479 ;
        RECT 13.845 0.725 13.855 1.479 ;
        RECT 13.855 0.735 13.865 1.479 ;
        RECT 13.865 0.745 13.875 1.479 ;
        RECT 13.875 0.755 13.885 1.479 ;
        RECT 13.885 0.765 13.895 1.479 ;
        RECT 13.895 0.775 13.905 1.479 ;
        RECT 13.905 0.785 13.915 1.479 ;
        RECT 13.915 0.795 13.925 1.479 ;
        RECT 13.925 0.805 13.935 1.479 ;
        RECT 13.935 0.815 13.945 1.479 ;
        RECT 13.945 0.825 13.955 1.479 ;
        RECT 13.955 0.835 13.965 1.479 ;
        RECT 13.965 0.845 13.975 1.479 ;
        RECT 13.975 0.855 13.985 1.479 ;
        RECT 13.985 0.865 13.995 1.479 ;
        RECT 13.995 0.875 14.005 1.479 ;
        RECT 13.705 0.585 13.715 0.835 ;
        RECT 13.715 0.595 13.725 0.845 ;
        RECT 13.725 0.605 13.735 0.855 ;
        RECT 13.735 0.615 13.745 0.865 ;
        RECT 13.745 0.625 13.755 0.875 ;
        RECT 13.755 0.635 13.765 0.885 ;
        RECT 13.765 0.645 13.775 0.895 ;
        RECT 13.775 0.655 13.785 0.905 ;
        RECT 13.785 0.665 13.795 0.915 ;
        RECT 13.795 0.675 13.805 0.925 ;
        RECT 13.805 0.685 13.815 0.935 ;
        RECT 13.815 0.695 13.825 0.945 ;
        RECT 13.825 0.705 13.835 0.955 ;
        RECT 13.630 0.575 13.640 0.759 ;
        RECT 13.640 0.575 13.650 0.769 ;
        RECT 13.650 0.575 13.660 0.779 ;
        RECT 13.660 0.575 13.670 0.789 ;
        RECT 13.670 0.575 13.680 0.799 ;
        RECT 13.680 0.575 13.690 0.809 ;
        RECT 13.690 0.575 13.700 0.819 ;
        RECT 13.700 0.575 13.706 0.829 ;
        RECT 12.995 0.575 13.005 0.819 ;
        RECT 13.005 0.575 13.015 0.809 ;
        RECT 13.015 0.575 13.025 0.799 ;
        RECT 13.025 0.575 13.035 0.789 ;
        RECT 13.035 0.575 13.045 0.779 ;
        RECT 13.045 0.575 13.055 0.769 ;
        RECT 13.055 0.575 13.065 0.759 ;
        RECT 12.880 0.690 12.890 0.934 ;
        RECT 12.890 0.680 12.900 0.924 ;
        RECT 12.900 0.670 12.910 0.914 ;
        RECT 12.910 0.660 12.920 0.904 ;
        RECT 12.920 0.650 12.930 0.894 ;
        RECT 12.930 0.640 12.940 0.884 ;
        RECT 12.940 0.630 12.950 0.874 ;
        RECT 12.950 0.620 12.960 0.864 ;
        RECT 12.960 0.610 12.970 0.854 ;
        RECT 12.970 0.600 12.980 0.844 ;
        RECT 12.980 0.590 12.990 0.834 ;
        RECT 12.990 0.580 12.996 0.830 ;
        RECT 12.805 0.765 12.815 0.945 ;
        RECT 12.815 0.755 12.825 0.945 ;
        RECT 12.825 0.745 12.835 0.945 ;
        RECT 12.835 0.735 12.845 0.945 ;
        RECT 12.845 0.725 12.855 0.945 ;
        RECT 12.855 0.715 12.865 0.945 ;
        RECT 12.865 0.705 12.875 0.945 ;
        RECT 12.875 0.695 12.881 0.945 ;
        RECT 11.030 0.650 11.040 0.944 ;
        RECT 11.040 0.660 11.050 0.944 ;
        RECT 11.050 0.670 11.060 0.944 ;
        RECT 11.060 0.680 11.070 0.944 ;
        RECT 11.070 0.690 11.080 0.944 ;
        RECT 11.080 0.700 11.090 0.944 ;
        RECT 11.090 0.710 11.100 0.944 ;
        RECT 11.100 0.720 11.110 0.944 ;
        RECT 11.110 0.730 11.120 0.944 ;
        RECT 11.120 0.740 11.130 0.944 ;
        RECT 11.130 0.750 11.140 0.944 ;
        RECT 11.140 0.760 11.150 0.944 ;
        RECT 11.150 0.765 11.156 0.945 ;
        RECT 10.995 0.615 11.005 0.909 ;
        RECT 11.005 0.625 11.015 0.919 ;
        RECT 11.015 0.635 11.025 0.929 ;
        RECT 11.025 0.640 11.031 0.940 ;
        RECT 10.860 0.605 10.870 0.775 ;
        RECT 10.870 0.605 10.880 0.785 ;
        RECT 10.880 0.605 10.890 0.795 ;
        RECT 10.890 0.605 10.900 0.805 ;
        RECT 10.900 0.605 10.910 0.815 ;
        RECT 10.910 0.605 10.920 0.825 ;
        RECT 10.920 0.605 10.930 0.835 ;
        RECT 10.930 0.605 10.940 0.845 ;
        RECT 10.940 0.605 10.950 0.855 ;
        RECT 10.950 0.605 10.960 0.865 ;
        RECT 10.960 0.605 10.970 0.875 ;
        RECT 10.970 0.605 10.980 0.885 ;
        RECT 10.980 0.605 10.990 0.895 ;
        RECT 10.990 0.605 10.996 0.905 ;
        RECT 9.230 0.960 9.240 1.200 ;
        RECT 9.240 0.970 9.250 1.200 ;
        RECT 9.250 0.980 9.260 1.200 ;
        RECT 9.260 0.990 9.270 1.200 ;
        RECT 9.270 1.000 9.280 1.200 ;
        RECT 9.280 1.010 9.290 1.200 ;
        RECT 9.290 1.020 9.300 1.200 ;
        RECT 9.300 1.030 9.310 1.200 ;
        RECT 9.030 0.760 9.040 1.000 ;
        RECT 9.040 0.770 9.050 1.010 ;
        RECT 9.050 0.780 9.060 1.020 ;
        RECT 9.060 0.790 9.070 1.030 ;
        RECT 9.070 0.800 9.080 1.040 ;
        RECT 9.080 0.810 9.090 1.050 ;
        RECT 9.090 0.820 9.100 1.060 ;
        RECT 9.100 0.830 9.110 1.070 ;
        RECT 9.110 0.840 9.120 1.080 ;
        RECT 9.120 0.850 9.130 1.090 ;
        RECT 9.130 0.860 9.140 1.100 ;
        RECT 9.140 0.870 9.150 1.110 ;
        RECT 9.150 0.880 9.160 1.120 ;
        RECT 9.160 0.890 9.170 1.130 ;
        RECT 9.170 0.900 9.180 1.140 ;
        RECT 9.180 0.910 9.190 1.150 ;
        RECT 9.190 0.920 9.200 1.160 ;
        RECT 9.200 0.930 9.210 1.170 ;
        RECT 9.210 0.940 9.220 1.180 ;
        RECT 9.220 0.950 9.230 1.190 ;
        RECT 8.950 0.750 8.960 0.920 ;
        RECT 8.960 0.750 8.970 0.930 ;
        RECT 8.970 0.750 8.980 0.940 ;
        RECT 8.980 0.750 8.990 0.950 ;
        RECT 8.990 0.750 9.000 0.960 ;
        RECT 9.000 0.750 9.010 0.970 ;
        RECT 9.010 0.750 9.020 0.980 ;
        RECT 9.020 0.750 9.030 0.990 ;
        RECT 13.145 0.940 13.545 1.110 ;
        RECT 13.375 0.940 13.545 2.215 ;
        RECT 13.145 2.045 13.545 2.215 ;
        RECT 14.295 1.675 14.465 2.650 ;
        RECT 14.485 1.540 14.655 1.845 ;
        RECT 13.375 1.675 14.655 1.845 ;
        RECT 15.300 1.520 15.470 2.650 ;
        RECT 14.295 2.480 15.470 2.650 ;
  END 
END FFSEDHQHDMXHT

MACRO FFSEDCRHD2XHT
  CLASS  CORE ;
  FOREIGN FFSEDCRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.630 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 16.770 0.720 16.940 2.960 ;
        RECT 16.770 1.645 17.120 2.035 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 15.680 0.720 15.900 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.040 1.265 2.420 1.795 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 2.560 0.990 2.770 ;
        RECT 0.820 2.560 0.990 3.105 ;
        RECT 0.820 2.935 1.525 3.105 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.620 1.610 2.800 2.430 ;
        RECT 2.560 2.085 2.800 2.430 ;
        RECT 2.620 1.610 3.015 1.780 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.775 1.675 6.955 2.360 ;
        RECT 6.550 2.150 6.955 2.360 ;
        RECT 6.775 1.675 7.095 1.975 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.685 ;
        RECT 2.425 -0.300 2.725 0.745 ;
        RECT 3.470 -0.300 3.770 0.550 ;
        RECT 3.470 -0.300 4.870 0.315 ;
        RECT 4.570 -0.300 4.870 0.550 ;
        RECT 6.640 -0.300 6.940 0.595 ;
        RECT 8.195 -0.300 8.495 0.595 ;
        RECT 11.125 -0.300 11.295 0.585 ;
        RECT 12.190 -0.300 12.360 0.700 ;
        RECT 14.180 -0.300 14.350 1.060 ;
        RECT 15.145 -0.300 15.445 1.055 ;
        RECT 16.185 -0.300 16.485 1.055 ;
        RECT 17.225 -0.300 17.525 1.055 ;
        RECT 0.000 -0.300 17.630 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 7.715 1.530 8.170 1.950 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.170 1.515 6.595 1.950 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.405 2.960 0.640 3.990 ;
        RECT 2.425 2.970 2.725 3.990 ;
        RECT 3.325 2.695 3.625 3.990 ;
        RECT 4.780 2.405 5.080 3.990 ;
        RECT 6.690 2.995 6.990 3.990 ;
        RECT 8.155 2.915 8.455 3.990 ;
        RECT 10.975 3.170 11.275 3.990 ;
        RECT 12.125 3.170 12.425 3.990 ;
        RECT 14.085 2.825 14.385 3.990 ;
        RECT 15.145 2.975 15.445 3.990 ;
        RECT 16.185 2.975 16.485 3.990 ;
        RECT 17.225 2.295 17.525 3.990 ;
        RECT 0.000 3.390 17.630 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.010 0.340 2.300 ;
        RECT 0.170 1.585 1.340 1.755 ;
        RECT 1.170 0.605 1.340 2.755 ;
        RECT 1.170 0.605 1.525 0.775 ;
        RECT 1.170 2.585 1.940 2.755 ;
        RECT 1.770 2.585 1.940 3.170 ;
        RECT 1.520 1.010 1.690 2.405 ;
        RECT 1.520 2.225 2.330 2.405 ;
        RECT 2.160 2.225 2.330 2.780 ;
        RECT 2.160 2.610 3.130 2.780 ;
        RECT 2.960 2.610 3.130 3.080 ;
        RECT 2.900 1.125 3.770 1.295 ;
        RECT 3.600 1.125 3.770 2.300 ;
        RECT 2.980 2.000 3.770 2.300 ;
        RECT 4.020 1.125 4.490 1.295 ;
        RECT 4.310 1.125 4.480 2.505 ;
        RECT 4.310 1.125 4.490 1.945 ;
        RECT 5.025 1.645 5.195 1.945 ;
        RECT 4.310 1.775 5.195 1.945 ;
        RECT 5.490 0.830 5.555 3.085 ;
        RECT 5.580 0.830 5.930 1.000 ;
        RECT 5.490 2.915 6.250 3.085 ;
        RECT 6.315 1.125 7.455 1.295 ;
        RECT 7.285 1.125 7.455 2.415 ;
        RECT 7.135 2.245 7.455 2.415 ;
        RECT 6.225 1.045 6.235 1.295 ;
        RECT 6.235 1.055 6.245 1.295 ;
        RECT 6.245 1.065 6.255 1.295 ;
        RECT 6.255 1.075 6.265 1.295 ;
        RECT 6.265 1.085 6.275 1.295 ;
        RECT 6.275 1.095 6.285 1.295 ;
        RECT 6.285 1.105 6.295 1.295 ;
        RECT 6.295 1.115 6.305 1.295 ;
        RECT 6.305 1.125 6.315 1.295 ;
        RECT 6.020 0.840 6.030 1.090 ;
        RECT 6.030 0.850 6.040 1.100 ;
        RECT 6.040 0.860 6.050 1.110 ;
        RECT 6.050 0.870 6.060 1.120 ;
        RECT 6.060 0.880 6.070 1.130 ;
        RECT 6.070 0.890 6.080 1.140 ;
        RECT 6.080 0.900 6.090 1.150 ;
        RECT 6.090 0.910 6.100 1.160 ;
        RECT 6.100 0.920 6.110 1.170 ;
        RECT 6.110 0.930 6.120 1.180 ;
        RECT 6.120 0.940 6.130 1.190 ;
        RECT 6.130 0.950 6.140 1.200 ;
        RECT 6.140 0.960 6.150 1.210 ;
        RECT 6.150 0.970 6.160 1.220 ;
        RECT 6.160 0.980 6.170 1.230 ;
        RECT 6.170 0.990 6.180 1.240 ;
        RECT 6.180 1.000 6.190 1.250 ;
        RECT 6.190 1.010 6.200 1.260 ;
        RECT 6.200 1.020 6.210 1.270 ;
        RECT 6.210 1.030 6.220 1.280 ;
        RECT 6.220 1.035 6.226 1.289 ;
        RECT 5.930 0.830 5.940 1.000 ;
        RECT 5.940 0.830 5.950 1.010 ;
        RECT 5.950 0.830 5.960 1.020 ;
        RECT 5.960 0.830 5.970 1.030 ;
        RECT 5.970 0.830 5.980 1.040 ;
        RECT 5.980 0.830 5.990 1.050 ;
        RECT 5.990 0.830 6.000 1.060 ;
        RECT 6.000 0.830 6.010 1.070 ;
        RECT 6.010 0.830 6.020 1.080 ;
        RECT 5.555 0.830 5.565 1.014 ;
        RECT 5.565 0.830 5.575 1.004 ;
        RECT 5.575 0.830 5.581 1.000 ;
        RECT 5.385 0.935 5.395 3.085 ;
        RECT 5.395 0.925 5.405 3.085 ;
        RECT 5.405 0.915 5.415 3.085 ;
        RECT 5.415 0.905 5.425 3.085 ;
        RECT 5.425 0.895 5.435 3.085 ;
        RECT 5.435 0.885 5.445 3.085 ;
        RECT 5.445 0.875 5.455 3.085 ;
        RECT 5.455 0.865 5.465 3.085 ;
        RECT 5.465 0.855 5.475 3.085 ;
        RECT 5.475 0.845 5.485 3.085 ;
        RECT 5.485 0.835 5.491 3.085 ;
        RECT 7.645 1.125 8.530 1.295 ;
        RECT 8.350 1.125 8.530 2.335 ;
        RECT 7.645 2.165 8.530 2.335 ;
        RECT 8.350 1.535 8.610 1.835 ;
        RECT 8.790 1.125 8.960 2.365 ;
        RECT 8.730 1.125 9.030 1.295 ;
        RECT 5.735 1.235 5.905 2.735 ;
        RECT 6.350 2.605 7.860 2.745 ;
        RECT 6.360 2.605 7.860 2.755 ;
        RECT 6.370 2.605 7.860 2.765 ;
        RECT 5.735 2.565 6.445 2.735 ;
        RECT 5.735 2.575 6.455 2.735 ;
        RECT 5.735 2.585 6.465 2.735 ;
        RECT 5.735 2.595 6.475 2.735 ;
        RECT 7.670 2.545 7.860 2.775 ;
        RECT 6.380 2.605 7.860 2.775 ;
        RECT 9.240 1.200 9.540 1.370 ;
        RECT 7.670 2.545 9.540 2.715 ;
        RECT 9.370 1.200 9.540 2.715 ;
        RECT 10.070 1.200 10.370 1.370 ;
        RECT 10.200 1.200 10.370 2.290 ;
        RECT 10.070 2.120 10.370 2.290 ;
        RECT 10.200 1.960 11.190 2.130 ;
        RECT 11.310 1.595 11.320 2.089 ;
        RECT 11.320 1.595 11.330 2.079 ;
        RECT 11.330 1.595 11.340 2.069 ;
        RECT 11.340 1.595 11.350 2.059 ;
        RECT 11.350 1.595 11.360 2.049 ;
        RECT 11.360 1.595 11.370 2.039 ;
        RECT 11.370 1.595 11.380 2.029 ;
        RECT 11.380 1.595 11.390 2.019 ;
        RECT 11.390 1.595 11.400 2.009 ;
        RECT 11.400 1.595 11.410 1.999 ;
        RECT 11.410 1.595 11.420 1.989 ;
        RECT 11.420 1.595 11.430 1.979 ;
        RECT 11.430 1.595 11.440 1.969 ;
        RECT 11.440 1.595 11.450 1.959 ;
        RECT 11.450 1.595 11.460 1.949 ;
        RECT 11.460 1.595 11.470 1.939 ;
        RECT 11.470 1.595 11.480 1.929 ;
        RECT 11.480 1.595 11.490 1.919 ;
        RECT 11.490 1.595 11.500 1.909 ;
        RECT 11.280 1.870 11.290 2.120 ;
        RECT 11.290 1.860 11.300 2.110 ;
        RECT 11.300 1.850 11.310 2.100 ;
        RECT 11.190 1.960 11.200 2.130 ;
        RECT 11.200 1.950 11.210 2.130 ;
        RECT 11.210 1.940 11.220 2.130 ;
        RECT 11.220 1.930 11.230 2.130 ;
        RECT 11.230 1.920 11.240 2.130 ;
        RECT 11.240 1.910 11.250 2.130 ;
        RECT 11.250 1.900 11.260 2.130 ;
        RECT 11.260 1.890 11.270 2.130 ;
        RECT 11.270 1.880 11.280 2.130 ;
        RECT 10.915 1.200 11.085 1.740 ;
        RECT 10.785 1.570 11.085 1.740 ;
        RECT 10.915 1.200 11.830 1.370 ;
        RECT 10.915 1.210 11.840 1.370 ;
        RECT 11.680 1.220 11.850 2.290 ;
        RECT 11.550 2.120 11.850 2.290 ;
        RECT 11.680 1.570 12.605 1.740 ;
        RECT 10.250 2.820 12.560 2.990 ;
        RECT 12.870 3.040 13.715 3.210 ;
        RECT 12.780 2.960 12.790 3.210 ;
        RECT 12.790 2.970 12.800 3.210 ;
        RECT 12.800 2.980 12.810 3.210 ;
        RECT 12.810 2.990 12.820 3.210 ;
        RECT 12.820 3.000 12.830 3.210 ;
        RECT 12.830 3.010 12.840 3.210 ;
        RECT 12.840 3.020 12.850 3.210 ;
        RECT 12.850 3.030 12.860 3.210 ;
        RECT 12.860 3.040 12.870 3.210 ;
        RECT 12.650 2.830 12.660 3.080 ;
        RECT 12.660 2.840 12.670 3.090 ;
        RECT 12.670 2.850 12.680 3.100 ;
        RECT 12.680 2.860 12.690 3.110 ;
        RECT 12.690 2.870 12.700 3.120 ;
        RECT 12.700 2.880 12.710 3.130 ;
        RECT 12.710 2.890 12.720 3.140 ;
        RECT 12.720 2.900 12.730 3.150 ;
        RECT 12.730 2.910 12.740 3.160 ;
        RECT 12.740 2.920 12.750 3.170 ;
        RECT 12.750 2.930 12.760 3.180 ;
        RECT 12.760 2.940 12.770 3.190 ;
        RECT 12.770 2.950 12.780 3.200 ;
        RECT 12.560 2.820 12.570 2.990 ;
        RECT 12.570 2.820 12.580 3.000 ;
        RECT 12.580 2.820 12.590 3.010 ;
        RECT 12.590 2.820 12.600 3.020 ;
        RECT 12.600 2.820 12.610 3.030 ;
        RECT 12.610 2.820 12.620 3.040 ;
        RECT 12.620 2.820 12.630 3.050 ;
        RECT 12.630 2.820 12.640 3.060 ;
        RECT 12.640 2.820 12.650 3.070 ;
        RECT 8.775 2.895 9.720 3.065 ;
        RECT 9.890 2.470 10.020 2.760 ;
        RECT 10.015 0.830 10.480 1.000 ;
        RECT 12.785 1.315 12.815 2.640 ;
        RECT 9.890 2.470 12.815 2.640 ;
        RECT 12.905 1.315 12.955 2.730 ;
        RECT 12.905 1.315 13.050 1.615 ;
        RECT 13.035 2.560 13.755 2.730 ;
        RECT 12.955 2.490 12.965 2.730 ;
        RECT 12.965 2.500 12.975 2.730 ;
        RECT 12.975 2.510 12.985 2.730 ;
        RECT 12.985 2.520 12.995 2.730 ;
        RECT 12.995 2.530 13.005 2.730 ;
        RECT 13.005 2.540 13.015 2.730 ;
        RECT 13.015 2.550 13.025 2.730 ;
        RECT 13.025 2.560 13.035 2.730 ;
        RECT 12.815 1.315 12.825 2.639 ;
        RECT 12.825 1.315 12.835 2.649 ;
        RECT 12.835 1.315 12.845 2.659 ;
        RECT 12.845 1.315 12.855 2.669 ;
        RECT 12.855 1.315 12.865 2.679 ;
        RECT 12.865 1.315 12.875 2.689 ;
        RECT 12.875 1.315 12.885 2.699 ;
        RECT 12.885 1.315 12.895 2.709 ;
        RECT 12.895 1.315 12.905 2.719 ;
        RECT 9.940 0.830 9.950 1.064 ;
        RECT 9.950 0.830 9.960 1.054 ;
        RECT 9.960 0.830 9.970 1.044 ;
        RECT 9.970 0.830 9.980 1.034 ;
        RECT 9.980 0.830 9.990 1.024 ;
        RECT 9.990 0.830 10.000 1.014 ;
        RECT 10.000 0.830 10.010 1.004 ;
        RECT 10.010 0.830 10.016 1.000 ;
        RECT 9.890 0.880 9.900 1.114 ;
        RECT 9.900 0.870 9.910 1.104 ;
        RECT 9.910 0.860 9.920 1.094 ;
        RECT 9.920 0.850 9.930 1.084 ;
        RECT 9.930 0.840 9.940 1.074 ;
        RECT 9.720 1.050 9.730 3.064 ;
        RECT 9.730 1.040 9.740 3.064 ;
        RECT 9.740 1.030 9.750 3.064 ;
        RECT 9.750 1.020 9.760 3.064 ;
        RECT 9.760 1.010 9.770 3.064 ;
        RECT 9.770 1.000 9.780 3.064 ;
        RECT 9.780 0.990 9.790 3.064 ;
        RECT 9.790 0.980 9.800 3.064 ;
        RECT 9.800 0.970 9.810 3.064 ;
        RECT 9.810 0.960 9.820 3.064 ;
        RECT 9.820 0.950 9.830 3.064 ;
        RECT 9.830 0.940 9.840 3.064 ;
        RECT 9.840 0.930 9.850 3.064 ;
        RECT 9.850 0.920 9.860 3.064 ;
        RECT 9.860 0.910 9.870 3.064 ;
        RECT 9.870 0.900 9.880 3.064 ;
        RECT 9.880 0.890 9.890 3.064 ;
        RECT 2.990 0.490 3.290 0.945 ;
        RECT 2.990 0.775 4.970 0.945 ;
        RECT 5.400 0.480 6.105 0.650 ;
        RECT 6.490 0.775 9.410 0.945 ;
        RECT 9.790 0.480 10.560 0.650 ;
        RECT 10.985 0.810 11.885 0.980 ;
        RECT 11.965 0.810 11.980 1.060 ;
        RECT 12.705 0.615 12.875 1.060 ;
        RECT 12.050 0.880 12.875 1.060 ;
        RECT 12.705 0.615 13.980 0.785 ;
        RECT 13.810 0.500 13.980 1.410 ;
        RECT 14.700 1.060 14.955 1.410 ;
        RECT 13.810 1.240 14.955 1.410 ;
        RECT 14.785 1.060 14.955 2.285 ;
        RECT 14.635 2.115 14.955 2.285 ;
        RECT 14.785 1.675 15.500 1.845 ;
        RECT 11.980 0.820 11.990 1.060 ;
        RECT 11.990 0.830 12.000 1.060 ;
        RECT 12.000 0.840 12.010 1.060 ;
        RECT 12.010 0.850 12.020 1.060 ;
        RECT 12.020 0.860 12.030 1.060 ;
        RECT 12.030 0.870 12.040 1.060 ;
        RECT 12.040 0.880 12.050 1.060 ;
        RECT 11.885 0.810 11.895 0.980 ;
        RECT 11.895 0.810 11.905 0.990 ;
        RECT 11.905 0.810 11.915 1.000 ;
        RECT 11.915 0.810 11.925 1.010 ;
        RECT 11.925 0.810 11.935 1.020 ;
        RECT 11.935 0.810 11.945 1.030 ;
        RECT 11.945 0.810 11.955 1.040 ;
        RECT 11.955 0.810 11.965 1.050 ;
        RECT 10.890 0.725 10.900 0.979 ;
        RECT 10.900 0.735 10.910 0.979 ;
        RECT 10.910 0.745 10.920 0.979 ;
        RECT 10.920 0.755 10.930 0.979 ;
        RECT 10.930 0.765 10.940 0.979 ;
        RECT 10.940 0.775 10.950 0.979 ;
        RECT 10.950 0.785 10.960 0.979 ;
        RECT 10.960 0.795 10.970 0.979 ;
        RECT 10.970 0.805 10.980 0.979 ;
        RECT 10.980 0.810 10.986 0.980 ;
        RECT 10.655 0.490 10.665 0.744 ;
        RECT 10.665 0.500 10.675 0.754 ;
        RECT 10.675 0.510 10.685 0.764 ;
        RECT 10.685 0.520 10.695 0.774 ;
        RECT 10.695 0.530 10.705 0.784 ;
        RECT 10.705 0.540 10.715 0.794 ;
        RECT 10.715 0.550 10.725 0.804 ;
        RECT 10.725 0.560 10.735 0.814 ;
        RECT 10.735 0.570 10.745 0.824 ;
        RECT 10.745 0.580 10.755 0.834 ;
        RECT 10.755 0.590 10.765 0.844 ;
        RECT 10.765 0.600 10.775 0.854 ;
        RECT 10.775 0.610 10.785 0.864 ;
        RECT 10.785 0.620 10.795 0.874 ;
        RECT 10.795 0.630 10.805 0.884 ;
        RECT 10.805 0.640 10.815 0.894 ;
        RECT 10.815 0.650 10.825 0.904 ;
        RECT 10.825 0.660 10.835 0.914 ;
        RECT 10.835 0.670 10.845 0.924 ;
        RECT 10.845 0.680 10.855 0.934 ;
        RECT 10.855 0.690 10.865 0.944 ;
        RECT 10.865 0.700 10.875 0.954 ;
        RECT 10.875 0.710 10.885 0.964 ;
        RECT 10.885 0.715 10.891 0.975 ;
        RECT 10.560 0.480 10.570 0.650 ;
        RECT 10.570 0.480 10.580 0.660 ;
        RECT 10.580 0.480 10.590 0.670 ;
        RECT 10.590 0.480 10.600 0.680 ;
        RECT 10.600 0.480 10.610 0.690 ;
        RECT 10.610 0.480 10.620 0.700 ;
        RECT 10.620 0.480 10.630 0.710 ;
        RECT 10.630 0.480 10.640 0.720 ;
        RECT 10.640 0.480 10.650 0.730 ;
        RECT 10.650 0.480 10.656 0.740 ;
        RECT 9.705 0.480 9.715 0.724 ;
        RECT 9.715 0.480 9.725 0.714 ;
        RECT 9.725 0.480 9.735 0.704 ;
        RECT 9.735 0.480 9.745 0.694 ;
        RECT 9.745 0.480 9.755 0.684 ;
        RECT 9.755 0.480 9.765 0.674 ;
        RECT 9.765 0.480 9.775 0.664 ;
        RECT 9.775 0.480 9.785 0.654 ;
        RECT 9.785 0.480 9.791 0.650 ;
        RECT 9.495 0.690 9.505 0.934 ;
        RECT 9.505 0.680 9.515 0.924 ;
        RECT 9.515 0.670 9.525 0.914 ;
        RECT 9.525 0.660 9.535 0.904 ;
        RECT 9.535 0.650 9.545 0.894 ;
        RECT 9.545 0.640 9.555 0.884 ;
        RECT 9.555 0.630 9.565 0.874 ;
        RECT 9.565 0.620 9.575 0.864 ;
        RECT 9.575 0.610 9.585 0.854 ;
        RECT 9.585 0.600 9.595 0.844 ;
        RECT 9.595 0.590 9.605 0.834 ;
        RECT 9.605 0.580 9.615 0.824 ;
        RECT 9.615 0.570 9.625 0.814 ;
        RECT 9.625 0.560 9.635 0.804 ;
        RECT 9.635 0.550 9.645 0.794 ;
        RECT 9.645 0.540 9.655 0.784 ;
        RECT 9.655 0.530 9.665 0.774 ;
        RECT 9.665 0.520 9.675 0.764 ;
        RECT 9.675 0.510 9.685 0.754 ;
        RECT 9.685 0.500 9.695 0.744 ;
        RECT 9.695 0.490 9.705 0.734 ;
        RECT 9.410 0.775 9.420 0.945 ;
        RECT 9.420 0.765 9.430 0.945 ;
        RECT 9.430 0.755 9.440 0.945 ;
        RECT 9.440 0.745 9.450 0.945 ;
        RECT 9.450 0.735 9.460 0.945 ;
        RECT 9.460 0.725 9.470 0.945 ;
        RECT 9.470 0.715 9.480 0.945 ;
        RECT 9.480 0.705 9.490 0.945 ;
        RECT 9.490 0.695 9.496 0.945 ;
        RECT 6.400 0.695 6.410 0.945 ;
        RECT 6.410 0.705 6.420 0.945 ;
        RECT 6.420 0.715 6.430 0.945 ;
        RECT 6.430 0.725 6.440 0.945 ;
        RECT 6.440 0.735 6.450 0.945 ;
        RECT 6.450 0.745 6.460 0.945 ;
        RECT 6.460 0.755 6.470 0.945 ;
        RECT 6.470 0.765 6.480 0.945 ;
        RECT 6.480 0.775 6.490 0.945 ;
        RECT 6.195 0.490 6.205 0.740 ;
        RECT 6.205 0.500 6.215 0.750 ;
        RECT 6.215 0.510 6.225 0.760 ;
        RECT 6.225 0.520 6.235 0.770 ;
        RECT 6.235 0.530 6.245 0.780 ;
        RECT 6.245 0.540 6.255 0.790 ;
        RECT 6.255 0.550 6.265 0.800 ;
        RECT 6.265 0.560 6.275 0.810 ;
        RECT 6.275 0.570 6.285 0.820 ;
        RECT 6.285 0.580 6.295 0.830 ;
        RECT 6.295 0.590 6.305 0.840 ;
        RECT 6.305 0.600 6.315 0.850 ;
        RECT 6.315 0.610 6.325 0.860 ;
        RECT 6.325 0.620 6.335 0.870 ;
        RECT 6.335 0.630 6.345 0.880 ;
        RECT 6.345 0.640 6.355 0.890 ;
        RECT 6.355 0.650 6.365 0.900 ;
        RECT 6.365 0.660 6.375 0.910 ;
        RECT 6.375 0.670 6.385 0.920 ;
        RECT 6.385 0.680 6.395 0.930 ;
        RECT 6.395 0.685 6.401 0.939 ;
        RECT 6.105 0.480 6.115 0.650 ;
        RECT 6.115 0.480 6.125 0.660 ;
        RECT 6.125 0.480 6.135 0.670 ;
        RECT 6.135 0.480 6.145 0.680 ;
        RECT 6.145 0.480 6.155 0.690 ;
        RECT 6.155 0.480 6.165 0.700 ;
        RECT 6.165 0.480 6.175 0.710 ;
        RECT 6.175 0.480 6.185 0.720 ;
        RECT 6.185 0.480 6.195 0.730 ;
        RECT 5.265 0.480 5.275 0.774 ;
        RECT 5.275 0.480 5.285 0.764 ;
        RECT 5.285 0.480 5.295 0.754 ;
        RECT 5.295 0.480 5.305 0.744 ;
        RECT 5.305 0.480 5.315 0.734 ;
        RECT 5.315 0.480 5.325 0.724 ;
        RECT 5.325 0.480 5.335 0.714 ;
        RECT 5.335 0.480 5.345 0.704 ;
        RECT 5.345 0.480 5.355 0.694 ;
        RECT 5.355 0.480 5.365 0.684 ;
        RECT 5.365 0.480 5.375 0.674 ;
        RECT 5.375 0.480 5.385 0.664 ;
        RECT 5.385 0.480 5.395 0.654 ;
        RECT 5.395 0.480 5.401 0.650 ;
        RECT 5.105 0.640 5.115 0.934 ;
        RECT 5.115 0.630 5.125 0.924 ;
        RECT 5.125 0.620 5.135 0.914 ;
        RECT 5.135 0.610 5.145 0.904 ;
        RECT 5.145 0.600 5.155 0.894 ;
        RECT 5.155 0.590 5.165 0.884 ;
        RECT 5.165 0.580 5.175 0.874 ;
        RECT 5.175 0.570 5.185 0.864 ;
        RECT 5.185 0.560 5.195 0.854 ;
        RECT 5.195 0.550 5.205 0.844 ;
        RECT 5.205 0.540 5.215 0.834 ;
        RECT 5.215 0.530 5.225 0.824 ;
        RECT 5.225 0.520 5.235 0.814 ;
        RECT 5.235 0.510 5.245 0.804 ;
        RECT 5.245 0.500 5.255 0.794 ;
        RECT 5.255 0.490 5.265 0.784 ;
        RECT 4.970 0.775 4.980 0.945 ;
        RECT 4.980 0.765 4.990 0.945 ;
        RECT 4.990 0.755 5.000 0.945 ;
        RECT 5.000 0.745 5.010 0.945 ;
        RECT 5.010 0.735 5.020 0.945 ;
        RECT 5.020 0.725 5.030 0.945 ;
        RECT 5.030 0.715 5.040 0.945 ;
        RECT 5.040 0.705 5.050 0.945 ;
        RECT 5.050 0.695 5.060 0.945 ;
        RECT 5.060 0.685 5.070 0.945 ;
        RECT 5.070 0.675 5.080 0.945 ;
        RECT 5.080 0.665 5.090 0.945 ;
        RECT 5.090 0.655 5.100 0.945 ;
        RECT 5.100 0.645 5.106 0.945 ;
        RECT 13.075 0.965 13.410 1.135 ;
        RECT 13.230 0.965 13.410 2.330 ;
        RECT 13.150 2.030 13.410 2.330 ;
        RECT 14.175 1.700 14.345 2.645 ;
        RECT 13.230 1.700 14.605 1.870 ;
        RECT 16.415 1.540 16.585 2.645 ;
        RECT 14.175 2.475 16.585 2.645 ;
  END 
END FFSEDCRHD2XHT

MACRO FFSDSRHDMXHT
  CLASS  CORE ;
  FOREIGN FFSDSRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.760 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.410 0.995 14.580 2.845 ;
        RECT 14.410 2.490 14.660 2.845 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.145 0.920 13.680 1.230 ;
        RECT 13.510 0.920 13.680 2.215 ;
        RECT 13.245 2.045 13.680 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 1.290 1.605 1.540 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.760 1.510 6.385 1.955 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.520 1.735 0.690 2.100 ;
        RECT 0.815 1.930 1.230 2.360 ;
        RECT 1.400 1.735 1.570 2.100 ;
        RECT 0.520 1.930 1.570 2.100 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.995 ;
        RECT 2.495 -0.300 2.795 0.785 ;
        RECT 3.230 -0.300 3.530 0.745 ;
        RECT 5.970 -0.300 6.270 1.130 ;
        RECT 8.765 -0.300 8.935 1.360 ;
        RECT 10.645 -0.300 10.945 0.795 ;
        RECT 12.665 -0.300 12.965 1.280 ;
        RECT 13.860 -0.300 14.030 1.145 ;
        RECT 0.000 -0.300 14.760 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.965 1.550 3.305 2.015 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.290 1.610 2.775 2.015 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 12.175 1.540 12.675 1.950 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.905 0.895 3.990 ;
        RECT 2.540 2.895 3.520 3.990 ;
        RECT 6.145 2.995 7.125 3.990 ;
        RECT 8.675 2.995 8.975 3.990 ;
        RECT 10.700 2.315 11.000 3.990 ;
        RECT 12.605 2.975 12.905 3.990 ;
        RECT 13.795 2.790 14.095 3.990 ;
        RECT 0.000 3.390 14.760 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.170 0.340 2.470 ;
        RECT 0.105 0.825 0.275 2.470 ;
        RECT 0.170 2.170 0.340 2.725 ;
        RECT 0.105 0.825 0.405 0.995 ;
        RECT 0.170 2.555 1.305 2.725 ;
        RECT 1.135 2.555 1.305 3.130 ;
        RECT 1.135 2.960 1.995 3.130 ;
        RECT 2.770 1.125 3.310 1.295 ;
        RECT 2.825 2.195 3.580 2.365 ;
        RECT 3.580 1.290 3.590 2.364 ;
        RECT 3.590 1.300 3.600 2.364 ;
        RECT 3.600 1.310 3.610 2.364 ;
        RECT 3.610 1.320 3.620 2.364 ;
        RECT 3.620 1.330 3.630 2.364 ;
        RECT 3.630 1.340 3.640 2.364 ;
        RECT 3.640 1.350 3.650 2.364 ;
        RECT 3.650 1.360 3.660 2.364 ;
        RECT 3.660 1.370 3.670 2.364 ;
        RECT 3.670 1.380 3.680 2.364 ;
        RECT 3.680 1.390 3.690 2.364 ;
        RECT 3.690 1.400 3.700 2.364 ;
        RECT 3.700 1.410 3.710 2.364 ;
        RECT 3.710 1.420 3.720 2.364 ;
        RECT 3.720 1.430 3.730 2.364 ;
        RECT 3.730 1.440 3.740 2.364 ;
        RECT 3.740 1.450 3.750 2.364 ;
        RECT 3.425 1.135 3.435 1.409 ;
        RECT 3.435 1.145 3.445 1.419 ;
        RECT 3.445 1.155 3.455 1.429 ;
        RECT 3.455 1.165 3.465 1.439 ;
        RECT 3.465 1.175 3.475 1.449 ;
        RECT 3.475 1.185 3.485 1.459 ;
        RECT 3.485 1.195 3.495 1.469 ;
        RECT 3.495 1.205 3.505 1.479 ;
        RECT 3.505 1.215 3.515 1.489 ;
        RECT 3.515 1.225 3.525 1.499 ;
        RECT 3.525 1.235 3.535 1.509 ;
        RECT 3.535 1.245 3.545 1.519 ;
        RECT 3.545 1.255 3.555 1.529 ;
        RECT 3.555 1.265 3.565 1.539 ;
        RECT 3.565 1.275 3.575 1.549 ;
        RECT 3.575 1.280 3.581 1.560 ;
        RECT 3.310 1.125 3.320 1.295 ;
        RECT 3.320 1.125 3.330 1.305 ;
        RECT 3.330 1.125 3.340 1.315 ;
        RECT 3.340 1.125 3.350 1.325 ;
        RECT 3.350 1.125 3.360 1.335 ;
        RECT 3.360 1.125 3.370 1.345 ;
        RECT 3.370 1.125 3.380 1.355 ;
        RECT 3.380 1.125 3.390 1.365 ;
        RECT 3.390 1.125 3.400 1.375 ;
        RECT 3.400 1.125 3.410 1.385 ;
        RECT 3.410 1.125 3.420 1.395 ;
        RECT 3.420 1.125 3.426 1.405 ;
        RECT 1.545 0.790 1.985 0.960 ;
        RECT 1.815 0.790 1.985 2.715 ;
        RECT 1.580 2.370 1.985 2.715 ;
        RECT 1.580 2.545 3.655 2.715 ;
        RECT 4.445 0.895 4.555 2.830 ;
        RECT 3.845 2.660 4.555 2.830 ;
        RECT 4.555 1.575 4.565 2.829 ;
        RECT 4.565 1.585 4.575 2.829 ;
        RECT 4.575 1.595 4.585 2.829 ;
        RECT 4.585 1.605 4.595 2.829 ;
        RECT 4.595 1.615 4.605 2.829 ;
        RECT 4.605 1.625 4.615 2.829 ;
        RECT 4.385 0.895 4.395 1.659 ;
        RECT 4.395 0.895 4.405 1.669 ;
        RECT 4.405 0.895 4.415 1.679 ;
        RECT 4.415 0.895 4.425 1.689 ;
        RECT 4.425 0.895 4.435 1.699 ;
        RECT 4.435 0.895 4.445 1.709 ;
        RECT 3.770 2.595 3.780 2.829 ;
        RECT 3.780 2.605 3.790 2.829 ;
        RECT 3.790 2.615 3.800 2.829 ;
        RECT 3.800 2.625 3.810 2.829 ;
        RECT 3.810 2.635 3.820 2.829 ;
        RECT 3.820 2.645 3.830 2.829 ;
        RECT 3.830 2.655 3.840 2.829 ;
        RECT 3.840 2.660 3.846 2.830 ;
        RECT 3.730 2.555 3.740 2.789 ;
        RECT 3.740 2.565 3.750 2.799 ;
        RECT 3.750 2.575 3.760 2.809 ;
        RECT 3.760 2.585 3.770 2.819 ;
        RECT 3.655 2.545 3.665 2.715 ;
        RECT 3.665 2.545 3.675 2.725 ;
        RECT 3.675 2.545 3.685 2.735 ;
        RECT 3.685 2.545 3.695 2.745 ;
        RECT 3.695 2.545 3.705 2.755 ;
        RECT 3.705 2.545 3.715 2.765 ;
        RECT 3.715 2.545 3.725 2.775 ;
        RECT 3.725 2.545 3.731 2.785 ;
        RECT 6.585 0.960 6.755 2.115 ;
        RECT 6.490 0.960 6.790 1.130 ;
        RECT 6.585 1.500 7.360 1.670 ;
        RECT 5.085 0.895 5.315 1.195 ;
        RECT 5.095 0.895 5.315 1.205 ;
        RECT 5.105 0.895 5.315 1.215 ;
        RECT 5.115 0.895 5.315 1.225 ;
        RECT 5.125 0.895 5.315 1.235 ;
        RECT 5.135 0.895 5.315 1.245 ;
        RECT 5.145 0.895 5.315 2.465 ;
        RECT 7.540 1.680 7.710 2.465 ;
        RECT 5.145 2.295 7.710 2.465 ;
        RECT 7.775 1.550 7.945 1.850 ;
        RECT 7.540 1.680 7.945 1.850 ;
        RECT 7.000 0.960 7.300 1.230 ;
        RECT 7.000 1.060 8.235 1.230 ;
        RECT 8.065 1.060 8.235 1.360 ;
        RECT 6.630 0.480 6.930 0.730 ;
        RECT 7.890 2.045 8.015 2.215 ;
        RECT 8.125 1.580 8.190 2.215 ;
        RECT 6.630 0.560 8.585 0.730 ;
        RECT 8.415 0.560 8.585 1.750 ;
        RECT 8.295 1.580 9.180 1.750 ;
        RECT 8.190 1.580 8.200 2.104 ;
        RECT 8.200 1.580 8.210 2.094 ;
        RECT 8.210 1.580 8.220 2.084 ;
        RECT 8.220 1.580 8.230 2.074 ;
        RECT 8.230 1.580 8.240 2.064 ;
        RECT 8.240 1.580 8.250 2.054 ;
        RECT 8.250 1.580 8.260 2.044 ;
        RECT 8.260 1.580 8.270 2.034 ;
        RECT 8.270 1.580 8.280 2.024 ;
        RECT 8.280 1.580 8.290 2.014 ;
        RECT 8.290 1.580 8.296 2.010 ;
        RECT 8.015 2.045 8.025 2.215 ;
        RECT 8.025 2.035 8.035 2.215 ;
        RECT 8.035 2.025 8.045 2.215 ;
        RECT 8.045 2.015 8.055 2.215 ;
        RECT 8.055 2.005 8.065 2.215 ;
        RECT 8.065 1.995 8.075 2.215 ;
        RECT 8.075 1.985 8.085 2.215 ;
        RECT 8.085 1.975 8.095 2.215 ;
        RECT 8.095 1.965 8.105 2.215 ;
        RECT 8.105 1.955 8.115 2.215 ;
        RECT 8.115 1.945 8.125 2.215 ;
        RECT 3.875 0.895 4.205 1.195 ;
        RECT 3.970 0.895 4.205 2.430 ;
        RECT 4.000 0.545 4.205 2.430 ;
        RECT 3.930 2.130 4.205 2.430 ;
        RECT 4.000 0.545 4.735 0.715 ;
        RECT 4.795 0.545 4.905 2.835 ;
        RECT 4.795 0.545 5.530 0.715 ;
        RECT 4.965 2.645 8.020 2.815 ;
        RECT 8.445 2.295 9.205 2.465 ;
        RECT 9.380 2.395 10.105 2.565 ;
        RECT 9.935 2.395 10.105 2.695 ;
        RECT 9.305 2.330 9.315 2.564 ;
        RECT 9.315 2.340 9.325 2.564 ;
        RECT 9.325 2.350 9.335 2.564 ;
        RECT 9.335 2.360 9.345 2.564 ;
        RECT 9.345 2.370 9.355 2.564 ;
        RECT 9.355 2.380 9.365 2.564 ;
        RECT 9.365 2.390 9.375 2.564 ;
        RECT 9.375 2.395 9.381 2.565 ;
        RECT 9.280 2.305 9.290 2.539 ;
        RECT 9.290 2.315 9.300 2.549 ;
        RECT 9.300 2.320 9.306 2.560 ;
        RECT 9.205 2.295 9.215 2.465 ;
        RECT 9.215 2.295 9.225 2.475 ;
        RECT 9.225 2.295 9.235 2.485 ;
        RECT 9.235 2.295 9.245 2.495 ;
        RECT 9.245 2.295 9.255 2.505 ;
        RECT 9.255 2.295 9.265 2.515 ;
        RECT 9.265 2.295 9.275 2.525 ;
        RECT 9.275 2.295 9.281 2.535 ;
        RECT 8.370 2.295 8.380 2.529 ;
        RECT 8.380 2.295 8.390 2.519 ;
        RECT 8.390 2.295 8.400 2.509 ;
        RECT 8.400 2.295 8.410 2.499 ;
        RECT 8.410 2.295 8.420 2.489 ;
        RECT 8.420 2.295 8.430 2.479 ;
        RECT 8.430 2.295 8.440 2.469 ;
        RECT 8.440 2.295 8.446 2.465 ;
        RECT 8.095 2.570 8.105 2.804 ;
        RECT 8.105 2.560 8.115 2.794 ;
        RECT 8.115 2.550 8.125 2.784 ;
        RECT 8.125 2.540 8.135 2.774 ;
        RECT 8.135 2.530 8.145 2.764 ;
        RECT 8.145 2.520 8.155 2.754 ;
        RECT 8.155 2.510 8.165 2.744 ;
        RECT 8.165 2.500 8.175 2.734 ;
        RECT 8.175 2.490 8.185 2.724 ;
        RECT 8.185 2.480 8.195 2.714 ;
        RECT 8.195 2.470 8.205 2.704 ;
        RECT 8.205 2.460 8.215 2.694 ;
        RECT 8.215 2.450 8.225 2.684 ;
        RECT 8.225 2.440 8.235 2.674 ;
        RECT 8.235 2.430 8.245 2.664 ;
        RECT 8.245 2.420 8.255 2.654 ;
        RECT 8.255 2.410 8.265 2.644 ;
        RECT 8.265 2.400 8.275 2.634 ;
        RECT 8.275 2.390 8.285 2.624 ;
        RECT 8.285 2.380 8.295 2.614 ;
        RECT 8.295 2.370 8.305 2.604 ;
        RECT 8.305 2.360 8.315 2.594 ;
        RECT 8.315 2.350 8.325 2.584 ;
        RECT 8.325 2.340 8.335 2.574 ;
        RECT 8.335 2.330 8.345 2.564 ;
        RECT 8.345 2.320 8.355 2.554 ;
        RECT 8.355 2.310 8.365 2.544 ;
        RECT 8.365 2.300 8.371 2.540 ;
        RECT 8.020 2.645 8.030 2.815 ;
        RECT 8.030 2.635 8.040 2.815 ;
        RECT 8.040 2.625 8.050 2.815 ;
        RECT 8.050 2.615 8.060 2.815 ;
        RECT 8.060 2.605 8.070 2.815 ;
        RECT 8.070 2.595 8.080 2.815 ;
        RECT 8.080 2.585 8.090 2.815 ;
        RECT 8.090 2.575 8.096 2.815 ;
        RECT 4.905 1.340 4.915 2.834 ;
        RECT 4.915 1.350 4.925 2.834 ;
        RECT 4.925 1.360 4.935 2.834 ;
        RECT 4.935 1.370 4.945 2.834 ;
        RECT 4.945 1.380 4.955 2.834 ;
        RECT 4.955 1.390 4.965 2.834 ;
        RECT 4.735 0.545 4.745 1.425 ;
        RECT 4.745 0.545 4.755 1.435 ;
        RECT 4.755 0.545 4.765 1.445 ;
        RECT 4.765 0.545 4.775 1.455 ;
        RECT 4.775 0.545 4.785 1.465 ;
        RECT 4.785 0.545 4.795 1.475 ;
        RECT 7.340 2.995 7.640 3.210 ;
        RECT 7.340 2.995 8.325 3.165 ;
        RECT 8.595 2.645 9.050 2.815 ;
        RECT 9.495 2.745 9.665 3.045 ;
        RECT 9.225 2.745 9.665 2.915 ;
        RECT 9.955 1.270 10.255 1.440 ;
        RECT 10.085 1.270 10.255 1.825 ;
        RECT 10.085 1.655 10.455 1.825 ;
        RECT 10.285 1.655 10.455 3.045 ;
        RECT 9.495 2.875 10.455 3.045 ;
        RECT 9.150 2.680 9.160 2.914 ;
        RECT 9.160 2.690 9.170 2.914 ;
        RECT 9.170 2.700 9.180 2.914 ;
        RECT 9.180 2.710 9.190 2.914 ;
        RECT 9.190 2.720 9.200 2.914 ;
        RECT 9.200 2.730 9.210 2.914 ;
        RECT 9.210 2.740 9.220 2.914 ;
        RECT 9.220 2.745 9.226 2.915 ;
        RECT 9.125 2.655 9.135 2.889 ;
        RECT 9.135 2.665 9.145 2.899 ;
        RECT 9.145 2.670 9.151 2.910 ;
        RECT 9.050 2.645 9.060 2.815 ;
        RECT 9.060 2.645 9.070 2.825 ;
        RECT 9.070 2.645 9.080 2.835 ;
        RECT 9.080 2.645 9.090 2.845 ;
        RECT 9.090 2.645 9.100 2.855 ;
        RECT 9.100 2.645 9.110 2.865 ;
        RECT 9.110 2.645 9.120 2.875 ;
        RECT 9.120 2.645 9.126 2.885 ;
        RECT 8.520 2.645 8.530 2.879 ;
        RECT 8.530 2.645 8.540 2.869 ;
        RECT 8.540 2.645 8.550 2.859 ;
        RECT 8.550 2.645 8.560 2.849 ;
        RECT 8.560 2.645 8.570 2.839 ;
        RECT 8.570 2.645 8.580 2.829 ;
        RECT 8.580 2.645 8.590 2.819 ;
        RECT 8.590 2.645 8.596 2.815 ;
        RECT 8.495 2.670 8.505 2.904 ;
        RECT 8.505 2.660 8.515 2.894 ;
        RECT 8.515 2.650 8.521 2.890 ;
        RECT 8.325 2.840 8.335 3.164 ;
        RECT 8.335 2.830 8.345 3.164 ;
        RECT 8.345 2.820 8.355 3.164 ;
        RECT 8.355 2.810 8.365 3.164 ;
        RECT 8.365 2.800 8.375 3.164 ;
        RECT 8.375 2.790 8.385 3.164 ;
        RECT 8.385 2.780 8.395 3.164 ;
        RECT 8.395 2.770 8.405 3.164 ;
        RECT 8.405 2.760 8.415 3.164 ;
        RECT 8.415 2.750 8.425 3.164 ;
        RECT 8.425 2.740 8.435 3.164 ;
        RECT 8.435 2.730 8.445 3.164 ;
        RECT 8.445 2.720 8.455 3.164 ;
        RECT 8.455 2.710 8.465 3.164 ;
        RECT 8.465 2.700 8.475 3.164 ;
        RECT 8.475 2.690 8.485 3.164 ;
        RECT 8.485 2.680 8.495 3.164 ;
        RECT 11.205 0.760 11.375 1.280 ;
        RECT 11.075 1.110 11.375 1.280 ;
        RECT 11.205 0.760 12.285 0.930 ;
        RECT 12.115 0.760 12.285 1.280 ;
        RECT 12.115 1.110 12.415 1.280 ;
        RECT 10.985 1.460 11.155 1.760 ;
        RECT 11.595 1.110 11.895 1.630 ;
        RECT 10.985 1.460 11.895 1.630 ;
        RECT 11.725 1.110 11.895 2.300 ;
        RECT 12.110 2.130 12.295 2.345 ;
        RECT 11.725 2.130 12.295 2.300 ;
        RECT 12.895 1.475 13.065 2.345 ;
        RECT 12.110 2.175 13.065 2.345 ;
        RECT 12.895 1.475 13.330 1.775 ;
        RECT 9.545 0.900 9.715 2.215 ;
        RECT 9.545 2.045 9.845 2.215 ;
        RECT 9.545 0.900 10.330 1.070 ;
        RECT 10.565 1.060 10.805 1.230 ;
        RECT 10.635 1.060 10.805 2.110 ;
        RECT 10.635 1.940 11.390 2.110 ;
        RECT 11.220 1.940 11.390 2.795 ;
        RECT 11.815 2.625 12.115 2.855 ;
        RECT 13.335 2.440 13.505 2.795 ;
        RECT 11.220 2.625 13.505 2.795 ;
        RECT 13.990 1.520 14.160 2.610 ;
        RECT 13.335 2.440 14.160 2.610 ;
        RECT 13.990 1.520 14.230 1.820 ;
        RECT 10.490 0.995 10.500 1.229 ;
        RECT 10.500 1.005 10.510 1.229 ;
        RECT 10.510 1.015 10.520 1.229 ;
        RECT 10.520 1.025 10.530 1.229 ;
        RECT 10.530 1.035 10.540 1.229 ;
        RECT 10.540 1.045 10.550 1.229 ;
        RECT 10.550 1.055 10.560 1.229 ;
        RECT 10.560 1.060 10.566 1.230 ;
        RECT 10.405 0.910 10.415 1.144 ;
        RECT 10.415 0.920 10.425 1.154 ;
        RECT 10.425 0.930 10.435 1.164 ;
        RECT 10.435 0.940 10.445 1.174 ;
        RECT 10.445 0.950 10.455 1.184 ;
        RECT 10.455 0.960 10.465 1.194 ;
        RECT 10.465 0.970 10.475 1.204 ;
        RECT 10.475 0.980 10.485 1.214 ;
        RECT 10.485 0.985 10.491 1.225 ;
        RECT 10.330 0.900 10.340 1.070 ;
        RECT 10.340 0.900 10.350 1.080 ;
        RECT 10.350 0.900 10.360 1.090 ;
        RECT 10.360 0.900 10.370 1.100 ;
        RECT 10.370 0.900 10.380 1.110 ;
        RECT 10.380 0.900 10.390 1.120 ;
        RECT 10.390 0.900 10.400 1.130 ;
        RECT 10.400 0.900 10.406 1.140 ;
  END 
END FFSDSRHDMXHT

MACRO FFSDSHQHD2XHT
  CLASS  CORE ;
  FOREIGN FFSDSHQHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.760 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.870 0.595 14.135 2.960 ;
        RECT 13.870 1.265 14.250 1.980 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.150 1.165 1.775 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.545 0.380 2.020 ;
        RECT 0.285 2.580 0.470 2.840 ;
        RECT 0.170 2.670 0.470 2.840 ;
        RECT 0.285 2.580 1.340 2.750 ;
        RECT 0.170 2.670 1.340 2.750 ;
        RECT 1.170 2.580 1.340 3.190 ;
        RECT 1.170 3.020 2.245 3.190 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.955 ;
        RECT 2.540 -0.300 2.850 0.435 ;
        RECT 3.450 -0.300 3.750 0.435 ;
        RECT 4.510 -0.300 4.810 0.435 ;
        RECT 7.480 -0.300 7.780 0.595 ;
        RECT 10.135 -0.300 10.440 0.665 ;
        RECT 12.120 -0.300 12.295 0.850 ;
        RECT 13.320 -0.300 13.490 0.780 ;
        RECT 14.420 -0.300 14.590 1.120 ;
        RECT 0.000 -0.300 14.760 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 4.510 1.570 5.025 2.020 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.145 1.435 2.500 2.055 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 8.850 2.340 9.020 2.880 ;
        RECT 8.850 2.710 12.915 2.880 ;
        RECT 12.400 2.490 12.615 2.880 ;
        RECT 12.615 2.690 12.915 2.925 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.945 0.955 3.990 ;
        RECT 2.560 2.830 2.740 3.990 ;
        RECT 3.580 2.745 3.880 3.990 ;
        RECT 4.395 2.745 4.695 3.990 ;
        RECT 7.380 3.065 7.680 3.990 ;
        RECT 8.480 3.095 8.780 3.990 ;
        RECT 10.135 3.095 10.435 3.990 ;
        RECT 12.055 3.095 12.355 3.990 ;
        RECT 13.320 2.910 13.490 3.990 ;
        RECT 14.420 2.230 14.590 3.990 ;
        RECT 0.000 3.390 14.760 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.020 0.340 1.320 ;
        RECT 0.170 1.150 0.730 1.320 ;
        RECT 0.560 1.150 0.730 2.370 ;
        RECT 0.105 2.200 0.730 2.370 ;
        RECT 1.780 1.460 1.950 2.125 ;
        RECT 0.560 1.955 1.950 2.125 ;
        RECT 3.405 1.605 3.575 1.905 ;
        RECT 3.405 1.605 4.300 1.780 ;
        RECT 4.000 1.125 4.300 2.215 ;
        RECT 5.070 1.125 5.700 1.295 ;
        RECT 5.530 1.125 5.700 2.215 ;
        RECT 5.315 2.045 5.700 2.215 ;
        RECT 1.575 2.330 1.875 2.840 ;
        RECT 1.575 0.825 2.850 1.005 ;
        RECT 2.680 0.615 2.850 2.500 ;
        RECT 1.575 2.330 2.850 2.500 ;
        RECT 2.680 0.615 6.115 0.785 ;
        RECT 5.945 0.615 6.115 2.415 ;
        RECT 6.645 1.060 6.815 2.365 ;
        RECT 7.785 1.695 7.955 2.080 ;
        RECT 6.645 1.910 7.955 2.080 ;
        RECT 7.305 1.125 7.475 1.730 ;
        RECT 8.135 1.125 8.305 2.520 ;
        RECT 7.930 2.350 8.305 2.520 ;
        RECT 7.305 1.125 8.750 1.295 ;
        RECT 8.135 1.570 10.565 1.740 ;
        RECT 3.030 1.060 3.200 2.735 ;
        RECT 3.030 1.060 3.255 1.360 ;
        RECT 3.030 2.095 3.320 2.735 ;
        RECT 3.030 2.395 5.435 2.565 ;
        RECT 5.135 2.395 5.435 2.825 ;
        RECT 6.295 0.550 6.465 2.825 ;
        RECT 5.135 2.655 6.465 2.825 ;
        RECT 6.295 0.550 7.205 0.730 ;
        RECT 6.985 0.550 7.205 0.945 ;
        RECT 6.985 0.775 8.830 0.945 ;
        RECT 9.100 0.970 9.500 1.140 ;
        RECT 9.330 0.970 9.500 1.365 ;
        RECT 9.330 1.195 11.060 1.365 ;
        RECT 10.890 1.195 11.060 1.675 ;
        RECT 9.025 0.905 9.035 1.139 ;
        RECT 9.035 0.915 9.045 1.139 ;
        RECT 9.045 0.925 9.055 1.139 ;
        RECT 9.055 0.935 9.065 1.139 ;
        RECT 9.065 0.945 9.075 1.139 ;
        RECT 9.075 0.955 9.085 1.139 ;
        RECT 9.085 0.965 9.095 1.139 ;
        RECT 9.095 0.970 9.101 1.140 ;
        RECT 8.905 0.785 8.915 1.019 ;
        RECT 8.915 0.795 8.925 1.029 ;
        RECT 8.925 0.805 8.935 1.039 ;
        RECT 8.935 0.815 8.945 1.049 ;
        RECT 8.945 0.825 8.955 1.059 ;
        RECT 8.955 0.835 8.965 1.069 ;
        RECT 8.965 0.845 8.975 1.079 ;
        RECT 8.975 0.855 8.985 1.089 ;
        RECT 8.985 0.865 8.995 1.099 ;
        RECT 8.995 0.875 9.005 1.109 ;
        RECT 9.005 0.885 9.015 1.119 ;
        RECT 9.015 0.895 9.025 1.129 ;
        RECT 8.830 0.775 8.840 0.945 ;
        RECT 8.840 0.775 8.850 0.955 ;
        RECT 8.850 0.775 8.860 0.965 ;
        RECT 8.860 0.775 8.870 0.975 ;
        RECT 8.870 0.775 8.880 0.985 ;
        RECT 8.880 0.775 8.890 0.995 ;
        RECT 8.890 0.775 8.900 1.005 ;
        RECT 8.900 0.775 8.906 1.015 ;
        RECT 8.485 1.990 8.655 2.875 ;
        RECT 6.755 2.705 8.655 2.875 ;
        RECT 11.260 0.985 11.430 2.160 ;
        RECT 8.485 1.990 11.430 2.160 ;
        RECT 11.260 0.985 11.590 1.285 ;
        RECT 9.150 0.590 9.910 0.760 ;
        RECT 9.740 0.590 9.910 1.015 ;
        RECT 10.850 0.615 11.020 1.015 ;
        RECT 9.740 0.845 11.020 1.015 ;
        RECT 10.850 0.615 11.940 0.785 ;
        RECT 11.610 1.540 11.780 2.530 ;
        RECT 9.215 2.360 11.780 2.530 ;
        RECT 11.770 0.615 11.940 1.710 ;
        RECT 11.610 1.540 13.310 1.710 ;
        RECT 13.140 1.475 13.310 1.775 ;
        RECT 11.960 1.890 12.130 2.245 ;
        RECT 11.960 2.075 12.965 2.245 ;
        RECT 12.795 2.075 12.965 2.505 ;
        RECT 12.415 1.125 13.680 1.295 ;
        RECT 13.490 1.125 13.680 2.505 ;
        RECT 12.795 2.335 13.680 2.505 ;
  END 
END FFSDSHQHD2XHT

MACRO FFSDQSRHDLXHT
  CLASS  CORE ;
  FOREIGN FFSDQSRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.530 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.190 1.045 13.430 2.430 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.835 1.290 1.605 1.540 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.760 1.740 6.385 2.055 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.520 1.735 0.690 2.100 ;
        RECT 0.815 1.930 1.230 2.360 ;
        RECT 1.370 1.735 1.540 2.100 ;
        RECT 0.520 1.930 1.540 2.100 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.090 ;
        RECT 2.525 -0.300 2.825 0.785 ;
        RECT 3.285 -0.300 3.585 0.745 ;
        RECT 5.930 -0.300 6.230 0.460 ;
        RECT 8.805 -0.300 9.380 0.795 ;
        RECT 10.645 -0.300 10.945 0.770 ;
        RECT 12.695 -0.300 12.995 0.715 ;
        RECT 0.000 -0.300 13.530 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.965 1.550 3.305 2.015 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.290 1.610 2.775 2.015 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 12.185 1.540 12.640 2.015 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 2.905 0.865 3.990 ;
        RECT 2.540 2.895 3.520 3.990 ;
        RECT 6.145 2.995 7.125 3.990 ;
        RECT 8.675 2.995 8.975 3.990 ;
        RECT 10.700 2.315 11.000 3.990 ;
        RECT 12.605 2.975 12.905 3.990 ;
        RECT 0.000 3.390 13.530 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.920 0.275 2.590 ;
        RECT 0.170 2.290 0.340 2.725 ;
        RECT 0.105 2.290 0.340 2.590 ;
        RECT 0.105 0.920 0.405 1.090 ;
        RECT 0.170 2.555 1.305 2.725 ;
        RECT 1.135 2.555 1.305 3.075 ;
        RECT 1.135 2.905 1.995 3.075 ;
        RECT 2.825 1.125 3.750 1.295 ;
        RECT 3.580 1.125 3.750 2.365 ;
        RECT 2.825 2.195 3.750 2.365 ;
        RECT 1.640 0.690 1.810 1.020 ;
        RECT 1.640 0.850 1.985 1.020 ;
        RECT 1.815 0.850 1.985 2.715 ;
        RECT 1.550 2.310 1.985 2.715 ;
        RECT 1.550 2.545 3.730 2.715 ;
        RECT 3.665 2.610 4.615 2.725 ;
        RECT 3.675 2.610 4.615 2.735 ;
        RECT 3.685 2.610 4.615 2.745 ;
        RECT 3.695 2.610 4.615 2.755 ;
        RECT 3.705 2.610 4.615 2.765 ;
        RECT 3.715 2.610 4.615 2.775 ;
        RECT 3.720 2.545 3.730 2.780 ;
        RECT 1.550 2.555 3.740 2.715 ;
        RECT 1.550 2.565 3.750 2.715 ;
        RECT 1.550 2.575 3.760 2.715 ;
        RECT 1.550 2.585 3.770 2.715 ;
        RECT 1.550 2.595 3.780 2.715 ;
        RECT 3.720 2.610 4.615 2.779 ;
        RECT 1.550 2.605 3.790 2.715 ;
        RECT 4.445 0.895 4.615 2.780 ;
        RECT 3.790 2.610 4.615 2.780 ;
        RECT 6.585 0.960 6.755 2.115 ;
        RECT 6.490 0.960 6.790 1.130 ;
        RECT 6.585 1.500 7.360 1.670 ;
        RECT 5.145 0.895 5.315 2.465 ;
        RECT 5.145 0.895 5.345 1.195 ;
        RECT 7.540 1.680 7.710 2.465 ;
        RECT 5.145 2.295 7.710 2.465 ;
        RECT 7.775 1.550 7.945 1.850 ;
        RECT 7.540 1.680 7.945 1.850 ;
        RECT 7.000 0.960 7.300 1.230 ;
        RECT 7.000 1.060 8.275 1.230 ;
        RECT 8.105 1.060 8.275 1.360 ;
        RECT 5.930 0.805 6.100 1.500 ;
        RECT 5.800 1.330 6.100 1.500 ;
        RECT 5.930 0.805 6.140 0.975 ;
        RECT 7.890 2.045 8.015 2.215 ;
        RECT 8.125 1.580 8.190 2.215 ;
        RECT 6.465 0.560 8.625 0.730 ;
        RECT 8.455 0.560 8.625 1.750 ;
        RECT 8.295 1.580 9.180 1.750 ;
        RECT 8.190 1.580 8.200 2.104 ;
        RECT 8.200 1.580 8.210 2.094 ;
        RECT 8.210 1.580 8.220 2.084 ;
        RECT 8.220 1.580 8.230 2.074 ;
        RECT 8.230 1.580 8.240 2.064 ;
        RECT 8.240 1.580 8.250 2.054 ;
        RECT 8.250 1.580 8.260 2.044 ;
        RECT 8.260 1.580 8.270 2.034 ;
        RECT 8.270 1.580 8.280 2.024 ;
        RECT 8.280 1.580 8.290 2.014 ;
        RECT 8.290 1.580 8.296 2.010 ;
        RECT 8.015 2.045 8.025 2.215 ;
        RECT 8.025 2.035 8.035 2.215 ;
        RECT 8.035 2.025 8.045 2.215 ;
        RECT 8.045 2.015 8.055 2.215 ;
        RECT 8.055 2.005 8.065 2.215 ;
        RECT 8.065 1.995 8.075 2.215 ;
        RECT 8.075 1.985 8.085 2.215 ;
        RECT 8.085 1.975 8.095 2.215 ;
        RECT 8.095 1.965 8.105 2.215 ;
        RECT 8.105 1.955 8.115 2.215 ;
        RECT 8.115 1.945 8.125 2.215 ;
        RECT 6.385 0.560 6.395 0.800 ;
        RECT 6.395 0.560 6.405 0.790 ;
        RECT 6.405 0.560 6.415 0.780 ;
        RECT 6.415 0.560 6.425 0.770 ;
        RECT 6.425 0.560 6.435 0.760 ;
        RECT 6.435 0.560 6.445 0.750 ;
        RECT 6.445 0.560 6.455 0.740 ;
        RECT 6.455 0.560 6.465 0.730 ;
        RECT 6.220 0.725 6.230 0.965 ;
        RECT 6.230 0.715 6.240 0.955 ;
        RECT 6.240 0.705 6.250 0.945 ;
        RECT 6.250 0.695 6.260 0.935 ;
        RECT 6.260 0.685 6.270 0.925 ;
        RECT 6.270 0.675 6.280 0.915 ;
        RECT 6.280 0.665 6.290 0.905 ;
        RECT 6.290 0.655 6.300 0.895 ;
        RECT 6.300 0.645 6.310 0.885 ;
        RECT 6.310 0.635 6.320 0.875 ;
        RECT 6.320 0.625 6.330 0.865 ;
        RECT 6.330 0.615 6.340 0.855 ;
        RECT 6.340 0.605 6.350 0.845 ;
        RECT 6.350 0.595 6.360 0.835 ;
        RECT 6.360 0.585 6.370 0.825 ;
        RECT 6.370 0.575 6.380 0.815 ;
        RECT 6.380 0.565 6.386 0.809 ;
        RECT 6.140 0.805 6.150 0.975 ;
        RECT 6.150 0.795 6.160 0.975 ;
        RECT 6.160 0.785 6.170 0.975 ;
        RECT 6.170 0.775 6.180 0.975 ;
        RECT 6.180 0.765 6.190 0.975 ;
        RECT 6.190 0.755 6.200 0.975 ;
        RECT 6.200 0.745 6.210 0.975 ;
        RECT 6.210 0.735 6.220 0.975 ;
        RECT 3.930 0.545 4.100 2.430 ;
        RECT 4.795 0.545 4.965 2.835 ;
        RECT 3.930 0.545 5.620 0.715 ;
        RECT 4.795 2.645 8.020 2.815 ;
        RECT 8.445 2.295 9.205 2.465 ;
        RECT 9.380 2.395 10.105 2.565 ;
        RECT 9.935 2.395 10.105 2.695 ;
        RECT 9.305 2.330 9.315 2.564 ;
        RECT 9.315 2.340 9.325 2.564 ;
        RECT 9.325 2.350 9.335 2.564 ;
        RECT 9.335 2.360 9.345 2.564 ;
        RECT 9.345 2.370 9.355 2.564 ;
        RECT 9.355 2.380 9.365 2.564 ;
        RECT 9.365 2.390 9.375 2.564 ;
        RECT 9.375 2.395 9.381 2.565 ;
        RECT 9.280 2.305 9.290 2.539 ;
        RECT 9.290 2.315 9.300 2.549 ;
        RECT 9.300 2.320 9.306 2.560 ;
        RECT 9.205 2.295 9.215 2.465 ;
        RECT 9.215 2.295 9.225 2.475 ;
        RECT 9.225 2.295 9.235 2.485 ;
        RECT 9.235 2.295 9.245 2.495 ;
        RECT 9.245 2.295 9.255 2.505 ;
        RECT 9.255 2.295 9.265 2.515 ;
        RECT 9.265 2.295 9.275 2.525 ;
        RECT 9.275 2.295 9.281 2.535 ;
        RECT 8.370 2.295 8.380 2.529 ;
        RECT 8.380 2.295 8.390 2.519 ;
        RECT 8.390 2.295 8.400 2.509 ;
        RECT 8.400 2.295 8.410 2.499 ;
        RECT 8.410 2.295 8.420 2.489 ;
        RECT 8.420 2.295 8.430 2.479 ;
        RECT 8.430 2.295 8.440 2.469 ;
        RECT 8.440 2.295 8.446 2.465 ;
        RECT 8.095 2.570 8.105 2.804 ;
        RECT 8.105 2.560 8.115 2.794 ;
        RECT 8.115 2.550 8.125 2.784 ;
        RECT 8.125 2.540 8.135 2.774 ;
        RECT 8.135 2.530 8.145 2.764 ;
        RECT 8.145 2.520 8.155 2.754 ;
        RECT 8.155 2.510 8.165 2.744 ;
        RECT 8.165 2.500 8.175 2.734 ;
        RECT 8.175 2.490 8.185 2.724 ;
        RECT 8.185 2.480 8.195 2.714 ;
        RECT 8.195 2.470 8.205 2.704 ;
        RECT 8.205 2.460 8.215 2.694 ;
        RECT 8.215 2.450 8.225 2.684 ;
        RECT 8.225 2.440 8.235 2.674 ;
        RECT 8.235 2.430 8.245 2.664 ;
        RECT 8.245 2.420 8.255 2.654 ;
        RECT 8.255 2.410 8.265 2.644 ;
        RECT 8.265 2.400 8.275 2.634 ;
        RECT 8.275 2.390 8.285 2.624 ;
        RECT 8.285 2.380 8.295 2.614 ;
        RECT 8.295 2.370 8.305 2.604 ;
        RECT 8.305 2.360 8.315 2.594 ;
        RECT 8.315 2.350 8.325 2.584 ;
        RECT 8.325 2.340 8.335 2.574 ;
        RECT 8.335 2.330 8.345 2.564 ;
        RECT 8.345 2.320 8.355 2.554 ;
        RECT 8.355 2.310 8.365 2.544 ;
        RECT 8.365 2.300 8.371 2.540 ;
        RECT 8.020 2.645 8.030 2.815 ;
        RECT 8.030 2.635 8.040 2.815 ;
        RECT 8.040 2.625 8.050 2.815 ;
        RECT 8.050 2.615 8.060 2.815 ;
        RECT 8.060 2.605 8.070 2.815 ;
        RECT 8.070 2.595 8.080 2.815 ;
        RECT 8.080 2.585 8.090 2.815 ;
        RECT 8.090 2.575 8.096 2.815 ;
        RECT 7.340 2.995 7.640 3.210 ;
        RECT 7.340 2.995 8.325 3.165 ;
        RECT 8.595 2.645 9.050 2.815 ;
        RECT 9.495 2.745 9.665 3.045 ;
        RECT 9.225 2.745 9.665 2.915 ;
        RECT 9.955 1.270 10.255 1.440 ;
        RECT 10.085 1.270 10.255 1.825 ;
        RECT 10.085 1.655 10.455 1.825 ;
        RECT 10.285 1.655 10.455 3.045 ;
        RECT 9.495 2.875 10.455 3.045 ;
        RECT 9.150 2.680 9.160 2.914 ;
        RECT 9.160 2.690 9.170 2.914 ;
        RECT 9.170 2.700 9.180 2.914 ;
        RECT 9.180 2.710 9.190 2.914 ;
        RECT 9.190 2.720 9.200 2.914 ;
        RECT 9.200 2.730 9.210 2.914 ;
        RECT 9.210 2.740 9.220 2.914 ;
        RECT 9.220 2.745 9.226 2.915 ;
        RECT 9.125 2.655 9.135 2.889 ;
        RECT 9.135 2.665 9.145 2.899 ;
        RECT 9.145 2.670 9.151 2.910 ;
        RECT 9.050 2.645 9.060 2.815 ;
        RECT 9.060 2.645 9.070 2.825 ;
        RECT 9.070 2.645 9.080 2.835 ;
        RECT 9.080 2.645 9.090 2.845 ;
        RECT 9.090 2.645 9.100 2.855 ;
        RECT 9.100 2.645 9.110 2.865 ;
        RECT 9.110 2.645 9.120 2.875 ;
        RECT 9.120 2.645 9.126 2.885 ;
        RECT 8.520 2.645 8.530 2.879 ;
        RECT 8.530 2.645 8.540 2.869 ;
        RECT 8.540 2.645 8.550 2.859 ;
        RECT 8.550 2.645 8.560 2.849 ;
        RECT 8.560 2.645 8.570 2.839 ;
        RECT 8.570 2.645 8.580 2.829 ;
        RECT 8.580 2.645 8.590 2.819 ;
        RECT 8.590 2.645 8.596 2.815 ;
        RECT 8.495 2.670 8.505 2.904 ;
        RECT 8.505 2.660 8.515 2.894 ;
        RECT 8.515 2.650 8.521 2.890 ;
        RECT 8.325 2.840 8.335 3.164 ;
        RECT 8.335 2.830 8.345 3.164 ;
        RECT 8.345 2.820 8.355 3.164 ;
        RECT 8.355 2.810 8.365 3.164 ;
        RECT 8.365 2.800 8.375 3.164 ;
        RECT 8.375 2.790 8.385 3.164 ;
        RECT 8.385 2.780 8.395 3.164 ;
        RECT 8.395 2.770 8.405 3.164 ;
        RECT 8.405 2.760 8.415 3.164 ;
        RECT 8.415 2.750 8.425 3.164 ;
        RECT 8.425 2.740 8.435 3.164 ;
        RECT 8.435 2.730 8.445 3.164 ;
        RECT 8.445 2.720 8.455 3.164 ;
        RECT 8.455 2.710 8.465 3.164 ;
        RECT 8.465 2.700 8.475 3.164 ;
        RECT 8.475 2.690 8.485 3.164 ;
        RECT 8.485 2.680 8.495 3.164 ;
        RECT 10.985 1.460 11.155 1.760 ;
        RECT 11.615 1.110 11.915 1.630 ;
        RECT 10.985 1.460 11.915 1.630 ;
        RECT 11.725 1.110 11.915 2.365 ;
        RECT 11.725 2.195 12.325 2.365 ;
        RECT 11.205 0.520 11.375 1.280 ;
        RECT 11.035 1.110 11.375 1.280 ;
        RECT 11.205 0.520 12.385 0.690 ;
        RECT 9.650 0.900 9.715 2.215 ;
        RECT 9.650 2.045 9.875 2.215 ;
        RECT 9.780 0.900 10.330 1.070 ;
        RECT 10.565 1.060 10.805 1.230 ;
        RECT 10.635 1.060 10.805 2.110 ;
        RECT 10.635 1.940 11.390 2.110 ;
        RECT 11.220 1.940 11.390 2.795 ;
        RECT 12.840 1.610 13.010 2.795 ;
        RECT 11.220 2.625 13.010 2.795 ;
        RECT 10.490 0.995 10.500 1.229 ;
        RECT 10.500 1.005 10.510 1.229 ;
        RECT 10.510 1.015 10.520 1.229 ;
        RECT 10.520 1.025 10.530 1.229 ;
        RECT 10.530 1.035 10.540 1.229 ;
        RECT 10.540 1.045 10.550 1.229 ;
        RECT 10.550 1.055 10.560 1.229 ;
        RECT 10.560 1.060 10.566 1.230 ;
        RECT 10.405 0.910 10.415 1.144 ;
        RECT 10.415 0.920 10.425 1.154 ;
        RECT 10.425 0.930 10.435 1.164 ;
        RECT 10.435 0.940 10.445 1.174 ;
        RECT 10.445 0.950 10.455 1.184 ;
        RECT 10.455 0.960 10.465 1.194 ;
        RECT 10.465 0.970 10.475 1.204 ;
        RECT 10.475 0.980 10.485 1.214 ;
        RECT 10.485 0.985 10.491 1.225 ;
        RECT 10.330 0.900 10.340 1.070 ;
        RECT 10.340 0.900 10.350 1.080 ;
        RECT 10.350 0.900 10.360 1.090 ;
        RECT 10.360 0.900 10.370 1.100 ;
        RECT 10.370 0.900 10.380 1.110 ;
        RECT 10.380 0.900 10.390 1.120 ;
        RECT 10.390 0.900 10.400 1.130 ;
        RECT 10.400 0.900 10.406 1.140 ;
        RECT 9.715 0.900 9.725 1.124 ;
        RECT 9.725 0.900 9.735 1.114 ;
        RECT 9.735 0.900 9.745 1.104 ;
        RECT 9.745 0.900 9.755 1.094 ;
        RECT 9.755 0.900 9.765 1.084 ;
        RECT 9.765 0.900 9.775 1.074 ;
        RECT 9.775 0.900 9.781 1.070 ;
        RECT 9.545 1.005 9.555 2.215 ;
        RECT 9.555 0.995 9.565 2.215 ;
        RECT 9.565 0.985 9.575 2.215 ;
        RECT 9.575 0.975 9.585 2.215 ;
        RECT 9.585 0.965 9.595 2.215 ;
        RECT 9.595 0.955 9.605 2.215 ;
        RECT 9.605 0.945 9.615 2.215 ;
        RECT 9.615 0.935 9.625 2.215 ;
        RECT 9.625 0.925 9.635 2.215 ;
        RECT 9.635 0.915 9.645 2.215 ;
        RECT 9.645 0.905 9.651 2.215 ;
  END 
END FFSDQSRHDLXHT

MACRO FFSDQSHD1XHT
  CLASS  CORE ;
  FOREIGN FFSDQSHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.480 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.140 0.720 11.380 1.360 ;
        RECT 11.170 0.720 11.380 2.960 ;
        RECT 11.140 1.980 11.380 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.385 -0.300 2.685 0.595 ;
        RECT 3.390 -0.300 3.690 0.595 ;
        RECT 6.950 -0.300 7.460 0.780 ;
        RECT 9.260 -0.300 9.430 0.640 ;
        RECT 10.555 -0.300 10.855 1.055 ;
        RECT 0.000 -0.300 11.480 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.850 1.525 3.340 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.245 2.410 1.800 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.640 0.605 7.810 1.910 ;
        RECT 6.995 1.610 7.810 1.910 ;
        RECT 7.640 0.605 9.015 0.775 ;
        RECT 8.845 0.605 9.015 1.145 ;
        RECT 9.705 0.540 9.875 1.145 ;
        RECT 8.845 0.920 9.875 1.145 ;
        RECT 9.705 0.540 10.165 0.710 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.355 2.345 2.655 3.990 ;
        RECT 3.235 2.675 3.405 3.990 ;
        RECT 5.965 3.160 6.265 3.990 ;
        RECT 7.140 3.160 7.440 3.990 ;
        RECT 9.215 2.770 9.515 3.990 ;
        RECT 9.855 2.945 10.155 3.990 ;
        RECT 10.555 2.975 10.855 3.990 ;
        RECT 0.000 3.390 11.480 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.555 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.150 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.985 0.775 2.155 1.035 ;
        RECT 1.530 0.865 2.155 1.035 ;
        RECT 1.985 0.775 4.620 0.945 ;
        RECT 4.450 0.775 4.620 2.280 ;
        RECT 5.150 0.900 5.320 2.280 ;
        RECT 5.150 1.605 6.465 1.775 ;
        RECT 6.645 1.060 6.815 2.215 ;
        RECT 6.515 2.045 6.815 2.215 ;
        RECT 6.645 1.060 7.460 1.360 ;
        RECT 2.840 1.125 3.695 1.295 ;
        RECT 2.865 2.190 3.755 2.360 ;
        RECT 3.525 1.125 3.695 2.360 ;
        RECT 3.585 1.525 3.755 2.980 ;
        RECT 3.525 1.525 3.770 1.825 ;
        RECT 3.585 2.810 8.315 2.980 ;
        RECT 3.875 1.125 4.195 1.295 ;
        RECT 3.940 1.980 4.195 2.280 ;
        RECT 4.025 1.125 4.195 2.630 ;
        RECT 4.800 0.535 4.970 2.630 ;
        RECT 4.800 0.535 5.595 0.705 ;
        RECT 7.990 1.645 8.160 2.630 ;
        RECT 8.020 1.245 8.190 1.815 ;
        RECT 7.990 1.645 8.190 1.815 ;
        RECT 4.025 2.460 8.830 2.630 ;
        RECT 8.660 2.460 8.830 2.795 ;
        RECT 9.015 1.325 10.280 1.495 ;
        RECT 10.110 0.890 10.280 2.215 ;
        RECT 9.795 2.045 10.280 2.215 ;
        RECT 8.415 0.955 8.585 2.215 ;
        RECT 8.325 0.955 8.625 1.125 ;
        RECT 8.340 2.045 8.640 2.215 ;
        RECT 9.120 1.675 9.290 2.590 ;
        RECT 8.415 1.675 9.865 1.845 ;
        RECT 10.790 1.610 10.960 2.590 ;
        RECT 9.120 2.420 10.960 2.590 ;
        RECT 10.790 1.610 10.970 1.910 ;
  END 
END FFSDQSHD1XHT

MACRO FFSDNSRHDLXHT
  CLASS  CORE ;
  FOREIGN FFSDNSRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.760 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.965 1.550 3.305 2.015 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.405 0.850 14.575 2.280 ;
        RECT 14.405 0.850 14.660 1.195 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.220 0.830 13.430 1.295 ;
        RECT 13.220 1.125 13.875 1.295 ;
        RECT 13.705 1.125 13.875 2.215 ;
        RECT 13.300 2.045 13.875 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.325 0.855 1.545 1.460 ;
        RECT 0.855 1.290 1.545 1.460 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.760 1.735 6.385 2.110 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.455 1.640 0.625 1.945 ;
        RECT 0.815 1.775 1.290 2.365 ;
        RECT 1.370 1.640 1.540 1.945 ;
        RECT 0.455 1.775 1.540 1.945 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.060 ;
        RECT 2.625 -0.300 2.925 0.785 ;
        RECT 3.285 -0.300 3.585 0.745 ;
        RECT 5.970 -0.300 6.270 1.130 ;
        RECT 8.860 -0.300 9.435 0.825 ;
        RECT 10.745 -0.300 11.045 0.795 ;
        RECT 12.740 -0.300 13.040 0.720 ;
        RECT 13.910 -0.300 14.210 0.715 ;
        RECT 0.000 -0.300 14.760 0.300 ;
    END
  END GND
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.290 1.610 2.775 2.015 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 12.330 1.540 12.760 1.950 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.545 2.975 0.845 3.990 ;
        RECT 2.470 2.995 3.450 3.990 ;
        RECT 6.170 2.995 7.150 3.990 ;
        RECT 8.675 2.995 8.975 3.990 ;
        RECT 10.800 2.535 11.100 3.990 ;
        RECT 12.860 2.830 13.115 3.990 ;
        RECT 13.790 2.830 14.090 3.990 ;
        RECT 0.000 3.390 14.760 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.130 0.340 2.430 ;
        RECT 0.105 0.890 0.275 2.430 ;
        RECT 0.170 2.130 0.340 2.795 ;
        RECT 0.105 0.890 0.405 1.060 ;
        RECT 0.170 2.625 1.305 2.795 ;
        RECT 1.135 2.625 1.305 3.065 ;
        RECT 1.135 2.895 1.995 3.065 ;
        RECT 2.795 1.125 3.750 1.295 ;
        RECT 3.580 1.125 3.750 2.365 ;
        RECT 2.825 2.195 3.750 2.365 ;
        RECT 1.740 0.825 1.985 1.125 ;
        RECT 1.815 0.825 1.985 2.715 ;
        RECT 1.580 2.150 1.985 2.715 ;
        RECT 4.445 1.045 4.615 2.715 ;
        RECT 1.580 2.545 4.615 2.715 ;
        RECT 3.930 0.695 4.100 2.290 ;
        RECT 3.930 0.695 5.545 0.865 ;
        RECT 5.375 0.695 5.545 2.245 ;
        RECT 6.555 0.895 6.755 1.195 ;
        RECT 6.585 0.895 6.755 2.115 ;
        RECT 6.585 1.445 6.795 2.115 ;
        RECT 6.585 1.445 7.345 1.745 ;
        RECT 5.025 1.045 5.195 2.595 ;
        RECT 5.025 2.425 5.715 2.595 ;
        RECT 7.525 1.680 7.695 2.465 ;
        RECT 5.920 2.295 7.695 2.465 ;
        RECT 7.775 1.550 7.945 1.850 ;
        RECT 7.525 1.680 7.945 1.850 ;
        RECT 5.845 2.295 5.855 2.529 ;
        RECT 5.855 2.295 5.865 2.519 ;
        RECT 5.865 2.295 5.875 2.509 ;
        RECT 5.875 2.295 5.885 2.499 ;
        RECT 5.885 2.295 5.895 2.489 ;
        RECT 5.895 2.295 5.905 2.479 ;
        RECT 5.905 2.295 5.915 2.469 ;
        RECT 5.915 2.295 5.921 2.465 ;
        RECT 5.790 2.350 5.800 2.584 ;
        RECT 5.800 2.340 5.810 2.574 ;
        RECT 5.810 2.330 5.820 2.564 ;
        RECT 5.820 2.320 5.830 2.554 ;
        RECT 5.830 2.310 5.840 2.544 ;
        RECT 5.840 2.300 5.846 2.540 ;
        RECT 5.715 2.425 5.725 2.595 ;
        RECT 5.725 2.415 5.735 2.595 ;
        RECT 5.735 2.405 5.745 2.595 ;
        RECT 5.745 2.395 5.755 2.595 ;
        RECT 5.755 2.385 5.765 2.595 ;
        RECT 5.765 2.375 5.775 2.595 ;
        RECT 5.775 2.365 5.785 2.595 ;
        RECT 5.785 2.355 5.791 2.595 ;
        RECT 7.000 0.960 7.300 1.215 ;
        RECT 7.000 1.045 8.275 1.215 ;
        RECT 8.105 1.045 8.275 1.345 ;
        RECT 6.990 0.525 7.160 0.730 ;
        RECT 6.630 0.525 7.160 0.695 ;
        RECT 7.890 2.045 8.015 2.215 ;
        RECT 8.125 1.535 8.190 2.215 ;
        RECT 6.990 0.560 8.625 0.730 ;
        RECT 8.455 0.560 8.625 1.705 ;
        RECT 8.295 1.535 9.210 1.705 ;
        RECT 8.190 1.535 8.200 2.105 ;
        RECT 8.200 1.535 8.210 2.095 ;
        RECT 8.210 1.535 8.220 2.085 ;
        RECT 8.220 1.535 8.230 2.075 ;
        RECT 8.230 1.535 8.240 2.065 ;
        RECT 8.240 1.535 8.250 2.055 ;
        RECT 8.250 1.535 8.260 2.045 ;
        RECT 8.260 1.535 8.270 2.035 ;
        RECT 8.270 1.535 8.280 2.025 ;
        RECT 8.280 1.535 8.290 2.015 ;
        RECT 8.290 1.535 8.296 2.009 ;
        RECT 8.015 2.045 8.025 2.215 ;
        RECT 8.025 2.035 8.035 2.215 ;
        RECT 8.035 2.025 8.045 2.215 ;
        RECT 8.045 2.015 8.055 2.215 ;
        RECT 8.055 2.005 8.065 2.215 ;
        RECT 8.065 1.995 8.075 2.215 ;
        RECT 8.075 1.985 8.085 2.215 ;
        RECT 8.085 1.975 8.095 2.215 ;
        RECT 8.095 1.965 8.105 2.215 ;
        RECT 8.105 1.955 8.115 2.215 ;
        RECT 8.115 1.945 8.125 2.215 ;
        RECT 3.655 2.895 5.745 3.065 ;
        RECT 7.900 2.395 8.070 2.815 ;
        RECT 6.095 2.645 8.070 2.815 ;
        RECT 7.900 2.395 8.270 2.565 ;
        RECT 8.445 2.295 9.260 2.465 ;
        RECT 10.100 1.810 10.270 2.565 ;
        RECT 9.435 2.395 10.270 2.565 ;
        RECT 9.360 2.330 9.370 2.564 ;
        RECT 9.370 2.340 9.380 2.564 ;
        RECT 9.380 2.350 9.390 2.564 ;
        RECT 9.390 2.360 9.400 2.564 ;
        RECT 9.400 2.370 9.410 2.564 ;
        RECT 9.410 2.380 9.420 2.564 ;
        RECT 9.420 2.390 9.430 2.564 ;
        RECT 9.430 2.395 9.436 2.565 ;
        RECT 9.335 2.305 9.345 2.539 ;
        RECT 9.345 2.315 9.355 2.549 ;
        RECT 9.355 2.320 9.361 2.560 ;
        RECT 9.260 2.295 9.270 2.465 ;
        RECT 9.270 2.295 9.280 2.475 ;
        RECT 9.280 2.295 9.290 2.485 ;
        RECT 9.290 2.295 9.300 2.495 ;
        RECT 9.300 2.295 9.310 2.505 ;
        RECT 9.310 2.295 9.320 2.515 ;
        RECT 9.320 2.295 9.330 2.525 ;
        RECT 9.330 2.295 9.336 2.535 ;
        RECT 8.370 2.295 8.380 2.529 ;
        RECT 8.380 2.295 8.390 2.519 ;
        RECT 8.390 2.295 8.400 2.509 ;
        RECT 8.400 2.295 8.410 2.499 ;
        RECT 8.410 2.295 8.420 2.489 ;
        RECT 8.420 2.295 8.430 2.479 ;
        RECT 8.430 2.295 8.440 2.469 ;
        RECT 8.440 2.295 8.446 2.465 ;
        RECT 8.345 2.320 8.355 2.554 ;
        RECT 8.355 2.310 8.365 2.544 ;
        RECT 8.365 2.300 8.371 2.540 ;
        RECT 8.270 2.395 8.280 2.565 ;
        RECT 8.280 2.385 8.290 2.565 ;
        RECT 8.290 2.375 8.300 2.565 ;
        RECT 8.300 2.365 8.310 2.565 ;
        RECT 8.310 2.355 8.320 2.565 ;
        RECT 8.320 2.345 8.330 2.565 ;
        RECT 8.330 2.335 8.340 2.565 ;
        RECT 8.340 2.325 8.346 2.565 ;
        RECT 5.995 2.645 6.005 2.905 ;
        RECT 6.005 2.645 6.015 2.895 ;
        RECT 6.015 2.645 6.025 2.885 ;
        RECT 6.025 2.645 6.035 2.875 ;
        RECT 6.035 2.645 6.045 2.865 ;
        RECT 6.045 2.645 6.055 2.855 ;
        RECT 6.055 2.645 6.065 2.845 ;
        RECT 6.065 2.645 6.075 2.835 ;
        RECT 6.075 2.645 6.085 2.825 ;
        RECT 6.085 2.645 6.095 2.815 ;
        RECT 5.845 2.795 5.855 3.055 ;
        RECT 5.855 2.785 5.865 3.045 ;
        RECT 5.865 2.775 5.875 3.035 ;
        RECT 5.875 2.765 5.885 3.025 ;
        RECT 5.885 2.755 5.895 3.015 ;
        RECT 5.895 2.745 5.905 3.005 ;
        RECT 5.905 2.735 5.915 2.995 ;
        RECT 5.915 2.725 5.925 2.985 ;
        RECT 5.925 2.715 5.935 2.975 ;
        RECT 5.935 2.705 5.945 2.965 ;
        RECT 5.945 2.695 5.955 2.955 ;
        RECT 5.955 2.685 5.965 2.945 ;
        RECT 5.965 2.675 5.975 2.935 ;
        RECT 5.975 2.665 5.985 2.925 ;
        RECT 5.985 2.655 5.995 2.915 ;
        RECT 5.745 2.895 5.755 3.065 ;
        RECT 5.755 2.885 5.765 3.065 ;
        RECT 5.765 2.875 5.775 3.065 ;
        RECT 5.775 2.865 5.785 3.065 ;
        RECT 5.785 2.855 5.795 3.065 ;
        RECT 5.795 2.845 5.805 3.065 ;
        RECT 5.805 2.835 5.815 3.065 ;
        RECT 5.815 2.825 5.825 3.065 ;
        RECT 5.825 2.815 5.835 3.065 ;
        RECT 5.835 2.805 5.845 3.065 ;
        RECT 7.485 3.040 8.275 3.210 ;
        RECT 8.600 2.645 9.105 2.815 ;
        RECT 10.055 1.325 10.350 1.495 ;
        RECT 9.280 2.745 10.450 2.915 ;
        RECT 10.450 1.360 10.460 2.914 ;
        RECT 10.460 1.370 10.470 2.914 ;
        RECT 10.470 1.380 10.480 2.914 ;
        RECT 10.480 1.390 10.490 2.914 ;
        RECT 10.490 1.400 10.500 2.914 ;
        RECT 10.500 1.410 10.510 2.914 ;
        RECT 10.510 1.420 10.520 2.914 ;
        RECT 10.520 1.430 10.530 2.914 ;
        RECT 10.530 1.440 10.540 2.914 ;
        RECT 10.540 1.450 10.550 2.914 ;
        RECT 10.550 1.460 10.560 2.914 ;
        RECT 10.560 1.470 10.570 2.914 ;
        RECT 10.570 1.480 10.580 2.914 ;
        RECT 10.580 1.490 10.590 2.914 ;
        RECT 10.590 1.500 10.600 2.914 ;
        RECT 10.600 1.510 10.610 2.914 ;
        RECT 10.610 1.520 10.620 2.914 ;
        RECT 10.425 1.335 10.435 1.569 ;
        RECT 10.435 1.345 10.445 1.579 ;
        RECT 10.445 1.350 10.451 1.590 ;
        RECT 10.350 1.325 10.360 1.495 ;
        RECT 10.360 1.325 10.370 1.505 ;
        RECT 10.370 1.325 10.380 1.515 ;
        RECT 10.380 1.325 10.390 1.525 ;
        RECT 10.390 1.325 10.400 1.535 ;
        RECT 10.400 1.325 10.410 1.545 ;
        RECT 10.410 1.325 10.420 1.555 ;
        RECT 10.420 1.325 10.426 1.565 ;
        RECT 9.205 2.680 9.215 2.914 ;
        RECT 9.215 2.690 9.225 2.914 ;
        RECT 9.225 2.700 9.235 2.914 ;
        RECT 9.235 2.710 9.245 2.914 ;
        RECT 9.245 2.720 9.255 2.914 ;
        RECT 9.255 2.730 9.265 2.914 ;
        RECT 9.265 2.740 9.275 2.914 ;
        RECT 9.275 2.745 9.281 2.915 ;
        RECT 9.180 2.655 9.190 2.889 ;
        RECT 9.190 2.665 9.200 2.899 ;
        RECT 9.200 2.670 9.206 2.910 ;
        RECT 9.105 2.645 9.115 2.815 ;
        RECT 9.115 2.645 9.125 2.825 ;
        RECT 9.125 2.645 9.135 2.835 ;
        RECT 9.135 2.645 9.145 2.845 ;
        RECT 9.145 2.645 9.155 2.855 ;
        RECT 9.155 2.645 9.165 2.865 ;
        RECT 9.165 2.645 9.175 2.875 ;
        RECT 9.175 2.645 9.181 2.885 ;
        RECT 8.525 2.645 8.535 2.879 ;
        RECT 8.535 2.645 8.545 2.869 ;
        RECT 8.545 2.645 8.555 2.859 ;
        RECT 8.555 2.645 8.565 2.849 ;
        RECT 8.565 2.645 8.575 2.839 ;
        RECT 8.575 2.645 8.585 2.829 ;
        RECT 8.585 2.645 8.595 2.819 ;
        RECT 8.595 2.645 8.601 2.815 ;
        RECT 8.445 2.725 8.455 2.959 ;
        RECT 8.455 2.715 8.465 2.949 ;
        RECT 8.465 2.705 8.475 2.939 ;
        RECT 8.475 2.695 8.485 2.929 ;
        RECT 8.485 2.685 8.495 2.919 ;
        RECT 8.495 2.675 8.505 2.909 ;
        RECT 8.505 2.665 8.515 2.899 ;
        RECT 8.515 2.655 8.525 2.889 ;
        RECT 8.275 2.895 8.285 3.209 ;
        RECT 8.285 2.885 8.295 3.209 ;
        RECT 8.295 2.875 8.305 3.209 ;
        RECT 8.305 2.865 8.315 3.209 ;
        RECT 8.315 2.855 8.325 3.209 ;
        RECT 8.325 2.845 8.335 3.209 ;
        RECT 8.335 2.835 8.345 3.209 ;
        RECT 8.345 2.825 8.355 3.209 ;
        RECT 8.355 2.815 8.365 3.209 ;
        RECT 8.365 2.805 8.375 3.209 ;
        RECT 8.375 2.795 8.385 3.209 ;
        RECT 8.385 2.785 8.395 3.209 ;
        RECT 8.395 2.775 8.405 3.209 ;
        RECT 8.405 2.765 8.415 3.209 ;
        RECT 8.415 2.755 8.425 3.209 ;
        RECT 8.425 2.745 8.435 3.209 ;
        RECT 8.435 2.735 8.445 3.209 ;
        RECT 11.355 0.760 11.525 1.280 ;
        RECT 11.150 1.110 11.525 1.280 ;
        RECT 11.355 0.760 12.435 0.930 ;
        RECT 12.265 0.760 12.435 1.280 ;
        RECT 12.265 1.110 12.610 1.280 ;
        RECT 11.150 1.460 11.320 2.005 ;
        RECT 11.730 1.110 12.030 1.630 ;
        RECT 11.150 1.460 12.030 1.630 ;
        RECT 11.860 1.110 12.030 2.415 ;
        RECT 11.860 2.245 12.330 2.415 ;
        RECT 12.940 1.540 13.110 2.300 ;
        RECT 12.530 2.130 13.110 2.300 ;
        RECT 12.940 1.540 13.525 1.840 ;
        RECT 12.445 2.130 12.455 2.374 ;
        RECT 12.455 2.130 12.465 2.364 ;
        RECT 12.465 2.130 12.475 2.354 ;
        RECT 12.475 2.130 12.485 2.344 ;
        RECT 12.485 2.130 12.495 2.334 ;
        RECT 12.495 2.130 12.505 2.324 ;
        RECT 12.505 2.130 12.515 2.314 ;
        RECT 12.515 2.130 12.525 2.304 ;
        RECT 12.525 2.130 12.531 2.300 ;
        RECT 12.415 2.160 12.425 2.404 ;
        RECT 12.425 2.150 12.435 2.394 ;
        RECT 12.435 2.140 12.445 2.384 ;
        RECT 12.330 2.245 12.340 2.415 ;
        RECT 12.340 2.235 12.350 2.415 ;
        RECT 12.350 2.225 12.360 2.415 ;
        RECT 12.360 2.215 12.370 2.415 ;
        RECT 12.370 2.205 12.380 2.415 ;
        RECT 12.380 2.195 12.390 2.415 ;
        RECT 12.390 2.185 12.400 2.415 ;
        RECT 12.400 2.175 12.410 2.415 ;
        RECT 12.410 2.165 12.416 2.415 ;
        RECT 9.620 0.900 9.790 2.215 ;
        RECT 9.620 2.045 9.920 2.215 ;
        RECT 9.620 0.900 10.430 1.070 ;
        RECT 10.645 1.040 10.970 1.210 ;
        RECT 10.800 1.040 10.970 2.355 ;
        RECT 10.800 2.185 11.530 2.355 ;
        RECT 11.360 2.185 11.530 2.810 ;
        RECT 11.935 2.640 12.235 2.970 ;
        RECT 11.360 2.640 12.445 2.810 ;
        RECT 14.055 1.540 14.225 2.650 ;
        RECT 12.720 2.480 14.225 2.650 ;
        RECT 12.605 2.480 12.615 2.754 ;
        RECT 12.615 2.480 12.625 2.744 ;
        RECT 12.625 2.480 12.635 2.734 ;
        RECT 12.635 2.480 12.645 2.724 ;
        RECT 12.645 2.480 12.655 2.714 ;
        RECT 12.655 2.480 12.665 2.704 ;
        RECT 12.665 2.480 12.675 2.694 ;
        RECT 12.675 2.480 12.685 2.684 ;
        RECT 12.685 2.480 12.695 2.674 ;
        RECT 12.695 2.480 12.705 2.664 ;
        RECT 12.705 2.480 12.715 2.654 ;
        RECT 12.715 2.480 12.721 2.650 ;
        RECT 12.560 2.525 12.570 2.799 ;
        RECT 12.570 2.515 12.580 2.789 ;
        RECT 12.580 2.505 12.590 2.779 ;
        RECT 12.590 2.495 12.600 2.769 ;
        RECT 12.600 2.485 12.606 2.765 ;
        RECT 12.445 2.640 12.455 2.810 ;
        RECT 12.455 2.630 12.465 2.810 ;
        RECT 12.465 2.620 12.475 2.810 ;
        RECT 12.475 2.610 12.485 2.810 ;
        RECT 12.485 2.600 12.495 2.810 ;
        RECT 12.495 2.590 12.505 2.810 ;
        RECT 12.505 2.580 12.515 2.810 ;
        RECT 12.515 2.570 12.525 2.810 ;
        RECT 12.525 2.560 12.535 2.810 ;
        RECT 12.535 2.550 12.545 2.810 ;
        RECT 12.545 2.540 12.555 2.810 ;
        RECT 12.555 2.530 12.561 2.810 ;
        RECT 10.570 0.975 10.580 1.209 ;
        RECT 10.580 0.985 10.590 1.209 ;
        RECT 10.590 0.995 10.600 1.209 ;
        RECT 10.600 1.005 10.610 1.209 ;
        RECT 10.610 1.015 10.620 1.209 ;
        RECT 10.620 1.025 10.630 1.209 ;
        RECT 10.630 1.035 10.640 1.209 ;
        RECT 10.640 1.040 10.646 1.210 ;
        RECT 10.505 0.910 10.515 1.144 ;
        RECT 10.515 0.920 10.525 1.154 ;
        RECT 10.525 0.930 10.535 1.164 ;
        RECT 10.535 0.940 10.545 1.174 ;
        RECT 10.545 0.950 10.555 1.184 ;
        RECT 10.555 0.960 10.565 1.194 ;
        RECT 10.565 0.965 10.571 1.205 ;
        RECT 10.430 0.900 10.440 1.070 ;
        RECT 10.440 0.900 10.450 1.080 ;
        RECT 10.450 0.900 10.460 1.090 ;
        RECT 10.460 0.900 10.470 1.100 ;
        RECT 10.470 0.900 10.480 1.110 ;
        RECT 10.480 0.900 10.490 1.120 ;
        RECT 10.490 0.900 10.500 1.130 ;
        RECT 10.500 0.900 10.506 1.140 ;
  END 
END FFSDNSRHDLXHT

MACRO FFSDNRHDLXHT
  CLASS  CORE ;
  FOREIGN FFSDNRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.120 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 3.680 1.525 4.170 2.010 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 12.780 1.060 13.020 1.360 ;
        RECT 12.810 1.060 13.020 2.445 ;
        RECT 12.780 1.980 13.020 2.445 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.580 0.860 11.910 1.470 ;
        RECT 11.580 1.300 12.250 1.470 ;
        RECT 12.080 1.300 12.250 2.215 ;
        RECT 11.675 2.045 12.250 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 8.030 1.610 8.510 2.010 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.110 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.435 -0.300 2.735 0.595 ;
        RECT 3.335 -0.300 3.635 0.595 ;
        RECT 6.035 -0.300 6.335 1.145 ;
        RECT 7.075 -0.300 7.375 0.595 ;
        RECT 8.105 -0.300 8.405 0.745 ;
        RECT 10.065 -0.300 10.365 0.525 ;
        RECT 11.195 -0.300 11.495 0.530 ;
        RECT 12.195 -0.300 12.495 0.745 ;
        RECT 0.000 -0.300 13.120 0.300 ;
    END
  END GND
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.450 2.510 2.620 3.990 ;
        RECT 3.340 2.890 3.510 3.990 ;
        RECT 6.035 3.195 6.335 3.990 ;
        RECT 8.165 3.195 8.465 3.990 ;
        RECT 10.165 2.810 10.465 3.990 ;
        RECT 12.195 2.810 12.495 3.990 ;
        RECT 0.000 3.390 13.120 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.555 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 2.965 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.530 0.865 1.720 1.185 ;
        RECT 2.005 0.775 2.175 1.035 ;
        RECT 1.530 0.865 2.175 1.035 ;
        RECT 2.005 0.775 4.600 0.945 ;
        RECT 4.365 0.565 4.600 0.945 ;
        RECT 4.430 0.565 4.600 2.280 ;
        RECT 5.130 0.900 5.300 2.280 ;
        RECT 6.235 1.675 6.535 1.865 ;
        RECT 5.130 1.695 6.535 1.865 ;
        RECT 5.755 1.325 6.055 1.515 ;
        RECT 6.650 0.775 6.885 1.495 ;
        RECT 5.755 1.325 6.885 1.495 ;
        RECT 6.715 0.775 6.885 2.215 ;
        RECT 6.715 2.045 7.255 2.215 ;
        RECT 7.630 0.480 7.800 0.945 ;
        RECT 6.650 0.775 7.800 0.945 ;
        RECT 2.795 1.985 3.050 2.285 ;
        RECT 2.795 1.125 2.990 2.285 ;
        RECT 2.880 1.985 3.050 2.710 ;
        RECT 2.795 1.125 3.125 1.295 ;
        RECT 2.880 2.540 3.900 2.710 ;
        RECT 3.730 2.540 3.900 3.015 ;
        RECT 8.460 2.745 8.630 3.015 ;
        RECT 3.730 2.845 8.630 3.015 ;
        RECT 8.460 2.745 9.045 2.915 ;
        RECT 3.170 1.525 3.495 1.825 ;
        RECT 3.325 1.125 3.495 2.360 ;
        RECT 3.325 2.190 4.250 2.360 ;
        RECT 3.325 1.125 4.165 1.295 ;
        RECT 4.080 2.190 4.250 2.635 ;
        RECT 4.780 0.535 4.950 2.635 ;
        RECT 4.780 0.535 5.575 0.705 ;
        RECT 8.105 2.395 8.275 2.635 ;
        RECT 4.080 2.465 8.275 2.635 ;
        RECT 8.845 1.330 9.015 2.565 ;
        RECT 8.825 1.330 9.125 1.500 ;
        RECT 8.105 2.395 9.720 2.565 ;
        RECT 9.550 2.395 9.720 2.695 ;
        RECT 7.065 1.600 7.810 1.770 ;
        RECT 7.640 1.125 7.810 2.280 ;
        RECT 7.640 1.125 8.475 1.295 ;
        RECT 9.690 0.605 9.860 0.945 ;
        RECT 8.975 0.605 9.860 0.775 ;
        RECT 9.690 0.775 11.335 0.945 ;
        RECT 11.165 0.775 11.335 1.515 ;
        RECT 8.860 0.605 8.870 0.879 ;
        RECT 8.870 0.605 8.880 0.869 ;
        RECT 8.880 0.605 8.890 0.859 ;
        RECT 8.890 0.605 8.900 0.849 ;
        RECT 8.900 0.605 8.910 0.839 ;
        RECT 8.910 0.605 8.920 0.829 ;
        RECT 8.920 0.605 8.930 0.819 ;
        RECT 8.930 0.605 8.940 0.809 ;
        RECT 8.940 0.605 8.950 0.799 ;
        RECT 8.950 0.605 8.960 0.789 ;
        RECT 8.960 0.605 8.970 0.779 ;
        RECT 8.970 0.605 8.976 0.775 ;
        RECT 8.645 0.820 8.655 1.094 ;
        RECT 8.655 0.810 8.665 1.084 ;
        RECT 8.665 0.800 8.675 1.074 ;
        RECT 8.675 0.790 8.685 1.064 ;
        RECT 8.685 0.780 8.695 1.054 ;
        RECT 8.695 0.770 8.705 1.044 ;
        RECT 8.705 0.760 8.715 1.034 ;
        RECT 8.715 0.750 8.725 1.024 ;
        RECT 8.725 0.740 8.735 1.014 ;
        RECT 8.735 0.730 8.745 1.004 ;
        RECT 8.745 0.720 8.755 0.994 ;
        RECT 8.755 0.710 8.765 0.984 ;
        RECT 8.765 0.700 8.775 0.974 ;
        RECT 8.775 0.690 8.785 0.964 ;
        RECT 8.785 0.680 8.795 0.954 ;
        RECT 8.795 0.670 8.805 0.944 ;
        RECT 8.805 0.660 8.815 0.934 ;
        RECT 8.815 0.650 8.825 0.924 ;
        RECT 8.825 0.640 8.835 0.914 ;
        RECT 8.835 0.630 8.845 0.904 ;
        RECT 8.845 0.620 8.855 0.894 ;
        RECT 8.855 0.610 8.861 0.890 ;
        RECT 8.475 0.990 8.485 1.294 ;
        RECT 8.485 0.980 8.495 1.294 ;
        RECT 8.495 0.970 8.505 1.294 ;
        RECT 8.505 0.960 8.515 1.294 ;
        RECT 8.515 0.950 8.525 1.294 ;
        RECT 8.525 0.940 8.535 1.294 ;
        RECT 8.535 0.930 8.545 1.294 ;
        RECT 8.545 0.920 8.555 1.294 ;
        RECT 8.555 0.910 8.565 1.294 ;
        RECT 8.565 0.900 8.575 1.294 ;
        RECT 8.575 0.890 8.585 1.294 ;
        RECT 8.585 0.880 8.595 1.294 ;
        RECT 8.595 0.870 8.605 1.294 ;
        RECT 8.605 0.860 8.615 1.294 ;
        RECT 8.615 0.850 8.625 1.294 ;
        RECT 8.625 0.840 8.635 1.294 ;
        RECT 8.635 0.830 8.645 1.294 ;
        RECT 10.615 1.125 10.985 1.495 ;
        RECT 9.855 1.325 10.985 1.495 ;
        RECT 10.815 1.125 10.985 1.865 ;
        RECT 11.150 1.695 11.320 2.280 ;
        RECT 11.600 1.675 11.900 1.865 ;
        RECT 10.815 1.695 11.900 1.865 ;
        RECT 9.115 0.955 9.475 1.125 ;
        RECT 9.305 0.955 9.475 2.215 ;
        RECT 9.220 2.045 9.520 2.215 ;
        RECT 9.305 1.675 10.635 1.845 ;
        RECT 10.465 1.675 10.635 2.630 ;
        RECT 12.430 1.610 12.600 2.630 ;
        RECT 10.465 2.460 12.600 2.630 ;
  END 
END FFSDNRHDLXHT

MACRO FFSDHQHD1XHT
  CLASS  CORE ;
  FOREIGN FFSDHQHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.300 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.800 0.720 12.200 1.360 ;
        RECT 11.950 0.720 12.200 2.895 ;
        RECT 11.800 1.980 12.200 2.895 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.240 1.175 1.775 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.575 0.380 2.010 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.045 ;
        RECT 2.545 -0.300 2.845 0.595 ;
        RECT 3.555 -0.300 3.855 0.595 ;
        RECT 4.495 -0.300 4.795 0.595 ;
        RECT 7.395 -0.300 7.695 0.595 ;
        RECT 8.430 -0.300 8.730 0.595 ;
        RECT 10.585 -0.300 10.755 0.805 ;
        RECT 11.280 -0.300 11.450 0.780 ;
        RECT 0.000 -0.300 12.300 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 4.495 1.470 5.010 2.020 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.365 1.435 2.775 2.020 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.540 0.955 3.990 ;
        RECT 2.555 2.470 2.730 3.990 ;
        RECT 3.555 2.745 3.855 3.990 ;
        RECT 4.460 2.745 4.760 3.990 ;
        RECT 7.410 2.890 7.710 3.990 ;
        RECT 8.465 2.970 8.765 3.990 ;
        RECT 10.415 2.610 10.585 3.990 ;
        RECT 11.305 2.635 11.605 3.990 ;
        RECT 0.000 3.390 12.300 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.010 0.340 1.395 ;
        RECT 0.170 2.190 0.340 2.490 ;
        RECT 0.170 1.225 0.730 1.395 ;
        RECT 0.560 1.225 0.730 2.360 ;
        RECT 0.170 2.190 0.730 2.360 ;
        RECT 1.355 1.510 1.525 2.125 ;
        RECT 0.560 1.955 1.525 2.125 ;
        RECT 1.355 1.510 1.630 1.810 ;
        RECT 3.390 1.605 3.560 1.905 ;
        RECT 3.390 1.605 4.285 1.775 ;
        RECT 3.985 1.125 4.285 2.215 ;
        RECT 5.080 1.125 5.655 1.295 ;
        RECT 5.485 1.125 5.655 2.215 ;
        RECT 5.350 2.045 5.655 2.215 ;
        RECT 5.485 1.430 5.720 1.730 ;
        RECT 1.640 2.330 1.810 2.970 ;
        RECT 1.810 1.025 1.980 2.515 ;
        RECT 1.640 2.330 1.980 2.515 ;
        RECT 2.485 0.775 2.655 1.195 ;
        RECT 1.575 1.025 2.655 1.195 ;
        RECT 2.485 0.775 6.095 0.945 ;
        RECT 5.925 0.775 6.095 2.320 ;
        RECT 6.625 1.060 6.795 2.320 ;
        RECT 7.635 1.585 7.805 2.210 ;
        RECT 6.625 2.040 7.805 2.210 ;
        RECT 7.635 1.585 8.030 1.755 ;
        RECT 7.285 1.220 7.455 1.820 ;
        RECT 8.050 1.970 8.220 2.280 ;
        RECT 7.985 1.125 8.525 1.390 ;
        RECT 7.285 1.220 8.525 1.390 ;
        RECT 8.355 1.125 8.525 2.140 ;
        RECT 8.050 1.970 8.525 2.140 ;
        RECT 8.355 1.515 8.655 1.815 ;
        RECT 3.005 1.125 3.185 2.565 ;
        RECT 3.005 2.135 3.240 2.565 ;
        RECT 3.005 1.125 3.305 1.370 ;
        RECT 5.170 2.395 5.470 2.670 ;
        RECT 3.005 2.395 5.470 2.565 ;
        RECT 6.275 0.650 6.445 2.670 ;
        RECT 5.170 2.500 6.445 2.670 ;
        RECT 6.965 0.650 7.135 0.945 ;
        RECT 6.275 0.650 7.135 0.830 ;
        RECT 6.965 0.775 9.045 0.945 ;
        RECT 8.875 0.775 9.045 1.610 ;
        RECT 8.875 1.310 9.440 1.610 ;
        RECT 6.740 2.530 7.040 2.705 ;
        RECT 8.835 1.925 9.005 2.700 ;
        RECT 6.740 2.530 9.005 2.700 ;
        RECT 9.645 0.985 9.815 2.095 ;
        RECT 8.835 1.925 9.815 2.095 ;
        RECT 9.645 0.985 9.945 1.285 ;
        RECT 9.420 2.435 9.590 3.075 ;
        RECT 9.995 1.550 10.165 2.605 ;
        RECT 9.420 2.435 10.165 2.605 ;
        RECT 9.420 0.570 10.365 0.740 ;
        RECT 10.195 0.570 10.365 1.720 ;
        RECT 9.995 1.550 11.190 1.720 ;
        RECT 10.380 1.915 10.550 2.215 ;
        RECT 10.665 1.125 11.560 1.295 ;
        RECT 11.370 1.125 11.560 2.215 ;
        RECT 10.380 2.045 11.560 2.215 ;
  END 
END FFSDHQHD1XHT

MACRO FFEDHQHDMXHT
  CLASS  CORE ;
  FOREIGN FFEDHQHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.890 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.415 0.720 11.585 2.280 ;
        RECT 11.415 1.675 11.790 2.280 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.865 1.265 1.130 2.015 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.585 2.015 ;
        RECT 0.285 2.645 1.365 2.815 ;
        RECT 1.195 2.645 1.365 3.210 ;
        RECT 1.195 3.040 2.075 3.210 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.735 ;
        RECT 2.415 -0.300 2.715 0.435 ;
        RECT 4.210 -0.300 4.510 0.435 ;
        RECT 6.960 -0.300 7.260 0.435 ;
        RECT 8.020 -0.300 8.320 0.435 ;
        RECT 9.890 -0.300 10.190 0.565 ;
        RECT 10.830 -0.300 11.130 1.055 ;
        RECT 0.000 -0.300 11.890 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 3.500 1.330 4.140 1.570 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.995 0.955 3.990 ;
        RECT 2.515 3.040 2.815 3.990 ;
        RECT 5.275 3.255 5.575 3.990 ;
        RECT 7.080 3.205 7.380 3.990 ;
        RECT 8.020 3.205 8.320 3.990 ;
        RECT 9.890 2.995 10.190 3.990 ;
        RECT 10.830 2.995 11.130 3.990 ;
        RECT 0.000 3.390 11.890 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.915 0.340 1.360 ;
        RECT 0.170 0.915 1.480 1.085 ;
        RECT 1.310 0.915 1.480 2.445 ;
        RECT 0.105 2.275 1.480 2.445 ;
        RECT 1.310 1.785 1.645 1.955 ;
        RECT 2.720 1.125 2.890 2.305 ;
        RECT 2.720 1.125 3.265 1.295 ;
        RECT 2.720 2.135 3.600 2.305 ;
        RECT 3.430 2.135 3.600 2.435 ;
        RECT 3.660 0.965 4.490 1.135 ;
        RECT 4.320 0.965 4.490 2.055 ;
        RECT 4.130 1.885 4.490 2.055 ;
        RECT 4.320 1.335 5.090 1.505 ;
        RECT 3.155 1.785 3.950 1.955 ;
        RECT 3.780 1.785 3.950 2.405 ;
        RECT 4.670 1.685 4.840 2.405 ;
        RECT 3.780 2.235 4.840 2.405 ;
        RECT 4.760 0.965 5.455 1.135 ;
        RECT 5.195 1.685 5.365 2.120 ;
        RECT 5.275 0.965 5.455 1.865 ;
        RECT 4.670 1.685 5.455 1.865 ;
        RECT 5.275 1.270 5.510 1.570 ;
        RECT 1.660 1.060 1.995 1.360 ;
        RECT 1.825 1.060 1.995 2.785 ;
        RECT 1.660 2.135 1.995 2.785 ;
        RECT 4.935 2.575 5.715 2.725 ;
        RECT 4.945 2.565 4.975 2.785 ;
        RECT 4.925 2.585 5.715 2.725 ;
        RECT 1.660 2.615 4.975 2.785 ;
        RECT 1.660 2.615 4.985 2.775 ;
        RECT 1.660 2.615 4.995 2.765 ;
        RECT 1.660 2.615 5.005 2.755 ;
        RECT 1.660 2.615 5.015 2.745 ;
        RECT 1.660 2.615 5.025 2.735 ;
        RECT 4.955 2.555 5.715 2.725 ;
        RECT 4.915 2.595 5.715 2.725 ;
        RECT 5.545 2.155 5.715 2.725 ;
        RECT 4.905 2.605 5.715 2.725 ;
        RECT 5.705 0.965 5.875 2.325 ;
        RECT 5.640 0.965 5.940 1.135 ;
        RECT 5.545 2.155 5.940 2.325 ;
        RECT 6.225 0.965 6.395 2.325 ;
        RECT 6.160 0.965 6.460 1.135 ;
        RECT 6.160 2.155 6.460 2.325 ;
        RECT 6.225 1.785 7.630 1.955 ;
        RECT 7.575 0.965 7.745 1.605 ;
        RECT 7.510 0.965 7.810 1.135 ;
        RECT 7.810 1.435 7.980 2.325 ;
        RECT 7.510 2.155 7.980 2.325 ;
        RECT 6.840 1.435 8.530 1.605 ;
        RECT 3.365 2.965 5.055 3.135 ;
        RECT 5.115 2.905 5.135 3.135 ;
        RECT 5.195 2.905 5.730 3.075 ;
        RECT 6.500 2.855 6.800 3.195 ;
        RECT 5.930 3.025 6.800 3.195 ;
        RECT 6.500 2.855 9.010 3.025 ;
        RECT 8.710 2.855 9.010 3.195 ;
        RECT 5.850 2.955 5.860 3.195 ;
        RECT 5.860 2.965 5.870 3.195 ;
        RECT 5.870 2.975 5.880 3.195 ;
        RECT 5.880 2.985 5.890 3.195 ;
        RECT 5.890 2.995 5.900 3.195 ;
        RECT 5.900 3.005 5.910 3.195 ;
        RECT 5.910 3.015 5.920 3.195 ;
        RECT 5.920 3.025 5.930 3.195 ;
        RECT 5.810 2.915 5.820 3.155 ;
        RECT 5.820 2.925 5.830 3.165 ;
        RECT 5.830 2.935 5.840 3.175 ;
        RECT 5.840 2.945 5.850 3.185 ;
        RECT 5.730 2.905 5.740 3.075 ;
        RECT 5.740 2.905 5.750 3.085 ;
        RECT 5.750 2.905 5.760 3.095 ;
        RECT 5.760 2.905 5.770 3.105 ;
        RECT 5.770 2.905 5.780 3.115 ;
        RECT 5.780 2.905 5.790 3.125 ;
        RECT 5.790 2.905 5.800 3.135 ;
        RECT 5.800 2.905 5.810 3.145 ;
        RECT 5.135 2.905 5.145 3.125 ;
        RECT 5.145 2.905 5.155 3.115 ;
        RECT 5.155 2.905 5.165 3.105 ;
        RECT 5.165 2.905 5.175 3.095 ;
        RECT 5.175 2.905 5.185 3.085 ;
        RECT 5.185 2.905 5.195 3.075 ;
        RECT 5.055 2.965 5.065 3.135 ;
        RECT 5.065 2.955 5.075 3.135 ;
        RECT 5.075 2.945 5.085 3.135 ;
        RECT 5.085 2.935 5.095 3.135 ;
        RECT 5.095 2.925 5.105 3.135 ;
        RECT 5.105 2.915 5.115 3.135 ;
        RECT 5.980 2.505 6.300 2.815 ;
        RECT 8.590 1.785 8.760 2.675 ;
        RECT 8.775 1.315 8.945 1.955 ;
        RECT 8.590 1.785 8.945 1.955 ;
        RECT 8.710 1.315 9.010 1.485 ;
        RECT 5.980 2.505 9.360 2.675 ;
        RECT 9.190 2.505 9.360 3.195 ;
        RECT 9.190 3.025 9.490 3.195 ;
        RECT 2.370 0.615 2.540 1.820 ;
        RECT 8.545 0.575 8.715 0.785 ;
        RECT 2.370 0.615 8.715 0.785 ;
        RECT 8.545 0.575 9.710 0.745 ;
        RECT 9.540 0.575 9.710 1.755 ;
        RECT 9.540 1.585 10.555 1.755 ;
        RECT 10.385 0.880 10.555 2.465 ;
        RECT 10.320 2.295 10.620 2.465 ;
        RECT 8.940 0.945 9.360 1.115 ;
        RECT 9.190 0.945 9.360 2.325 ;
        RECT 8.940 2.155 10.115 2.325 ;
        RECT 9.935 2.155 10.115 2.815 ;
        RECT 11.000 1.520 11.170 2.815 ;
        RECT 9.935 2.645 11.170 2.815 ;
  END 
END FFEDHQHDMXHT

MACRO FFEDCRHD2XHT
  CLASS  CORE ;
  FOREIGN FFEDCRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.170 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.210 0.720 14.380 2.960 ;
        RECT 14.210 1.740 14.755 1.950 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.170 0.720 13.340 2.280 ;
        RECT 13.170 0.720 13.430 1.230 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.115 1.265 2.425 1.795 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.195 2.560 0.835 2.770 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.605 1.625 2.780 2.430 ;
        RECT 2.560 2.085 2.780 2.430 ;
        RECT 2.605 1.625 2.980 1.795 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.685 ;
        RECT 2.425 -0.300 2.725 0.745 ;
        RECT 3.470 -0.300 3.770 0.595 ;
        RECT 4.350 -0.300 4.650 0.595 ;
        RECT 5.420 -0.300 5.720 0.595 ;
        RECT 6.335 -0.300 6.635 0.595 ;
        RECT 8.505 -0.300 8.675 0.620 ;
        RECT 9.630 -0.300 9.800 0.700 ;
        RECT 11.620 -0.300 11.790 1.060 ;
        RECT 12.585 -0.300 12.885 1.055 ;
        RECT 13.625 -0.300 13.925 1.055 ;
        RECT 14.665 -0.300 14.965 1.055 ;
        RECT 0.000 -0.300 15.170 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 4.870 1.545 5.300 1.950 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 2.960 0.835 3.990 ;
        RECT 2.425 2.970 2.725 3.990 ;
        RECT 3.285 2.970 3.585 3.990 ;
        RECT 5.305 2.830 5.605 3.990 ;
        RECT 6.345 3.170 6.645 3.990 ;
        RECT 8.410 3.170 8.710 3.990 ;
        RECT 9.565 3.170 9.865 3.990 ;
        RECT 11.525 2.825 11.825 3.990 ;
        RECT 12.585 2.975 12.885 3.990 ;
        RECT 13.625 2.975 13.925 3.990 ;
        RECT 14.665 2.295 14.965 3.990 ;
        RECT 0.000 3.390 15.170 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.010 0.340 2.300 ;
        RECT 0.170 1.585 1.340 1.755 ;
        RECT 1.170 0.605 1.340 3.040 ;
        RECT 1.170 0.605 1.525 0.775 ;
        RECT 1.170 2.870 1.940 3.040 ;
        RECT 1.770 2.870 1.940 3.170 ;
        RECT 2.960 2.000 3.130 2.300 ;
        RECT 2.900 1.125 3.520 1.295 ;
        RECT 3.350 1.125 3.520 2.170 ;
        RECT 2.960 2.000 3.520 2.170 ;
        RECT 3.350 1.580 3.820 1.750 ;
        RECT 1.520 1.010 1.740 1.310 ;
        RECT 1.570 1.010 1.740 2.640 ;
        RECT 2.160 2.460 2.330 2.780 ;
        RECT 1.570 2.460 2.330 2.640 ;
        RECT 2.160 2.610 3.990 2.780 ;
        RECT 3.810 2.610 3.990 3.045 ;
        RECT 3.810 2.875 4.325 3.045 ;
        RECT 4.785 2.130 5.390 2.300 ;
        RECT 4.870 1.125 5.490 1.295 ;
        RECT 5.480 1.125 5.490 2.300 ;
        RECT 5.660 1.540 5.765 1.840 ;
        RECT 5.490 1.125 5.500 2.289 ;
        RECT 5.500 1.125 5.510 2.279 ;
        RECT 5.510 1.125 5.520 2.269 ;
        RECT 5.520 1.125 5.530 2.259 ;
        RECT 5.530 1.125 5.540 2.249 ;
        RECT 5.540 1.125 5.550 2.239 ;
        RECT 5.550 1.125 5.560 2.229 ;
        RECT 5.560 1.125 5.570 2.219 ;
        RECT 5.570 1.125 5.580 2.209 ;
        RECT 5.580 1.125 5.590 2.199 ;
        RECT 5.590 1.125 5.600 2.189 ;
        RECT 5.600 1.125 5.610 2.179 ;
        RECT 5.610 1.125 5.620 2.169 ;
        RECT 5.620 1.125 5.630 2.159 ;
        RECT 5.630 1.125 5.640 2.149 ;
        RECT 5.640 1.125 5.650 2.139 ;
        RECT 5.650 1.125 5.660 2.129 ;
        RECT 5.390 2.130 5.400 2.300 ;
        RECT 5.400 2.120 5.410 2.300 ;
        RECT 5.410 2.110 5.420 2.300 ;
        RECT 5.420 2.100 5.430 2.300 ;
        RECT 5.430 2.090 5.440 2.300 ;
        RECT 5.440 2.080 5.450 2.300 ;
        RECT 5.450 2.070 5.460 2.300 ;
        RECT 5.460 2.060 5.470 2.300 ;
        RECT 5.470 2.050 5.480 2.300 ;
        RECT 3.860 1.125 4.440 1.295 ;
        RECT 4.270 1.125 4.440 2.650 ;
        RECT 5.635 2.440 5.705 2.650 ;
        RECT 5.625 2.450 6.765 2.595 ;
        RECT 5.645 2.430 5.705 2.650 ;
        RECT 5.615 2.460 6.765 2.595 ;
        RECT 4.270 2.480 5.705 2.650 ;
        RECT 4.270 2.480 5.715 2.639 ;
        RECT 4.270 2.480 5.725 2.629 ;
        RECT 4.270 2.480 5.735 2.619 ;
        RECT 4.270 2.480 5.745 2.609 ;
        RECT 4.270 2.480 5.755 2.599 ;
        RECT 5.650 2.425 6.765 2.595 ;
        RECT 5.605 2.470 6.765 2.595 ;
        RECT 6.595 1.580 6.765 2.595 ;
        RECT 7.450 1.200 7.620 2.290 ;
        RECT 7.450 1.200 7.795 1.370 ;
        RECT 7.450 2.120 8.545 2.290 ;
        RECT 8.840 1.595 8.925 1.895 ;
        RECT 8.755 1.595 8.765 1.969 ;
        RECT 8.765 1.595 8.775 1.959 ;
        RECT 8.775 1.595 8.785 1.949 ;
        RECT 8.785 1.595 8.795 1.939 ;
        RECT 8.795 1.595 8.805 1.929 ;
        RECT 8.805 1.595 8.815 1.919 ;
        RECT 8.815 1.595 8.825 1.909 ;
        RECT 8.825 1.595 8.835 1.899 ;
        RECT 8.835 1.595 8.841 1.895 ;
        RECT 8.725 1.735 8.735 1.999 ;
        RECT 8.735 1.725 8.745 1.989 ;
        RECT 8.745 1.715 8.755 1.979 ;
        RECT 8.545 1.915 8.555 2.289 ;
        RECT 8.555 1.905 8.565 2.289 ;
        RECT 8.565 1.895 8.575 2.289 ;
        RECT 8.575 1.885 8.585 2.289 ;
        RECT 8.585 1.875 8.595 2.289 ;
        RECT 8.595 1.865 8.605 2.289 ;
        RECT 8.605 1.855 8.615 2.289 ;
        RECT 8.615 1.845 8.625 2.289 ;
        RECT 8.625 1.835 8.635 2.289 ;
        RECT 8.635 1.825 8.645 2.289 ;
        RECT 8.645 1.815 8.655 2.289 ;
        RECT 8.655 1.805 8.665 2.289 ;
        RECT 8.665 1.795 8.675 2.289 ;
        RECT 8.675 1.785 8.685 2.289 ;
        RECT 8.685 1.775 8.695 2.289 ;
        RECT 8.695 1.765 8.705 2.289 ;
        RECT 8.705 1.755 8.715 2.289 ;
        RECT 8.715 1.745 8.725 2.289 ;
        RECT 8.295 1.165 8.465 1.740 ;
        RECT 8.165 1.570 8.465 1.740 ;
        RECT 8.295 1.165 9.290 1.335 ;
        RECT 9.120 1.165 9.290 2.290 ;
        RECT 8.960 2.120 9.290 2.290 ;
        RECT 9.120 1.570 10.015 1.740 ;
        RECT 5.830 2.820 6.105 3.195 ;
        RECT 7.790 2.820 8.090 3.005 ;
        RECT 5.830 2.820 10.000 2.990 ;
        RECT 10.310 3.040 11.155 3.210 ;
        RECT 10.220 2.960 10.230 3.210 ;
        RECT 10.230 2.970 10.240 3.210 ;
        RECT 10.240 2.980 10.250 3.210 ;
        RECT 10.250 2.990 10.260 3.210 ;
        RECT 10.260 3.000 10.270 3.210 ;
        RECT 10.270 3.010 10.280 3.210 ;
        RECT 10.280 3.020 10.290 3.210 ;
        RECT 10.290 3.030 10.300 3.210 ;
        RECT 10.300 3.040 10.310 3.210 ;
        RECT 10.090 2.830 10.100 3.080 ;
        RECT 10.100 2.840 10.110 3.090 ;
        RECT 10.110 2.850 10.120 3.100 ;
        RECT 10.120 2.860 10.130 3.110 ;
        RECT 10.130 2.870 10.140 3.120 ;
        RECT 10.140 2.880 10.150 3.130 ;
        RECT 10.150 2.890 10.160 3.140 ;
        RECT 10.160 2.900 10.170 3.150 ;
        RECT 10.170 2.910 10.180 3.160 ;
        RECT 10.180 2.920 10.190 3.170 ;
        RECT 10.190 2.930 10.200 3.180 ;
        RECT 10.200 2.940 10.210 3.190 ;
        RECT 10.210 2.950 10.220 3.200 ;
        RECT 10.000 2.820 10.010 2.990 ;
        RECT 10.010 2.820 10.020 3.000 ;
        RECT 10.020 2.820 10.030 3.010 ;
        RECT 10.030 2.820 10.040 3.020 ;
        RECT 10.040 2.820 10.050 3.030 ;
        RECT 10.050 2.820 10.060 3.040 ;
        RECT 10.060 2.820 10.070 3.050 ;
        RECT 10.070 2.820 10.080 3.060 ;
        RECT 10.080 2.820 10.090 3.070 ;
        RECT 5.805 2.845 5.815 3.195 ;
        RECT 5.815 2.835 5.825 3.195 ;
        RECT 5.825 2.825 5.831 3.195 ;
        RECT 5.985 1.125 6.155 2.225 ;
        RECT 5.855 2.055 6.155 2.225 ;
        RECT 5.860 1.125 7.020 1.295 ;
        RECT 6.965 1.125 7.020 2.125 ;
        RECT 7.135 1.825 7.270 2.640 ;
        RECT 7.635 0.830 7.935 1.020 ;
        RECT 7.370 0.850 7.935 1.020 ;
        RECT 10.225 1.315 10.255 2.640 ;
        RECT 7.135 2.470 10.255 2.640 ;
        RECT 10.345 1.315 10.395 2.730 ;
        RECT 10.345 1.315 10.490 1.615 ;
        RECT 10.475 2.560 11.195 2.730 ;
        RECT 10.395 2.490 10.405 2.730 ;
        RECT 10.405 2.500 10.415 2.730 ;
        RECT 10.415 2.510 10.425 2.730 ;
        RECT 10.425 2.520 10.435 2.730 ;
        RECT 10.435 2.530 10.445 2.730 ;
        RECT 10.445 2.540 10.455 2.730 ;
        RECT 10.455 2.550 10.465 2.730 ;
        RECT 10.465 2.560 10.475 2.730 ;
        RECT 10.255 1.315 10.265 2.639 ;
        RECT 10.265 1.315 10.275 2.649 ;
        RECT 10.275 1.315 10.285 2.659 ;
        RECT 10.285 1.315 10.295 2.669 ;
        RECT 10.295 1.315 10.305 2.679 ;
        RECT 10.305 1.315 10.315 2.689 ;
        RECT 10.315 1.315 10.325 2.699 ;
        RECT 10.325 1.315 10.335 2.709 ;
        RECT 10.335 1.315 10.345 2.719 ;
        RECT 7.295 0.850 7.305 1.084 ;
        RECT 7.305 0.850 7.315 1.074 ;
        RECT 7.315 0.850 7.325 1.064 ;
        RECT 7.325 0.850 7.335 1.054 ;
        RECT 7.335 0.850 7.345 1.044 ;
        RECT 7.345 0.850 7.355 1.034 ;
        RECT 7.355 0.850 7.365 1.024 ;
        RECT 7.365 0.850 7.371 1.020 ;
        RECT 7.135 1.010 7.145 1.244 ;
        RECT 7.145 1.000 7.155 1.234 ;
        RECT 7.155 0.990 7.165 1.224 ;
        RECT 7.165 0.980 7.175 1.214 ;
        RECT 7.175 0.970 7.185 1.204 ;
        RECT 7.185 0.960 7.195 1.194 ;
        RECT 7.195 0.950 7.205 1.184 ;
        RECT 7.205 0.940 7.215 1.174 ;
        RECT 7.215 0.930 7.225 1.164 ;
        RECT 7.225 0.920 7.235 1.154 ;
        RECT 7.235 0.910 7.245 1.144 ;
        RECT 7.245 0.900 7.255 1.134 ;
        RECT 7.255 0.890 7.265 1.124 ;
        RECT 7.265 0.880 7.275 1.114 ;
        RECT 7.275 0.870 7.285 1.104 ;
        RECT 7.285 0.860 7.295 1.094 ;
        RECT 7.100 1.045 7.110 2.639 ;
        RECT 7.110 1.035 7.120 2.639 ;
        RECT 7.120 1.025 7.130 2.639 ;
        RECT 7.130 1.015 7.136 2.639 ;
        RECT 7.020 1.125 7.030 2.125 ;
        RECT 7.030 1.115 7.040 2.125 ;
        RECT 7.040 1.105 7.050 2.125 ;
        RECT 7.050 1.095 7.060 2.125 ;
        RECT 7.060 1.085 7.070 2.125 ;
        RECT 7.070 1.075 7.080 2.125 ;
        RECT 7.080 1.065 7.090 2.125 ;
        RECT 7.090 1.055 7.100 2.125 ;
        RECT 2.990 0.490 3.290 0.945 ;
        RECT 2.990 0.775 6.865 0.945 ;
        RECT 7.235 0.480 8.015 0.650 ;
        RECT 8.285 0.810 9.390 0.980 ;
        RECT 9.470 0.810 9.475 1.060 ;
        RECT 10.145 0.615 10.315 1.060 ;
        RECT 9.545 0.880 10.315 1.060 ;
        RECT 10.145 0.615 11.420 0.785 ;
        RECT 11.250 0.500 11.420 1.415 ;
        RECT 11.250 1.245 12.395 1.415 ;
        RECT 12.140 1.060 12.310 1.415 ;
        RECT 12.225 1.245 12.395 2.285 ;
        RECT 12.075 2.115 12.395 2.285 ;
        RECT 12.225 1.540 12.990 1.840 ;
        RECT 9.475 0.820 9.485 1.060 ;
        RECT 9.485 0.830 9.495 1.060 ;
        RECT 9.495 0.840 9.505 1.060 ;
        RECT 9.505 0.850 9.515 1.060 ;
        RECT 9.515 0.860 9.525 1.060 ;
        RECT 9.525 0.870 9.535 1.060 ;
        RECT 9.535 0.880 9.545 1.060 ;
        RECT 9.390 0.810 9.400 0.980 ;
        RECT 9.400 0.810 9.410 0.990 ;
        RECT 9.410 0.810 9.420 1.000 ;
        RECT 9.420 0.810 9.430 1.010 ;
        RECT 9.430 0.810 9.440 1.020 ;
        RECT 9.440 0.810 9.450 1.030 ;
        RECT 9.450 0.810 9.460 1.040 ;
        RECT 9.460 0.810 9.470 1.050 ;
        RECT 8.115 0.515 8.125 0.979 ;
        RECT 8.125 0.525 8.135 0.979 ;
        RECT 8.135 0.535 8.145 0.979 ;
        RECT 8.145 0.545 8.155 0.979 ;
        RECT 8.155 0.555 8.165 0.979 ;
        RECT 8.165 0.565 8.175 0.979 ;
        RECT 8.175 0.575 8.185 0.979 ;
        RECT 8.185 0.585 8.195 0.979 ;
        RECT 8.195 0.595 8.205 0.979 ;
        RECT 8.205 0.605 8.215 0.979 ;
        RECT 8.215 0.615 8.225 0.979 ;
        RECT 8.225 0.625 8.235 0.979 ;
        RECT 8.235 0.635 8.245 0.979 ;
        RECT 8.245 0.645 8.255 0.979 ;
        RECT 8.255 0.655 8.265 0.979 ;
        RECT 8.265 0.665 8.275 0.979 ;
        RECT 8.275 0.675 8.285 0.979 ;
        RECT 8.090 0.490 8.100 0.724 ;
        RECT 8.100 0.500 8.110 0.734 ;
        RECT 8.110 0.505 8.116 0.745 ;
        RECT 8.015 0.480 8.025 0.650 ;
        RECT 8.025 0.480 8.035 0.660 ;
        RECT 8.035 0.480 8.045 0.670 ;
        RECT 8.045 0.480 8.055 0.680 ;
        RECT 8.055 0.480 8.065 0.690 ;
        RECT 8.065 0.480 8.075 0.700 ;
        RECT 8.075 0.480 8.085 0.710 ;
        RECT 8.085 0.480 8.091 0.720 ;
        RECT 7.160 0.480 7.170 0.714 ;
        RECT 7.170 0.480 7.180 0.704 ;
        RECT 7.180 0.480 7.190 0.694 ;
        RECT 7.190 0.480 7.200 0.684 ;
        RECT 7.200 0.480 7.210 0.674 ;
        RECT 7.210 0.480 7.220 0.664 ;
        RECT 7.220 0.480 7.230 0.654 ;
        RECT 7.230 0.480 7.236 0.650 ;
        RECT 6.940 0.700 6.950 0.934 ;
        RECT 6.950 0.690 6.960 0.924 ;
        RECT 6.960 0.680 6.970 0.914 ;
        RECT 6.970 0.670 6.980 0.904 ;
        RECT 6.980 0.660 6.990 0.894 ;
        RECT 6.990 0.650 7.000 0.884 ;
        RECT 7.000 0.640 7.010 0.874 ;
        RECT 7.010 0.630 7.020 0.864 ;
        RECT 7.020 0.620 7.030 0.854 ;
        RECT 7.030 0.610 7.040 0.844 ;
        RECT 7.040 0.600 7.050 0.834 ;
        RECT 7.050 0.590 7.060 0.824 ;
        RECT 7.060 0.580 7.070 0.814 ;
        RECT 7.070 0.570 7.080 0.804 ;
        RECT 7.080 0.560 7.090 0.794 ;
        RECT 7.090 0.550 7.100 0.784 ;
        RECT 7.100 0.540 7.110 0.774 ;
        RECT 7.110 0.530 7.120 0.764 ;
        RECT 7.120 0.520 7.130 0.754 ;
        RECT 7.130 0.510 7.140 0.744 ;
        RECT 7.140 0.500 7.150 0.734 ;
        RECT 7.150 0.490 7.160 0.724 ;
        RECT 6.865 0.775 6.875 0.945 ;
        RECT 6.875 0.765 6.885 0.945 ;
        RECT 6.885 0.755 6.895 0.945 ;
        RECT 6.895 0.745 6.905 0.945 ;
        RECT 6.905 0.735 6.915 0.945 ;
        RECT 6.915 0.725 6.925 0.945 ;
        RECT 6.925 0.715 6.935 0.945 ;
        RECT 6.935 0.705 6.941 0.945 ;
        RECT 10.515 0.965 10.850 1.135 ;
        RECT 10.670 0.965 10.850 2.330 ;
        RECT 10.590 2.030 10.850 2.330 ;
        RECT 11.445 1.700 11.615 2.645 ;
        RECT 10.670 1.700 12.045 1.870 ;
        RECT 13.840 1.545 14.010 2.645 ;
        RECT 11.445 2.475 14.010 2.645 ;
  END 
END FFEDCRHD2XHT

MACRO FFDSHQHDMXHT
  CLASS  CORE ;
  FOREIGN FFDSHQHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.430 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.025 0.630 9.330 2.280 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.600 2.560 2.050 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.995 ;
        RECT 2.175 -0.300 2.475 1.230 ;
        RECT 4.025 -0.300 4.325 1.065 ;
        RECT 5.345 -0.300 5.645 0.485 ;
        RECT 7.235 -0.300 7.535 0.745 ;
        RECT 8.505 -0.300 8.805 0.715 ;
        RECT 0.000 -0.300 9.430 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.870 1.260 1.130 1.785 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.610 0.710 4.840 1.200 ;
        RECT 4.670 0.710 4.840 1.845 ;
        RECT 4.670 1.675 5.065 1.845 ;
        RECT 5.945 0.545 6.115 0.880 ;
        RECT 4.610 0.710 6.115 0.880 ;
        RECT 5.945 0.545 7.035 0.715 ;
        RECT 4.610 0.710 7.035 0.715 ;
        RECT 6.865 0.545 7.035 1.095 ;
        RECT 7.715 0.755 7.885 1.095 ;
        RECT 6.865 0.925 7.885 1.095 ;
        RECT 7.715 0.755 8.235 0.925 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 1.980 0.340 3.990 ;
        RECT 2.145 3.215 2.445 3.990 ;
        RECT 4.035 3.095 4.335 3.990 ;
        RECT 5.135 3.095 5.435 3.990 ;
        RECT 7.235 2.745 7.535 3.990 ;
        RECT 8.570 2.310 8.805 3.990 ;
        RECT 0.000 3.390 9.430 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.000 1.965 1.170 2.215 ;
        RECT 0.870 2.045 1.170 2.215 ;
        RECT 1.145 0.825 1.480 0.995 ;
        RECT 1.000 1.965 1.480 2.135 ;
        RECT 1.310 0.825 1.480 2.135 ;
        RECT 1.310 1.610 1.540 1.910 ;
        RECT 3.115 2.165 3.285 2.335 ;
        RECT 3.130 0.995 3.300 1.495 ;
        RECT 3.130 1.325 3.415 1.495 ;
        RECT 3.315 1.325 3.415 2.335 ;
        RECT 3.485 1.325 4.150 1.495 ;
        RECT 4.320 1.405 4.330 1.865 ;
        RECT 4.330 1.415 4.340 1.865 ;
        RECT 4.340 1.425 4.350 1.865 ;
        RECT 4.350 1.435 4.360 1.865 ;
        RECT 4.360 1.445 4.370 1.865 ;
        RECT 4.370 1.455 4.380 1.865 ;
        RECT 4.380 1.465 4.390 1.865 ;
        RECT 4.390 1.475 4.400 1.865 ;
        RECT 4.400 1.485 4.410 1.865 ;
        RECT 4.410 1.495 4.420 1.865 ;
        RECT 4.420 1.505 4.430 1.865 ;
        RECT 4.430 1.515 4.440 1.865 ;
        RECT 4.440 1.525 4.450 1.865 ;
        RECT 4.450 1.535 4.460 1.865 ;
        RECT 4.460 1.545 4.470 1.865 ;
        RECT 4.470 1.555 4.480 1.865 ;
        RECT 4.480 1.565 4.490 1.865 ;
        RECT 4.250 1.335 4.260 1.595 ;
        RECT 4.260 1.345 4.270 1.605 ;
        RECT 4.270 1.355 4.280 1.615 ;
        RECT 4.280 1.365 4.290 1.625 ;
        RECT 4.290 1.375 4.300 1.635 ;
        RECT 4.300 1.385 4.310 1.645 ;
        RECT 4.310 1.395 4.320 1.655 ;
        RECT 4.150 1.325 4.160 1.495 ;
        RECT 4.160 1.325 4.170 1.505 ;
        RECT 4.170 1.325 4.180 1.515 ;
        RECT 4.180 1.325 4.190 1.525 ;
        RECT 4.190 1.325 4.200 1.535 ;
        RECT 4.200 1.325 4.210 1.545 ;
        RECT 4.210 1.325 4.220 1.555 ;
        RECT 4.220 1.325 4.230 1.565 ;
        RECT 4.230 1.325 4.240 1.575 ;
        RECT 4.240 1.325 4.250 1.585 ;
        RECT 3.415 1.325 3.425 2.325 ;
        RECT 3.425 1.325 3.435 2.315 ;
        RECT 3.435 1.325 3.445 2.305 ;
        RECT 3.445 1.325 3.455 2.295 ;
        RECT 3.455 1.325 3.465 2.285 ;
        RECT 3.465 1.325 3.475 2.275 ;
        RECT 3.475 1.325 3.485 2.265 ;
        RECT 3.285 2.165 3.295 2.335 ;
        RECT 3.295 2.155 3.305 2.335 ;
        RECT 3.305 2.145 3.315 2.335 ;
        RECT 3.775 1.675 4.075 2.215 ;
        RECT 5.020 1.060 5.190 1.360 ;
        RECT 5.020 1.190 5.760 1.360 ;
        RECT 5.590 1.190 5.760 2.215 ;
        RECT 3.770 2.045 5.760 2.215 ;
        RECT 0.170 1.060 0.340 1.790 ;
        RECT 0.170 1.620 0.690 1.790 ;
        RECT 0.520 1.620 0.690 2.565 ;
        RECT 0.520 2.395 1.230 2.565 ;
        RECT 1.060 2.395 1.230 3.035 ;
        RECT 1.060 2.865 3.640 3.035 ;
        RECT 5.615 2.745 5.785 3.035 ;
        RECT 3.835 2.745 5.785 2.915 ;
        RECT 5.615 2.865 6.335 3.035 ;
        RECT 3.760 2.745 3.770 2.979 ;
        RECT 3.770 2.745 3.780 2.969 ;
        RECT 3.780 2.745 3.790 2.959 ;
        RECT 3.790 2.745 3.800 2.949 ;
        RECT 3.800 2.745 3.810 2.939 ;
        RECT 3.810 2.745 3.820 2.929 ;
        RECT 3.820 2.745 3.830 2.919 ;
        RECT 3.830 2.745 3.836 2.915 ;
        RECT 3.715 2.790 3.725 3.024 ;
        RECT 3.725 2.780 3.735 3.014 ;
        RECT 3.735 2.770 3.745 3.004 ;
        RECT 3.745 2.760 3.755 2.994 ;
        RECT 3.755 2.750 3.761 2.990 ;
        RECT 3.640 2.865 3.650 3.035 ;
        RECT 3.650 2.855 3.660 3.035 ;
        RECT 3.660 2.845 3.670 3.035 ;
        RECT 3.670 2.835 3.680 3.035 ;
        RECT 3.680 2.825 3.690 3.035 ;
        RECT 3.690 2.815 3.700 3.035 ;
        RECT 3.700 2.805 3.710 3.035 ;
        RECT 3.710 2.795 3.716 3.035 ;
        RECT 1.720 0.995 1.890 2.685 ;
        RECT 1.440 2.350 1.890 2.685 ;
        RECT 2.765 0.525 2.935 2.685 ;
        RECT 2.765 1.795 3.135 1.965 ;
        RECT 1.440 2.515 3.490 2.685 ;
        RECT 2.765 0.525 3.595 0.695 ;
        RECT 5.965 1.265 6.135 2.685 ;
        RECT 3.685 2.395 6.135 2.565 ;
        RECT 5.965 1.265 6.335 1.435 ;
        RECT 5.965 2.515 6.780 2.685 ;
        RECT 6.610 2.515 6.780 2.890 ;
        RECT 3.610 2.395 3.620 2.629 ;
        RECT 3.620 2.395 3.630 2.619 ;
        RECT 3.630 2.395 3.640 2.609 ;
        RECT 3.640 2.395 3.650 2.599 ;
        RECT 3.650 2.395 3.660 2.589 ;
        RECT 3.660 2.395 3.670 2.579 ;
        RECT 3.670 2.395 3.680 2.569 ;
        RECT 3.680 2.395 3.686 2.565 ;
        RECT 3.565 2.440 3.575 2.674 ;
        RECT 3.575 2.430 3.585 2.664 ;
        RECT 3.585 2.420 3.595 2.654 ;
        RECT 3.595 2.410 3.605 2.644 ;
        RECT 3.605 2.400 3.611 2.640 ;
        RECT 3.490 2.515 3.500 2.685 ;
        RECT 3.500 2.505 3.510 2.685 ;
        RECT 3.510 2.495 3.520 2.685 ;
        RECT 3.520 2.485 3.530 2.685 ;
        RECT 3.530 2.475 3.540 2.685 ;
        RECT 3.540 2.465 3.550 2.685 ;
        RECT 3.550 2.455 3.560 2.685 ;
        RECT 3.560 2.445 3.566 2.685 ;
        RECT 7.870 1.455 8.040 2.215 ;
        RECT 7.490 2.045 8.040 2.215 ;
        RECT 8.065 1.125 8.235 1.625 ;
        RECT 7.870 1.455 8.235 1.625 ;
        RECT 8.065 1.125 8.415 1.295 ;
        RECT 7.320 1.885 7.330 2.215 ;
        RECT 7.330 1.895 7.340 2.215 ;
        RECT 7.340 1.905 7.350 2.215 ;
        RECT 7.350 1.915 7.360 2.215 ;
        RECT 7.360 1.925 7.370 2.215 ;
        RECT 7.370 1.935 7.380 2.215 ;
        RECT 7.380 1.945 7.390 2.215 ;
        RECT 7.390 1.955 7.400 2.215 ;
        RECT 7.400 1.965 7.410 2.215 ;
        RECT 7.410 1.975 7.420 2.215 ;
        RECT 7.420 1.985 7.430 2.215 ;
        RECT 7.430 1.995 7.440 2.215 ;
        RECT 7.440 2.005 7.450 2.215 ;
        RECT 7.450 2.015 7.460 2.215 ;
        RECT 7.460 2.025 7.470 2.215 ;
        RECT 7.470 2.035 7.480 2.215 ;
        RECT 7.480 2.045 7.490 2.215 ;
        RECT 7.275 1.840 7.285 2.170 ;
        RECT 7.285 1.850 7.295 2.180 ;
        RECT 7.295 1.860 7.305 2.190 ;
        RECT 7.305 1.870 7.315 2.200 ;
        RECT 7.315 1.875 7.321 2.209 ;
        RECT 6.975 1.675 6.985 1.869 ;
        RECT 6.985 1.675 6.995 1.879 ;
        RECT 6.995 1.675 7.005 1.889 ;
        RECT 7.005 1.675 7.015 1.899 ;
        RECT 7.015 1.675 7.025 1.909 ;
        RECT 7.025 1.675 7.035 1.919 ;
        RECT 7.035 1.675 7.045 1.929 ;
        RECT 7.045 1.675 7.055 1.939 ;
        RECT 7.055 1.675 7.065 1.949 ;
        RECT 7.065 1.675 7.075 1.959 ;
        RECT 7.075 1.675 7.085 1.969 ;
        RECT 7.085 1.675 7.095 1.979 ;
        RECT 7.095 1.675 7.105 1.989 ;
        RECT 7.105 1.675 7.115 1.999 ;
        RECT 7.115 1.675 7.125 2.009 ;
        RECT 7.125 1.675 7.135 2.019 ;
        RECT 7.135 1.675 7.145 2.029 ;
        RECT 7.145 1.675 7.155 2.039 ;
        RECT 7.155 1.675 7.165 2.049 ;
        RECT 7.165 1.675 7.175 2.059 ;
        RECT 7.175 1.675 7.185 2.069 ;
        RECT 7.185 1.675 7.195 2.079 ;
        RECT 7.195 1.675 7.205 2.089 ;
        RECT 7.205 1.675 7.215 2.099 ;
        RECT 7.215 1.675 7.225 2.109 ;
        RECT 7.225 1.675 7.235 2.119 ;
        RECT 7.235 1.675 7.245 2.129 ;
        RECT 7.245 1.675 7.255 2.139 ;
        RECT 7.255 1.675 7.265 2.149 ;
        RECT 7.265 1.675 7.275 2.159 ;
        RECT 6.295 0.895 6.685 1.065 ;
        RECT 6.515 0.895 6.685 2.335 ;
        RECT 6.315 2.165 6.855 2.335 ;
        RECT 6.515 1.325 7.690 1.495 ;
        RECT 7.520 1.325 7.690 1.730 ;
        RECT 8.220 1.860 8.390 2.565 ;
        RECT 7.185 2.395 8.390 2.565 ;
        RECT 8.675 1.370 8.845 2.030 ;
        RECT 8.220 1.860 8.845 2.030 ;
        RECT 7.085 2.305 7.095 2.565 ;
        RECT 7.095 2.315 7.105 2.565 ;
        RECT 7.105 2.325 7.115 2.565 ;
        RECT 7.115 2.335 7.125 2.565 ;
        RECT 7.125 2.345 7.135 2.565 ;
        RECT 7.135 2.355 7.145 2.565 ;
        RECT 7.145 2.365 7.155 2.565 ;
        RECT 7.155 2.375 7.165 2.565 ;
        RECT 7.165 2.385 7.175 2.565 ;
        RECT 7.175 2.395 7.185 2.565 ;
        RECT 6.955 2.175 6.965 2.435 ;
        RECT 6.965 2.185 6.975 2.445 ;
        RECT 6.975 2.195 6.985 2.455 ;
        RECT 6.985 2.205 6.995 2.465 ;
        RECT 6.995 2.215 7.005 2.475 ;
        RECT 7.005 2.225 7.015 2.485 ;
        RECT 7.015 2.235 7.025 2.495 ;
        RECT 7.025 2.245 7.035 2.505 ;
        RECT 7.035 2.255 7.045 2.515 ;
        RECT 7.045 2.265 7.055 2.525 ;
        RECT 7.055 2.275 7.065 2.535 ;
        RECT 7.065 2.285 7.075 2.545 ;
        RECT 7.075 2.295 7.085 2.555 ;
        RECT 6.855 2.165 6.865 2.335 ;
        RECT 6.865 2.165 6.875 2.345 ;
        RECT 6.875 2.165 6.885 2.355 ;
        RECT 6.885 2.165 6.895 2.365 ;
        RECT 6.895 2.165 6.905 2.375 ;
        RECT 6.905 2.165 6.915 2.385 ;
        RECT 6.915 2.165 6.925 2.395 ;
        RECT 6.925 2.165 6.935 2.405 ;
        RECT 6.935 2.165 6.945 2.415 ;
        RECT 6.945 2.165 6.955 2.425 ;
  END 
END FFDSHQHDMXHT

MACRO FFDHDLXHT
  CLASS  CORE ;
  FOREIGN FFDHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.610 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.270 1.060 8.510 1.360 ;
        RECT 8.300 1.060 8.510 2.445 ;
        RECT 8.270 1.980 8.510 2.445 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.230 1.060 7.400 1.405 ;
        RECT 7.230 2.000 7.400 2.300 ;
        RECT 7.230 1.225 7.690 1.405 ;
        RECT 7.480 1.225 7.690 2.235 ;
        RECT 7.230 2.000 7.690 2.235 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.600 1.265 1.985 1.765 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.855 ;
        RECT 1.535 -0.300 1.835 0.785 ;
        RECT 3.315 -0.300 3.615 0.645 ;
        RECT 4.410 -0.300 4.710 0.660 ;
        RECT 6.195 -0.300 6.495 0.550 ;
        RECT 7.685 -0.300 7.985 0.745 ;
        RECT 0.000 -0.300 8.610 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 2.745 0.865 3.990 ;
        RECT 1.500 2.745 1.670 3.990 ;
        RECT 3.435 3.160 3.735 3.990 ;
        RECT 4.295 3.160 4.595 3.990 ;
        RECT 6.195 2.830 6.495 3.990 ;
        RECT 7.685 2.860 7.985 3.990 ;
        RECT 0.000 3.390 8.610 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.550 0.920 2.720 2.280 ;
        RECT 2.550 1.675 3.955 1.845 ;
        RECT 3.960 0.840 4.130 1.445 ;
        RECT 3.175 1.275 4.705 1.445 ;
        RECT 4.535 1.275 4.705 2.215 ;
        RECT 3.865 2.045 4.705 2.215 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.195 0.965 2.365 ;
        RECT 0.795 1.125 0.965 2.565 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 2.395 2.020 2.565 ;
        RECT 1.850 2.395 2.020 2.995 ;
        RECT 2.855 2.810 3.155 2.995 ;
        RECT 1.850 2.825 3.155 2.995 ;
        RECT 2.855 2.810 5.175 2.980 ;
        RECT 1.210 1.060 1.400 1.360 ;
        RECT 1.230 1.060 1.400 2.215 ;
        RECT 1.145 2.045 2.370 2.215 ;
        RECT 2.200 0.570 2.370 2.645 ;
        RECT 2.200 2.460 2.575 2.645 ;
        RECT 2.200 0.570 2.995 0.740 ;
        RECT 4.885 1.425 5.055 2.630 ;
        RECT 4.950 0.500 5.120 1.595 ;
        RECT 4.885 1.425 5.120 1.595 ;
        RECT 4.950 0.500 5.285 0.670 ;
        RECT 4.885 2.440 5.755 2.630 ;
        RECT 2.200 2.460 5.755 2.630 ;
        RECT 5.945 1.220 7.050 1.390 ;
        RECT 6.720 0.785 6.890 1.390 ;
        RECT 6.880 1.220 7.050 2.215 ;
        RECT 6.625 2.045 7.050 2.215 ;
        RECT 6.880 1.585 7.275 1.755 ;
        RECT 5.310 0.875 5.480 2.215 ;
        RECT 5.245 2.045 5.545 2.215 ;
        RECT 6.275 1.675 6.445 2.650 ;
        RECT 5.310 1.675 6.700 1.845 ;
        RECT 7.920 1.520 8.090 2.650 ;
        RECT 6.275 2.480 8.090 2.650 ;
        RECT 7.920 1.520 8.110 1.820 ;
  END 
END FFDHDLXHT

MACRO FFDHD2XHT
  CLASS  CORE ;
  FOREIGN FFDHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.250 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.390 0.720 9.560 2.960 ;
        RECT 9.390 1.650 9.740 2.015 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.300 0.720 8.510 2.280 ;
        RECT 8.300 0.720 8.520 1.360 ;
        RECT 8.300 1.980 8.520 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.585 1.265 2.080 1.670 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.745 ;
        RECT 1.680 -0.300 1.980 1.020 ;
        RECT 3.650 -0.300 3.950 1.020 ;
        RECT 4.700 -0.300 5.000 1.055 ;
        RECT 6.475 -0.300 6.645 0.810 ;
        RECT 7.830 -0.300 8.000 1.120 ;
        RECT 8.805 -0.300 9.105 1.055 ;
        RECT 9.845 -0.300 10.145 1.055 ;
        RECT 0.000 -0.300 10.250 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.520 2.015 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.515 2.745 0.815 3.990 ;
        RECT 1.620 2.790 1.790 3.990 ;
        RECT 3.620 3.095 3.920 3.990 ;
        RECT 4.700 3.095 5.000 3.990 ;
        RECT 6.615 2.805 6.785 3.990 ;
        RECT 7.765 2.975 8.065 3.990 ;
        RECT 8.805 2.975 9.105 3.990 ;
        RECT 9.845 2.295 10.145 3.990 ;
        RECT 0.000 3.390 10.250 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.670 0.950 2.970 1.120 ;
        RECT 2.800 0.950 2.970 2.215 ;
        RECT 2.670 2.045 2.970 2.215 ;
        RECT 2.800 1.675 4.190 1.845 ;
        RECT 4.255 0.985 4.425 1.445 ;
        RECT 3.390 1.275 5.120 1.445 ;
        RECT 4.950 1.275 5.120 2.215 ;
        RECT 4.170 2.045 5.120 2.215 ;
        RECT 0.105 1.125 0.880 1.295 ;
        RECT 0.105 2.195 0.880 2.365 ;
        RECT 0.710 1.125 0.880 2.565 ;
        RECT 0.710 1.525 1.000 1.825 ;
        RECT 0.710 2.395 2.140 2.565 ;
        RECT 1.970 2.395 2.140 2.915 ;
        RECT 1.970 2.745 5.685 2.915 ;
        RECT 5.515 2.745 5.685 3.210 ;
        RECT 5.515 3.040 6.200 3.210 ;
        RECT 1.215 1.060 1.385 2.215 ;
        RECT 1.085 2.045 2.490 2.215 ;
        RECT 2.320 0.480 2.490 2.565 ;
        RECT 2.320 1.605 2.555 1.905 ;
        RECT 2.320 0.480 3.210 0.650 ;
        RECT 5.300 0.710 5.470 2.565 ;
        RECT 2.320 2.395 6.135 2.565 ;
        RECT 5.300 0.710 6.240 0.880 ;
        RECT 5.965 2.395 6.135 2.795 ;
        RECT 6.070 0.710 6.240 1.160 ;
        RECT 6.825 0.480 6.995 1.160 ;
        RECT 6.070 0.990 6.995 1.160 ;
        RECT 6.825 0.480 7.650 0.650 ;
        RECT 7.175 1.060 7.345 1.770 ;
        RECT 7.240 1.600 7.410 2.305 ;
        RECT 6.390 1.600 8.120 1.770 ;
        RECT 5.715 1.060 5.885 2.215 ;
        RECT 5.650 2.045 7.060 2.215 ;
        RECT 6.890 2.045 7.060 2.655 ;
        RECT 6.965 2.485 7.265 3.150 ;
        RECT 9.040 1.610 9.210 2.655 ;
        RECT 6.890 2.485 9.210 2.655 ;
  END 
END FFDHD2XHT

MACRO FAHHDLXHT
  CLASS  CORE ;
  FOREIGN FAHHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.250 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.485 0.720 1.820 ;
        RECT 0.510 1.485 0.720 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.135 1.275 4.485 1.840 ;
    END
  END B
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.905 1.060 10.150 1.360 ;
        RECT 9.970 1.060 10.150 2.865 ;
        RECT 9.905 2.100 10.150 2.865 ;
    END
  END S
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.600 1.170 8.100 1.820 ;
    END
  END CI
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.955 ;
        RECT 3.950 -0.300 4.250 0.665 ;
        RECT 7.615 -0.300 7.915 0.550 ;
        RECT 9.365 -0.300 9.535 0.705 ;
        RECT 0.000 -0.300 10.250 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.985 0.955 3.990 ;
        RECT 3.825 2.985 4.125 3.990 ;
        RECT 7.645 3.095 7.945 3.990 ;
        RECT 9.290 2.745 9.590 3.990 ;
        RECT 0.000 3.390 10.250 3.990 ;
    END
  END VDD
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.710 1.060 8.960 2.215 ;
        RECT 8.710 2.045 9.035 2.215 ;
    END
  END CO
  OBS 
      LAYER M1 ;
        RECT 1.270 1.060 1.505 1.360 ;
        RECT 1.335 1.060 1.505 2.455 ;
        RECT 1.205 2.285 1.505 2.455 ;
        RECT 0.090 1.125 0.260 2.805 ;
        RECT 0.090 2.110 0.340 2.805 ;
        RECT 0.090 1.125 0.405 1.305 ;
        RECT 0.090 1.135 1.090 1.305 ;
        RECT 0.920 1.135 1.090 1.850 ;
        RECT 2.310 1.060 2.480 2.805 ;
        RECT 0.090 2.635 2.480 2.805 ;
        RECT 1.235 2.985 3.615 3.155 ;
        RECT 3.180 1.125 3.350 2.455 ;
        RECT 3.180 2.285 3.585 2.455 ;
        RECT 3.180 1.125 3.615 1.295 ;
        RECT 3.530 1.625 3.935 1.795 ;
        RECT 3.765 1.625 3.935 2.250 ;
        RECT 4.820 0.855 4.990 2.250 ;
        RECT 3.765 2.045 4.990 2.250 ;
        RECT 3.765 2.055 5.310 2.250 ;
        RECT 1.790 0.710 1.960 2.455 ;
        RECT 1.725 2.280 2.025 2.455 ;
        RECT 1.790 0.710 3.635 0.880 ;
        RECT 4.470 0.500 4.640 1.020 ;
        RECT 3.850 0.850 4.640 1.020 ;
        RECT 4.470 0.500 5.395 0.670 ;
        RECT 3.775 0.785 3.785 1.019 ;
        RECT 3.785 0.795 3.795 1.019 ;
        RECT 3.795 0.805 3.805 1.019 ;
        RECT 3.805 0.815 3.815 1.019 ;
        RECT 3.815 0.825 3.825 1.019 ;
        RECT 3.825 0.835 3.835 1.019 ;
        RECT 3.835 0.845 3.845 1.019 ;
        RECT 3.845 0.850 3.851 1.020 ;
        RECT 3.710 0.720 3.720 0.954 ;
        RECT 3.720 0.730 3.730 0.964 ;
        RECT 3.730 0.740 3.740 0.974 ;
        RECT 3.740 0.750 3.750 0.984 ;
        RECT 3.750 0.760 3.760 0.994 ;
        RECT 3.760 0.770 3.770 1.004 ;
        RECT 3.770 0.775 3.776 1.015 ;
        RECT 3.635 0.710 3.645 0.880 ;
        RECT 3.645 0.710 3.655 0.890 ;
        RECT 3.655 0.710 3.665 0.900 ;
        RECT 3.665 0.710 3.675 0.910 ;
        RECT 3.675 0.710 3.685 0.920 ;
        RECT 3.685 0.710 3.695 0.930 ;
        RECT 3.695 0.710 3.705 0.940 ;
        RECT 3.705 0.710 3.711 0.950 ;
        RECT 2.830 1.060 3.000 2.805 ;
        RECT 3.890 2.480 4.060 2.805 ;
        RECT 2.830 2.635 4.060 2.805 ;
        RECT 3.890 2.480 5.490 2.650 ;
        RECT 5.935 2.675 6.105 3.000 ;
        RECT 4.640 2.830 6.105 3.000 ;
        RECT 7.185 1.060 7.355 2.215 ;
        RECT 7.120 2.045 7.420 2.215 ;
        RECT 8.280 1.060 8.450 2.215 ;
        RECT 8.200 2.045 8.500 2.215 ;
        RECT 6.115 2.165 6.455 2.335 ;
        RECT 6.115 0.920 6.285 2.335 ;
        RECT 6.050 0.920 6.350 1.090 ;
        RECT 6.285 2.165 6.455 2.915 ;
        RECT 6.285 2.745 8.525 2.915 ;
        RECT 5.420 0.920 5.765 1.090 ;
        RECT 5.595 0.570 5.765 2.315 ;
        RECT 5.595 0.570 7.295 0.740 ;
        RECT 7.625 0.820 7.925 0.990 ;
        RECT 8.110 0.710 9.035 0.880 ;
        RECT 9.140 0.750 9.150 1.820 ;
        RECT 9.150 0.760 9.160 1.820 ;
        RECT 9.160 0.770 9.170 1.820 ;
        RECT 9.170 0.780 9.180 1.820 ;
        RECT 9.180 0.790 9.190 1.820 ;
        RECT 9.190 0.800 9.200 1.820 ;
        RECT 9.200 0.810 9.210 1.820 ;
        RECT 9.210 0.820 9.220 1.820 ;
        RECT 9.220 0.830 9.230 1.820 ;
        RECT 9.230 0.840 9.240 1.820 ;
        RECT 9.240 0.850 9.250 1.820 ;
        RECT 9.250 0.860 9.260 1.820 ;
        RECT 9.260 0.870 9.270 1.820 ;
        RECT 9.270 0.880 9.280 1.820 ;
        RECT 9.280 0.890 9.290 1.820 ;
        RECT 9.290 0.900 9.300 1.820 ;
        RECT 9.300 0.910 9.310 1.820 ;
        RECT 9.110 0.720 9.120 0.954 ;
        RECT 9.120 0.730 9.130 0.964 ;
        RECT 9.130 0.740 9.140 0.974 ;
        RECT 9.035 0.710 9.045 0.880 ;
        RECT 9.045 0.710 9.055 0.890 ;
        RECT 9.055 0.710 9.065 0.900 ;
        RECT 9.065 0.710 9.075 0.910 ;
        RECT 9.075 0.710 9.085 0.920 ;
        RECT 9.085 0.710 9.095 0.930 ;
        RECT 9.095 0.710 9.105 0.940 ;
        RECT 9.105 0.710 9.111 0.950 ;
        RECT 8.035 0.710 8.045 0.944 ;
        RECT 8.045 0.710 8.055 0.934 ;
        RECT 8.055 0.710 8.065 0.924 ;
        RECT 8.065 0.710 8.075 0.914 ;
        RECT 8.075 0.710 8.085 0.904 ;
        RECT 8.085 0.710 8.095 0.894 ;
        RECT 8.095 0.710 8.105 0.884 ;
        RECT 8.105 0.710 8.111 0.880 ;
        RECT 8.000 0.745 8.010 0.979 ;
        RECT 8.010 0.735 8.020 0.969 ;
        RECT 8.020 0.725 8.030 0.959 ;
        RECT 8.030 0.715 8.036 0.955 ;
        RECT 7.925 0.820 7.935 0.990 ;
        RECT 7.935 0.810 7.945 0.990 ;
        RECT 7.945 0.800 7.955 0.990 ;
        RECT 7.955 0.790 7.965 0.990 ;
        RECT 7.965 0.780 7.975 0.990 ;
        RECT 7.975 0.770 7.985 0.990 ;
        RECT 7.985 0.760 7.995 0.990 ;
        RECT 7.995 0.750 8.001 0.990 ;
        RECT 7.545 0.750 7.555 0.990 ;
        RECT 7.555 0.760 7.565 0.990 ;
        RECT 7.565 0.770 7.575 0.990 ;
        RECT 7.575 0.780 7.585 0.990 ;
        RECT 7.585 0.790 7.595 0.990 ;
        RECT 7.595 0.800 7.605 0.990 ;
        RECT 7.605 0.810 7.615 0.990 ;
        RECT 7.615 0.820 7.625 0.990 ;
        RECT 7.375 0.580 7.385 0.820 ;
        RECT 7.385 0.590 7.395 0.830 ;
        RECT 7.395 0.600 7.405 0.840 ;
        RECT 7.405 0.610 7.415 0.850 ;
        RECT 7.415 0.620 7.425 0.860 ;
        RECT 7.425 0.630 7.435 0.870 ;
        RECT 7.435 0.640 7.445 0.880 ;
        RECT 7.445 0.650 7.455 0.890 ;
        RECT 7.455 0.660 7.465 0.900 ;
        RECT 7.465 0.670 7.475 0.910 ;
        RECT 7.475 0.680 7.485 0.920 ;
        RECT 7.485 0.690 7.495 0.930 ;
        RECT 7.495 0.700 7.505 0.940 ;
        RECT 7.505 0.710 7.515 0.950 ;
        RECT 7.515 0.720 7.525 0.960 ;
        RECT 7.525 0.730 7.535 0.970 ;
        RECT 7.535 0.740 7.545 0.980 ;
        RECT 7.295 0.570 7.305 0.740 ;
        RECT 7.305 0.570 7.315 0.750 ;
        RECT 7.315 0.570 7.325 0.760 ;
        RECT 7.325 0.570 7.335 0.770 ;
        RECT 7.335 0.570 7.345 0.780 ;
        RECT 7.345 0.570 7.355 0.790 ;
        RECT 7.355 0.570 7.365 0.800 ;
        RECT 7.365 0.570 7.375 0.810 ;
        RECT 6.635 0.920 6.805 2.565 ;
        RECT 6.570 0.920 6.870 1.090 ;
        RECT 9.545 1.520 9.715 2.565 ;
        RECT 6.635 2.395 9.715 2.565 ;
        RECT 9.545 1.520 9.790 1.820 ;
  END 
END FAHHDLXHT

MACRO FAHDLXHT
  CLASS  CORE ;
  FOREIGN FAHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.590 1.125 4.010 1.795 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 1.550 0.925 1.970 ;
    END
  END B
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.275 1.060 10.445 2.830 ;
        RECT 10.275 2.500 10.560 2.830 ;
    END
  END S
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.885 2.125 7.340 2.560 ;
    END
  END CI
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.075 ;
        RECT 1.175 -0.300 1.475 0.920 ;
        RECT 3.570 -0.300 3.870 0.460 ;
        RECT 7.375 -0.300 7.675 0.435 ;
        RECT 9.690 -0.300 9.990 1.295 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.465 0.405 3.990 ;
        RECT 1.135 3.070 1.435 3.990 ;
        RECT 3.585 3.025 3.885 3.990 ;
        RECT 6.930 3.090 7.230 3.990 ;
        RECT 9.660 2.810 9.960 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.120 0.860 9.330 2.280 ;
        RECT 9.120 0.860 9.405 1.360 ;
    END
  END CO
  OBS 
      LAYER M1 ;
        RECT 1.795 1.035 1.965 2.540 ;
        RECT 1.750 2.135 1.965 2.540 ;
        RECT 1.750 2.370 2.490 2.540 ;
        RECT 2.320 2.370 2.490 2.860 ;
        RECT 2.320 2.690 2.790 2.860 ;
        RECT 3.085 0.990 3.255 2.145 ;
        RECT 4.200 0.990 4.370 1.530 ;
        RECT 4.265 1.360 4.435 2.145 ;
        RECT 3.035 1.975 4.435 2.145 ;
        RECT 4.200 1.360 5.060 1.530 ;
        RECT 4.890 1.360 5.060 1.660 ;
        RECT 0.625 1.100 1.570 1.270 ;
        RECT 0.625 2.290 1.570 2.460 ;
        RECT 1.400 1.100 1.570 2.890 ;
        RECT 1.400 1.515 1.615 1.815 ;
        RECT 1.400 2.720 2.140 2.890 ;
        RECT 1.970 2.720 2.140 3.210 ;
        RECT 1.970 3.040 2.875 3.210 ;
        RECT 3.140 2.675 4.360 2.845 ;
        RECT 4.190 2.675 4.360 3.085 ;
        RECT 5.270 2.190 5.440 3.085 ;
        RECT 4.190 2.915 5.440 3.085 ;
        RECT 5.270 2.190 5.545 2.360 ;
        RECT 5.590 1.245 5.760 1.415 ;
        RECT 5.760 1.245 5.770 2.209 ;
        RECT 5.770 1.245 5.780 2.199 ;
        RECT 5.780 1.245 5.790 2.189 ;
        RECT 5.790 1.245 5.800 2.179 ;
        RECT 5.800 1.245 5.810 2.169 ;
        RECT 5.810 1.245 5.820 2.159 ;
        RECT 5.820 1.245 5.830 2.149 ;
        RECT 5.830 1.245 5.840 2.139 ;
        RECT 5.840 1.245 5.850 2.129 ;
        RECT 5.850 1.245 5.860 2.119 ;
        RECT 5.860 1.245 5.870 2.109 ;
        RECT 5.870 1.245 5.880 2.099 ;
        RECT 5.880 1.245 5.890 2.089 ;
        RECT 5.890 1.245 5.900 2.079 ;
        RECT 5.900 1.245 5.910 2.069 ;
        RECT 5.910 1.245 5.920 2.059 ;
        RECT 5.920 1.245 5.930 2.049 ;
        RECT 5.620 2.115 5.630 2.349 ;
        RECT 5.630 2.105 5.640 2.339 ;
        RECT 5.640 2.095 5.650 2.329 ;
        RECT 5.650 2.085 5.660 2.319 ;
        RECT 5.660 2.075 5.670 2.309 ;
        RECT 5.670 2.065 5.680 2.299 ;
        RECT 5.680 2.055 5.690 2.289 ;
        RECT 5.690 2.045 5.700 2.279 ;
        RECT 5.700 2.035 5.710 2.269 ;
        RECT 5.710 2.025 5.720 2.259 ;
        RECT 5.720 2.015 5.730 2.249 ;
        RECT 5.730 2.005 5.740 2.239 ;
        RECT 5.740 1.995 5.750 2.229 ;
        RECT 5.750 1.985 5.760 2.219 ;
        RECT 5.545 2.190 5.555 2.360 ;
        RECT 5.555 2.180 5.565 2.360 ;
        RECT 5.565 2.170 5.575 2.360 ;
        RECT 5.575 2.160 5.585 2.360 ;
        RECT 5.585 2.150 5.595 2.360 ;
        RECT 5.595 2.140 5.605 2.360 ;
        RECT 5.605 2.130 5.615 2.360 ;
        RECT 5.615 2.120 5.621 2.360 ;
        RECT 2.970 2.675 2.980 3.179 ;
        RECT 2.980 2.675 2.990 3.169 ;
        RECT 2.990 2.675 3.000 3.159 ;
        RECT 3.000 2.675 3.010 3.149 ;
        RECT 3.010 2.675 3.020 3.139 ;
        RECT 3.020 2.675 3.030 3.129 ;
        RECT 3.030 2.675 3.040 3.119 ;
        RECT 3.040 2.675 3.050 3.109 ;
        RECT 3.050 2.675 3.060 3.099 ;
        RECT 3.060 2.675 3.070 3.089 ;
        RECT 3.070 2.675 3.080 3.079 ;
        RECT 3.080 2.675 3.090 3.069 ;
        RECT 3.090 2.675 3.100 3.059 ;
        RECT 3.100 2.675 3.110 3.049 ;
        RECT 3.110 2.675 3.120 3.039 ;
        RECT 3.120 2.675 3.130 3.029 ;
        RECT 3.130 2.675 3.140 3.019 ;
        RECT 2.950 2.965 2.960 3.199 ;
        RECT 2.960 2.955 2.970 3.189 ;
        RECT 2.875 3.040 2.885 3.210 ;
        RECT 2.885 3.030 2.895 3.210 ;
        RECT 2.895 3.020 2.905 3.210 ;
        RECT 2.905 3.010 2.915 3.210 ;
        RECT 2.915 3.000 2.925 3.210 ;
        RECT 2.925 2.990 2.935 3.210 ;
        RECT 2.935 2.980 2.945 3.210 ;
        RECT 2.945 2.970 2.951 3.210 ;
        RECT 6.705 1.245 6.800 1.935 ;
        RECT 6.705 1.245 6.930 1.415 ;
        RECT 6.705 1.765 7.620 1.935 ;
        RECT 6.630 1.245 6.640 2.395 ;
        RECT 6.640 1.245 6.650 2.385 ;
        RECT 6.650 1.245 6.660 2.375 ;
        RECT 6.660 1.245 6.670 2.365 ;
        RECT 6.670 1.245 6.680 2.355 ;
        RECT 6.680 1.245 6.690 2.345 ;
        RECT 6.690 1.245 6.700 2.335 ;
        RECT 6.700 1.245 6.706 2.329 ;
        RECT 6.535 1.765 6.545 2.489 ;
        RECT 6.545 1.765 6.555 2.479 ;
        RECT 6.555 1.765 6.565 2.469 ;
        RECT 6.565 1.765 6.575 2.459 ;
        RECT 6.575 1.765 6.585 2.449 ;
        RECT 6.585 1.765 6.595 2.439 ;
        RECT 6.595 1.765 6.605 2.429 ;
        RECT 6.605 1.765 6.615 2.419 ;
        RECT 6.615 1.765 6.625 2.409 ;
        RECT 6.625 1.765 6.631 2.405 ;
        RECT 6.480 2.310 6.490 2.544 ;
        RECT 6.490 2.300 6.500 2.534 ;
        RECT 6.500 2.290 6.510 2.524 ;
        RECT 6.510 2.280 6.520 2.514 ;
        RECT 6.520 2.270 6.530 2.504 ;
        RECT 6.530 2.260 6.536 2.500 ;
        RECT 6.310 2.480 6.320 2.780 ;
        RECT 6.320 2.470 6.330 2.780 ;
        RECT 6.330 2.460 6.340 2.780 ;
        RECT 6.340 2.450 6.350 2.780 ;
        RECT 6.350 2.440 6.360 2.780 ;
        RECT 6.360 2.430 6.370 2.780 ;
        RECT 6.370 2.420 6.380 2.780 ;
        RECT 6.380 2.410 6.390 2.780 ;
        RECT 6.390 2.400 6.400 2.780 ;
        RECT 6.400 2.390 6.410 2.780 ;
        RECT 6.410 2.380 6.420 2.780 ;
        RECT 6.420 2.370 6.430 2.780 ;
        RECT 6.430 2.360 6.440 2.780 ;
        RECT 6.440 2.350 6.450 2.780 ;
        RECT 6.450 2.340 6.460 2.780 ;
        RECT 6.460 2.330 6.470 2.780 ;
        RECT 6.470 2.320 6.480 2.780 ;
        RECT 2.560 1.470 2.855 1.640 ;
        RECT 2.560 0.990 2.730 1.640 ;
        RECT 2.685 1.470 2.855 2.495 ;
        RECT 4.750 1.840 4.920 2.495 ;
        RECT 2.685 2.325 4.920 2.495 ;
        RECT 5.240 0.875 5.410 2.010 ;
        RECT 4.750 1.840 5.410 2.010 ;
        RECT 5.240 1.600 5.580 1.900 ;
        RECT 5.240 0.875 6.985 1.045 ;
        RECT 7.585 2.115 7.755 2.500 ;
        RECT 7.255 1.070 7.970 1.240 ;
        RECT 7.800 1.070 7.970 2.285 ;
        RECT 7.585 2.115 7.970 2.285 ;
        RECT 7.180 1.005 7.190 1.239 ;
        RECT 7.190 1.015 7.200 1.239 ;
        RECT 7.200 1.025 7.210 1.239 ;
        RECT 7.210 1.035 7.220 1.239 ;
        RECT 7.220 1.045 7.230 1.239 ;
        RECT 7.230 1.055 7.240 1.239 ;
        RECT 7.240 1.065 7.250 1.239 ;
        RECT 7.250 1.070 7.256 1.240 ;
        RECT 7.060 0.885 7.070 1.119 ;
        RECT 7.070 0.895 7.080 1.129 ;
        RECT 7.080 0.905 7.090 1.139 ;
        RECT 7.090 0.915 7.100 1.149 ;
        RECT 7.100 0.925 7.110 1.159 ;
        RECT 7.110 0.935 7.120 1.169 ;
        RECT 7.120 0.945 7.130 1.179 ;
        RECT 7.130 0.955 7.140 1.189 ;
        RECT 7.140 0.965 7.150 1.199 ;
        RECT 7.150 0.975 7.160 1.209 ;
        RECT 7.160 0.985 7.170 1.219 ;
        RECT 7.170 0.995 7.180 1.229 ;
        RECT 6.985 0.875 6.995 1.045 ;
        RECT 6.995 0.875 7.005 1.055 ;
        RECT 7.005 0.875 7.015 1.065 ;
        RECT 7.015 0.875 7.025 1.075 ;
        RECT 7.025 0.875 7.035 1.085 ;
        RECT 7.035 0.875 7.045 1.095 ;
        RECT 7.045 0.875 7.055 1.105 ;
        RECT 7.055 0.875 7.061 1.115 ;
        RECT 2.205 0.640 2.375 2.190 ;
        RECT 2.205 2.020 2.505 2.190 ;
        RECT 2.205 0.640 4.890 0.810 ;
        RECT 4.720 0.525 4.890 1.170 ;
        RECT 4.720 0.525 7.135 0.695 ;
        RECT 7.345 0.660 8.895 0.830 ;
        RECT 8.725 0.660 8.895 2.435 ;
        RECT 8.560 2.265 8.895 2.435 ;
        RECT 7.270 0.595 7.280 0.829 ;
        RECT 7.280 0.605 7.290 0.829 ;
        RECT 7.290 0.615 7.300 0.829 ;
        RECT 7.300 0.625 7.310 0.829 ;
        RECT 7.310 0.635 7.320 0.829 ;
        RECT 7.320 0.645 7.330 0.829 ;
        RECT 7.330 0.655 7.340 0.829 ;
        RECT 7.340 0.660 7.346 0.830 ;
        RECT 7.210 0.535 7.220 0.769 ;
        RECT 7.220 0.545 7.230 0.779 ;
        RECT 7.230 0.555 7.240 0.789 ;
        RECT 7.240 0.565 7.250 0.799 ;
        RECT 7.250 0.575 7.260 0.809 ;
        RECT 7.260 0.585 7.270 0.819 ;
        RECT 7.135 0.525 7.145 0.695 ;
        RECT 7.145 0.525 7.155 0.705 ;
        RECT 7.155 0.525 7.165 0.715 ;
        RECT 7.165 0.525 7.175 0.725 ;
        RECT 7.175 0.525 7.185 0.735 ;
        RECT 7.185 0.525 7.195 0.745 ;
        RECT 7.195 0.525 7.205 0.755 ;
        RECT 7.205 0.525 7.211 0.765 ;
        RECT 5.725 2.545 5.960 2.715 ;
        RECT 6.110 1.245 6.175 1.415 ;
        RECT 6.345 1.245 6.410 1.415 ;
        RECT 6.130 2.960 6.555 3.130 ;
        RECT 6.850 2.740 7.860 2.910 ;
        RECT 7.690 2.740 7.860 3.135 ;
        RECT 7.690 2.965 9.480 3.135 ;
        RECT 6.775 2.740 6.785 2.974 ;
        RECT 6.785 2.740 6.795 2.964 ;
        RECT 6.795 2.740 6.805 2.954 ;
        RECT 6.805 2.740 6.815 2.944 ;
        RECT 6.815 2.740 6.825 2.934 ;
        RECT 6.825 2.740 6.835 2.924 ;
        RECT 6.835 2.740 6.845 2.914 ;
        RECT 6.845 2.740 6.851 2.910 ;
        RECT 6.630 2.885 6.640 3.119 ;
        RECT 6.640 2.875 6.650 3.109 ;
        RECT 6.650 2.865 6.660 3.099 ;
        RECT 6.660 2.855 6.670 3.089 ;
        RECT 6.670 2.845 6.680 3.079 ;
        RECT 6.680 2.835 6.690 3.069 ;
        RECT 6.690 2.825 6.700 3.059 ;
        RECT 6.700 2.815 6.710 3.049 ;
        RECT 6.710 2.805 6.720 3.039 ;
        RECT 6.720 2.795 6.730 3.029 ;
        RECT 6.730 2.785 6.740 3.019 ;
        RECT 6.740 2.775 6.750 3.009 ;
        RECT 6.750 2.765 6.760 2.999 ;
        RECT 6.760 2.755 6.770 2.989 ;
        RECT 6.770 2.745 6.776 2.985 ;
        RECT 6.555 2.960 6.565 3.130 ;
        RECT 6.565 2.950 6.575 3.130 ;
        RECT 6.575 2.940 6.585 3.130 ;
        RECT 6.585 2.930 6.595 3.130 ;
        RECT 6.595 2.920 6.605 3.130 ;
        RECT 6.605 2.910 6.615 3.130 ;
        RECT 6.615 2.900 6.625 3.130 ;
        RECT 6.625 2.890 6.631 3.130 ;
        RECT 6.175 1.245 6.185 2.325 ;
        RECT 6.185 1.245 6.195 2.315 ;
        RECT 6.195 1.245 6.205 2.305 ;
        RECT 6.205 1.245 6.215 2.295 ;
        RECT 6.215 1.245 6.225 2.285 ;
        RECT 6.225 1.245 6.235 2.275 ;
        RECT 6.235 1.245 6.245 2.265 ;
        RECT 6.245 1.245 6.255 2.255 ;
        RECT 6.255 1.245 6.265 2.245 ;
        RECT 6.265 1.245 6.275 2.235 ;
        RECT 6.275 1.245 6.285 2.225 ;
        RECT 6.285 1.245 6.295 2.215 ;
        RECT 6.295 1.245 6.305 2.205 ;
        RECT 6.305 1.245 6.315 2.195 ;
        RECT 6.315 1.245 6.325 2.185 ;
        RECT 6.325 1.245 6.335 2.175 ;
        RECT 6.335 1.245 6.345 2.165 ;
        RECT 6.130 2.135 6.140 2.369 ;
        RECT 6.140 2.125 6.150 2.359 ;
        RECT 6.150 2.115 6.160 2.349 ;
        RECT 6.160 2.105 6.170 2.339 ;
        RECT 6.170 2.095 6.176 2.335 ;
        RECT 5.960 2.305 5.970 3.129 ;
        RECT 5.970 2.295 5.980 3.129 ;
        RECT 5.980 2.285 5.990 3.129 ;
        RECT 5.990 2.275 6.000 3.129 ;
        RECT 6.000 2.265 6.010 3.129 ;
        RECT 6.010 2.255 6.020 3.129 ;
        RECT 6.020 2.245 6.030 3.129 ;
        RECT 6.030 2.235 6.040 3.129 ;
        RECT 6.040 2.225 6.050 3.129 ;
        RECT 6.050 2.215 6.060 3.129 ;
        RECT 6.060 2.205 6.070 3.129 ;
        RECT 6.070 2.195 6.080 3.129 ;
        RECT 6.080 2.185 6.090 3.129 ;
        RECT 6.090 2.175 6.100 3.129 ;
        RECT 6.100 2.165 6.110 3.129 ;
        RECT 6.110 2.155 6.120 3.129 ;
        RECT 6.120 2.145 6.130 3.129 ;
        RECT 8.205 1.010 8.375 2.785 ;
        RECT 8.040 2.465 8.375 2.785 ;
        RECT 9.135 2.460 9.305 2.785 ;
        RECT 8.040 2.615 9.305 2.785 ;
        RECT 9.135 2.460 10.095 2.630 ;
        RECT 9.925 1.545 10.095 2.630 ;
  END 
END FAHDLXHT

MACRO FAHD2XHT
  CLASS  CORE ;
  FOREIGN FAHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.300 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.790 1.225 4.235 1.885 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.205 1.550 0.925 1.955 ;
    END
  END B
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.430 1.170 11.810 1.340 ;
        RECT 11.580 0.700 11.600 2.980 ;
        RECT 11.430 0.700 11.600 1.340 ;
        RECT 11.580 1.170 11.620 2.980 ;
        RECT 11.410 2.000 11.620 2.980 ;
        RECT 11.580 1.170 11.810 2.170 ;
        RECT 11.410 2.000 11.810 2.170 ;
    END
  END S
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.275 1.940 7.575 2.620 ;
        RECT 7.275 2.135 7.835 2.620 ;
    END
  END CI
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.205 ;
        RECT 1.145 -0.300 1.445 1.005 ;
        RECT 3.935 -0.300 4.235 0.595 ;
        RECT 7.685 -0.300 7.985 0.435 ;
        RECT 9.805 -0.300 10.105 1.065 ;
        RECT 10.845 -0.300 11.145 1.065 ;
        RECT 11.885 -0.300 12.185 0.715 ;
        RECT 0.000 -0.300 12.300 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 1.145 2.945 1.445 3.990 ;
        RECT 3.970 3.255 4.270 3.990 ;
        RECT 7.330 3.205 7.630 3.990 ;
        RECT 9.805 2.975 10.105 3.990 ;
        RECT 10.845 2.975 11.145 3.990 ;
        RECT 11.885 2.635 12.185 3.990 ;
        RECT 0.000 3.390 12.300 3.990 ;
    END
  END VDD
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.350 0.720 10.580 2.280 ;
    END
  END CO
  OBS 
      LAYER M1 ;
        RECT 1.730 0.480 1.900 2.430 ;
        RECT 1.730 0.480 2.230 0.650 ;
        RECT 2.780 1.655 2.950 1.955 ;
        RECT 2.780 1.785 3.545 1.955 ;
        RECT 3.375 1.060 3.545 2.375 ;
        RECT 3.375 1.060 3.610 1.360 ;
        RECT 4.580 1.060 4.750 1.530 ;
        RECT 4.715 1.360 4.885 2.375 ;
        RECT 3.375 2.205 4.885 2.375 ;
        RECT 4.580 1.360 5.460 1.530 ;
        RECT 5.290 1.360 5.460 1.660 ;
        RECT 0.690 0.720 0.860 1.365 ;
        RECT 0.690 2.135 0.860 3.115 ;
        RECT 0.690 1.185 1.380 1.365 ;
        RECT 0.690 2.135 1.380 2.305 ;
        RECT 3.595 2.905 3.765 3.150 ;
        RECT 1.795 2.980 3.765 3.150 ;
        RECT 4.865 2.905 5.165 3.210 ;
        RECT 3.595 2.905 5.900 3.075 ;
        RECT 5.730 2.190 5.900 3.075 ;
        RECT 5.730 2.190 6.115 2.360 ;
        RECT 5.990 1.355 6.225 1.525 ;
        RECT 6.225 1.355 6.235 2.315 ;
        RECT 6.235 1.355 6.245 2.305 ;
        RECT 6.245 1.355 6.255 2.295 ;
        RECT 6.255 1.355 6.265 2.285 ;
        RECT 6.265 1.355 6.275 2.275 ;
        RECT 6.275 1.355 6.285 2.265 ;
        RECT 6.285 1.355 6.295 2.255 ;
        RECT 6.295 1.355 6.305 2.245 ;
        RECT 6.305 1.355 6.315 2.235 ;
        RECT 6.315 1.355 6.325 2.225 ;
        RECT 6.325 1.355 6.335 2.215 ;
        RECT 6.335 1.355 6.345 2.205 ;
        RECT 6.345 1.355 6.355 2.195 ;
        RECT 6.355 1.355 6.365 2.185 ;
        RECT 6.365 1.355 6.375 2.175 ;
        RECT 6.375 1.355 6.385 2.165 ;
        RECT 6.385 1.355 6.395 2.155 ;
        RECT 6.190 2.115 6.200 2.349 ;
        RECT 6.200 2.105 6.210 2.339 ;
        RECT 6.210 2.095 6.220 2.329 ;
        RECT 6.220 2.085 6.226 2.325 ;
        RECT 6.115 2.190 6.125 2.360 ;
        RECT 6.125 2.180 6.135 2.360 ;
        RECT 6.135 2.170 6.145 2.360 ;
        RECT 6.145 2.160 6.155 2.360 ;
        RECT 6.155 2.150 6.165 2.360 ;
        RECT 6.165 2.140 6.175 2.360 ;
        RECT 6.175 2.130 6.185 2.360 ;
        RECT 6.185 2.120 6.191 2.360 ;
        RECT 1.625 2.610 1.635 3.150 ;
        RECT 1.635 2.620 1.645 3.150 ;
        RECT 1.645 2.630 1.655 3.150 ;
        RECT 1.655 2.640 1.665 3.150 ;
        RECT 1.665 2.650 1.675 3.150 ;
        RECT 1.675 2.660 1.685 3.150 ;
        RECT 1.685 2.670 1.695 3.150 ;
        RECT 1.695 2.680 1.705 3.150 ;
        RECT 1.705 2.690 1.715 3.150 ;
        RECT 1.715 2.700 1.725 3.150 ;
        RECT 1.725 2.710 1.735 3.150 ;
        RECT 1.735 2.720 1.745 3.150 ;
        RECT 1.745 2.730 1.755 3.150 ;
        RECT 1.755 2.740 1.765 3.150 ;
        RECT 1.765 2.750 1.775 3.150 ;
        RECT 1.775 2.760 1.785 3.150 ;
        RECT 1.785 2.770 1.795 3.150 ;
        RECT 1.550 2.535 1.560 2.769 ;
        RECT 1.560 2.545 1.570 2.779 ;
        RECT 1.570 2.555 1.580 2.789 ;
        RECT 1.580 2.565 1.590 2.799 ;
        RECT 1.590 2.575 1.600 2.809 ;
        RECT 1.600 2.585 1.610 2.819 ;
        RECT 1.610 2.595 1.620 2.829 ;
        RECT 1.620 2.600 1.626 2.840 ;
        RECT 1.380 1.185 1.390 2.599 ;
        RECT 1.390 1.185 1.400 2.609 ;
        RECT 1.400 1.185 1.410 2.619 ;
        RECT 1.410 1.185 1.420 2.629 ;
        RECT 1.420 1.185 1.430 2.639 ;
        RECT 1.430 1.185 1.440 2.649 ;
        RECT 1.440 1.185 1.450 2.659 ;
        RECT 1.450 1.185 1.460 2.669 ;
        RECT 1.460 1.185 1.470 2.679 ;
        RECT 1.470 1.185 1.480 2.689 ;
        RECT 1.480 1.185 1.490 2.699 ;
        RECT 1.490 1.185 1.500 2.709 ;
        RECT 1.500 1.185 1.510 2.719 ;
        RECT 1.510 1.185 1.520 2.729 ;
        RECT 1.520 1.185 1.530 2.739 ;
        RECT 1.530 1.185 1.540 2.749 ;
        RECT 1.540 1.185 1.550 2.759 ;
        RECT 6.925 1.590 6.940 2.840 ;
        RECT 7.095 1.290 7.265 1.760 ;
        RECT 7.095 1.590 8.055 1.760 ;
        RECT 7.755 1.590 8.055 1.935 ;
        RECT 6.940 1.590 6.950 2.604 ;
        RECT 6.950 1.590 6.960 2.594 ;
        RECT 6.960 1.590 6.970 2.584 ;
        RECT 6.970 1.590 6.980 2.574 ;
        RECT 6.980 1.590 6.990 2.564 ;
        RECT 6.990 1.590 7.000 2.554 ;
        RECT 7.000 1.590 7.010 2.544 ;
        RECT 7.010 1.590 7.020 2.534 ;
        RECT 7.020 1.590 7.030 2.524 ;
        RECT 7.030 1.590 7.040 2.514 ;
        RECT 7.040 1.590 7.050 2.504 ;
        RECT 7.050 1.590 7.060 2.494 ;
        RECT 7.060 1.590 7.070 2.484 ;
        RECT 7.070 1.590 7.080 2.474 ;
        RECT 7.080 1.590 7.090 2.464 ;
        RECT 7.090 1.590 7.096 2.460 ;
        RECT 6.770 2.540 6.780 2.840 ;
        RECT 6.780 2.530 6.790 2.840 ;
        RECT 6.790 2.520 6.800 2.840 ;
        RECT 6.800 2.510 6.810 2.840 ;
        RECT 6.810 2.500 6.820 2.840 ;
        RECT 6.820 2.490 6.830 2.840 ;
        RECT 6.830 2.480 6.840 2.840 ;
        RECT 6.840 2.470 6.850 2.840 ;
        RECT 6.850 2.460 6.860 2.840 ;
        RECT 6.860 2.450 6.870 2.840 ;
        RECT 6.870 2.440 6.880 2.840 ;
        RECT 6.880 2.430 6.890 2.840 ;
        RECT 6.890 2.420 6.900 2.840 ;
        RECT 6.900 2.410 6.910 2.840 ;
        RECT 6.910 2.400 6.920 2.840 ;
        RECT 6.920 2.390 6.926 2.840 ;
        RECT 2.430 1.275 2.600 2.305 ;
        RECT 2.430 2.135 3.190 2.305 ;
        RECT 2.920 1.060 3.090 1.445 ;
        RECT 2.430 1.275 3.090 1.445 ;
        RECT 3.020 2.135 3.190 2.725 ;
        RECT 5.190 1.840 5.360 2.725 ;
        RECT 3.020 2.555 5.360 2.725 ;
        RECT 5.640 0.875 5.810 2.010 ;
        RECT 5.640 1.710 6.040 2.010 ;
        RECT 5.190 1.840 6.040 2.010 ;
        RECT 5.640 0.875 7.290 1.045 ;
        RECT 8.070 2.115 8.240 2.500 ;
        RECT 7.500 1.010 8.430 1.180 ;
        RECT 8.260 1.010 8.430 2.285 ;
        RECT 8.070 2.115 8.430 2.285 ;
        RECT 7.425 0.945 7.435 1.179 ;
        RECT 7.435 0.955 7.445 1.179 ;
        RECT 7.445 0.965 7.455 1.179 ;
        RECT 7.455 0.975 7.465 1.179 ;
        RECT 7.465 0.985 7.475 1.179 ;
        RECT 7.475 0.995 7.485 1.179 ;
        RECT 7.485 1.005 7.495 1.179 ;
        RECT 7.495 1.010 7.501 1.180 ;
        RECT 7.365 0.885 7.375 1.119 ;
        RECT 7.375 0.895 7.385 1.129 ;
        RECT 7.385 0.905 7.395 1.139 ;
        RECT 7.395 0.915 7.405 1.149 ;
        RECT 7.405 0.925 7.415 1.159 ;
        RECT 7.415 0.935 7.425 1.169 ;
        RECT 7.290 0.875 7.300 1.045 ;
        RECT 7.300 0.875 7.310 1.055 ;
        RECT 7.310 0.875 7.320 1.065 ;
        RECT 7.320 0.875 7.330 1.075 ;
        RECT 7.330 0.875 7.340 1.085 ;
        RECT 7.340 0.875 7.350 1.095 ;
        RECT 7.350 0.875 7.360 1.105 ;
        RECT 7.360 0.875 7.366 1.115 ;
        RECT 2.080 0.925 2.250 2.795 ;
        RECT 2.510 0.710 2.680 1.095 ;
        RECT 2.080 0.925 2.680 1.095 ;
        RECT 2.080 2.495 2.825 2.795 ;
        RECT 2.510 0.710 3.695 0.880 ;
        RECT 3.760 0.710 3.770 0.945 ;
        RECT 3.835 0.775 4.360 0.945 ;
        RECT 4.425 0.710 4.435 0.945 ;
        RECT 4.500 0.710 5.300 0.880 ;
        RECT 5.130 0.525 5.300 0.960 ;
        RECT 5.130 0.525 7.440 0.695 ;
        RECT 7.650 0.660 9.470 0.830 ;
        RECT 9.300 0.660 9.470 2.435 ;
        RECT 9.045 2.265 9.470 2.435 ;
        RECT 7.575 0.595 7.585 0.829 ;
        RECT 7.585 0.605 7.595 0.829 ;
        RECT 7.595 0.615 7.605 0.829 ;
        RECT 7.605 0.625 7.615 0.829 ;
        RECT 7.615 0.635 7.625 0.829 ;
        RECT 7.625 0.645 7.635 0.829 ;
        RECT 7.635 0.655 7.645 0.829 ;
        RECT 7.645 0.660 7.651 0.830 ;
        RECT 7.515 0.535 7.525 0.769 ;
        RECT 7.525 0.545 7.535 0.779 ;
        RECT 7.535 0.555 7.545 0.789 ;
        RECT 7.545 0.565 7.555 0.799 ;
        RECT 7.555 0.575 7.565 0.809 ;
        RECT 7.565 0.585 7.575 0.819 ;
        RECT 7.440 0.525 7.450 0.695 ;
        RECT 7.450 0.525 7.460 0.705 ;
        RECT 7.460 0.525 7.470 0.715 ;
        RECT 7.470 0.525 7.480 0.725 ;
        RECT 7.480 0.525 7.490 0.735 ;
        RECT 7.490 0.525 7.500 0.745 ;
        RECT 7.500 0.525 7.510 0.755 ;
        RECT 7.510 0.525 7.516 0.765 ;
        RECT 4.435 0.710 4.445 0.934 ;
        RECT 4.445 0.710 4.455 0.924 ;
        RECT 4.455 0.710 4.465 0.914 ;
        RECT 4.465 0.710 4.475 0.904 ;
        RECT 4.475 0.710 4.485 0.894 ;
        RECT 4.485 0.710 4.495 0.884 ;
        RECT 4.495 0.710 4.501 0.880 ;
        RECT 4.360 0.775 4.370 0.945 ;
        RECT 4.370 0.765 4.380 0.945 ;
        RECT 4.380 0.755 4.390 0.945 ;
        RECT 4.390 0.745 4.400 0.945 ;
        RECT 4.400 0.735 4.410 0.945 ;
        RECT 4.410 0.725 4.420 0.945 ;
        RECT 4.420 0.715 4.426 0.945 ;
        RECT 3.770 0.720 3.780 0.944 ;
        RECT 3.780 0.730 3.790 0.944 ;
        RECT 3.790 0.740 3.800 0.944 ;
        RECT 3.800 0.750 3.810 0.944 ;
        RECT 3.810 0.760 3.820 0.944 ;
        RECT 3.820 0.770 3.830 0.944 ;
        RECT 3.830 0.775 3.836 0.945 ;
        RECT 3.695 0.710 3.705 0.880 ;
        RECT 3.705 0.710 3.715 0.890 ;
        RECT 3.715 0.710 3.725 0.900 ;
        RECT 3.725 0.710 3.735 0.910 ;
        RECT 3.735 0.710 3.745 0.920 ;
        RECT 3.745 0.710 3.755 0.930 ;
        RECT 3.755 0.710 3.761 0.940 ;
        RECT 6.185 2.605 6.360 2.775 ;
        RECT 6.530 3.020 7.015 3.190 ;
        RECT 8.175 2.800 8.345 3.140 ;
        RECT 7.310 2.800 8.345 2.970 ;
        RECT 8.175 2.970 9.625 3.140 ;
        RECT 7.235 2.800 7.245 3.034 ;
        RECT 7.245 2.800 7.255 3.024 ;
        RECT 7.255 2.800 7.265 3.014 ;
        RECT 7.265 2.800 7.275 3.004 ;
        RECT 7.275 2.800 7.285 2.994 ;
        RECT 7.285 2.800 7.295 2.984 ;
        RECT 7.295 2.800 7.305 2.974 ;
        RECT 7.305 2.800 7.311 2.970 ;
        RECT 7.090 2.945 7.100 3.179 ;
        RECT 7.100 2.935 7.110 3.169 ;
        RECT 7.110 2.925 7.120 3.159 ;
        RECT 7.120 2.915 7.130 3.149 ;
        RECT 7.130 2.905 7.140 3.139 ;
        RECT 7.140 2.895 7.150 3.129 ;
        RECT 7.150 2.885 7.160 3.119 ;
        RECT 7.160 2.875 7.170 3.109 ;
        RECT 7.170 2.865 7.180 3.099 ;
        RECT 7.180 2.855 7.190 3.089 ;
        RECT 7.190 2.845 7.200 3.079 ;
        RECT 7.200 2.835 7.210 3.069 ;
        RECT 7.210 2.825 7.220 3.059 ;
        RECT 7.220 2.815 7.230 3.049 ;
        RECT 7.230 2.805 7.236 3.045 ;
        RECT 7.015 3.020 7.025 3.190 ;
        RECT 7.025 3.010 7.035 3.190 ;
        RECT 7.035 3.000 7.045 3.190 ;
        RECT 7.045 2.990 7.055 3.190 ;
        RECT 7.055 2.980 7.065 3.190 ;
        RECT 7.065 2.970 7.075 3.190 ;
        RECT 7.075 2.960 7.085 3.190 ;
        RECT 7.085 2.950 7.091 3.190 ;
        RECT 6.575 1.290 6.585 2.464 ;
        RECT 6.585 1.290 6.595 2.454 ;
        RECT 6.595 1.290 6.605 2.444 ;
        RECT 6.605 1.290 6.615 2.434 ;
        RECT 6.615 1.290 6.625 2.424 ;
        RECT 6.625 1.290 6.635 2.414 ;
        RECT 6.635 1.290 6.645 2.404 ;
        RECT 6.645 1.290 6.655 2.394 ;
        RECT 6.655 1.290 6.665 2.384 ;
        RECT 6.665 1.290 6.675 2.374 ;
        RECT 6.675 1.290 6.685 2.364 ;
        RECT 6.685 1.290 6.695 2.354 ;
        RECT 6.695 1.290 6.705 2.344 ;
        RECT 6.705 1.290 6.715 2.334 ;
        RECT 6.715 1.290 6.725 2.324 ;
        RECT 6.725 1.290 6.735 2.314 ;
        RECT 6.735 1.290 6.745 2.304 ;
        RECT 6.530 2.275 6.540 2.509 ;
        RECT 6.540 2.265 6.550 2.499 ;
        RECT 6.550 2.255 6.560 2.489 ;
        RECT 6.560 2.245 6.570 2.479 ;
        RECT 6.570 2.235 6.576 2.475 ;
        RECT 6.360 2.445 6.370 3.189 ;
        RECT 6.370 2.435 6.380 3.189 ;
        RECT 6.380 2.425 6.390 3.189 ;
        RECT 6.390 2.415 6.400 3.189 ;
        RECT 6.400 2.405 6.410 3.189 ;
        RECT 6.410 2.395 6.420 3.189 ;
        RECT 6.420 2.385 6.430 3.189 ;
        RECT 6.430 2.375 6.440 3.189 ;
        RECT 6.440 2.365 6.450 3.189 ;
        RECT 6.450 2.355 6.460 3.189 ;
        RECT 6.460 2.345 6.470 3.189 ;
        RECT 6.470 2.335 6.480 3.189 ;
        RECT 6.480 2.325 6.490 3.189 ;
        RECT 6.490 2.315 6.500 3.189 ;
        RECT 6.500 2.305 6.510 3.189 ;
        RECT 6.510 2.295 6.520 3.189 ;
        RECT 6.520 2.285 6.530 3.189 ;
        RECT 8.690 1.010 8.860 2.790 ;
        RECT 8.590 2.490 8.860 2.790 ;
        RECT 8.690 1.010 8.950 1.310 ;
        RECT 10.810 1.520 10.980 2.790 ;
        RECT 8.590 2.620 10.980 2.790 ;
        RECT 10.810 1.520 11.400 1.820 ;
  END 
END FAHD2XHT

MACRO DEL2HDMXSPGHT
  CLASS  CORE ;
  FOREIGN DEL2HDMXSPGHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 0.345 0.425 0.885 3.085 ;
      LAYER V7 ;
        RECT 0.435 1.255 0.795 1.615 ;
      LAYER M7 ;
        RECT 0.255 1.245 0.980 1.625 ;
      LAYER V6 ;
        RECT 0.520 1.340 0.710 1.530 ;
      LAYER M4 ;
        RECT 0.515 1.255 0.715 2.030 ;
      LAYER V3 ;
        RECT 0.520 1.750 0.710 1.940 ;
      LAYER M3 ;
        RECT 0.105 1.660 0.820 2.030 ;
      LAYER V2 ;
        RECT 0.110 1.750 0.300 1.940 ;
      LAYER M2 ;
        RECT 0.105 1.625 0.305 2.865 ;
      LAYER V1 ;
        RECT 0.110 2.570 0.300 2.760 ;
      LAYER M1 ;
        RECT 0.095 2.470 0.510 2.865 ;
      LAYER M6 ;
        RECT 0.515 0.325 0.715 2.110 ;
      LAYER V5 ;
        RECT 0.520 1.340 0.710 1.530 ;
      LAYER M5 ;
        RECT 0.255 1.335 0.980 1.535 ;
      LAYER V4 ;
        RECT 0.520 1.340 0.710 1.530 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 -0.300 0.860 1.360 ;
        RECT 2.420 -0.300 2.590 0.870 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 1.985 0.325 2.525 3.080 ;
      LAYER V7 ;
        RECT 2.075 0.435 2.435 0.795 ;
      LAYER M7 ;
        RECT 1.935 0.425 3.050 0.805 ;
      LAYER V6 ;
        RECT 2.160 0.520 2.350 0.710 ;
      LAYER M4 ;
        RECT 2.565 0.420 2.765 1.210 ;
      LAYER V3 ;
        RECT 2.570 0.930 2.760 1.120 ;
      LAYER M3 ;
        RECT 2.450 0.840 3.175 1.210 ;
      LAYER V2 ;
        RECT 2.980 0.930 3.170 1.120 ;
      LAYER M2 ;
        RECT 2.975 0.825 3.175 1.670 ;
      LAYER V1 ;
        RECT 2.980 1.340 3.170 1.530 ;
      LAYER M1 ;
        RECT 2.940 0.720 3.110 2.470 ;
        RECT 2.940 1.250 3.180 1.600 ;
      LAYER M6 ;
        RECT 2.155 0.325 2.355 2.110 ;
      LAYER V5 ;
        RECT 2.160 0.520 2.350 0.710 ;
      LAYER M5 ;
        RECT 1.935 0.515 3.050 0.715 ;
      LAYER V4 ;
        RECT 2.570 0.520 2.760 0.710 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.100 0.860 3.990 ;
        RECT 2.355 2.500 2.655 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.540 1.170 1.840 ;
        RECT 1.350 1.060 1.520 2.280 ;
        RECT 1.350 1.520 2.175 1.820 ;
        RECT 1.760 0.570 1.930 1.220 ;
        RECT 1.760 2.055 1.930 2.800 ;
        RECT 1.760 1.050 2.760 1.220 ;
        RECT 2.590 1.050 2.760 2.225 ;
        RECT 1.760 2.055 2.760 2.225 ;
  END 
END DEL2HDMXSPGHT

MACRO BUFHDMXHT
  CLASS  CORE ;
  FOREIGN BUFHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.510 2.885 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.210 1.060 1.380 2.280 ;
        RECT 1.210 1.265 1.540 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.100 0.860 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.030 1.755 ;
        RECT 0.860 1.520 1.030 1.820 ;
  END 
END BUFHDMXHT

MACRO BUFTSHD16XHT
  CLASS  CORE ;
  FOREIGN BUFTSHD16XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.630 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 14.350 1.575 17.530 1.745 ;
        RECT 17.315 1.575 17.530 2.015 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.675 0.535 2.045 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.055 ;
        RECT 1.665 -0.300 1.965 0.715 ;
        RECT 5.445 -0.300 5.745 1.055 ;
        RECT 6.485 -0.300 6.785 1.055 ;
        RECT 7.525 -0.300 7.825 1.055 ;
        RECT 8.565 -0.300 8.865 1.055 ;
        RECT 9.605 -0.300 9.905 1.055 ;
        RECT 10.645 -0.300 10.945 1.055 ;
        RECT 11.685 -0.300 11.985 1.055 ;
        RECT 12.725 -0.300 13.025 1.055 ;
        RECT 13.985 -0.300 14.285 0.715 ;
        RECT 15.025 -0.300 15.325 0.760 ;
        RECT 16.065 -0.300 16.365 0.760 ;
        RECT 17.105 -0.300 17.405 1.055 ;
        RECT 0.000 -0.300 17.630 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 4.990 0.720 5.160 2.960 ;
        RECT 5.965 0.785 6.265 2.895 ;
        RECT 5.965 1.360 7.305 2.005 ;
        RECT 7.005 0.785 7.305 2.895 ;
        RECT 8.045 0.785 8.345 2.895 ;
        RECT 8.045 1.360 9.385 2.005 ;
        RECT 9.085 0.785 9.385 2.895 ;
        RECT 10.125 0.785 10.425 2.895 ;
        RECT 10.125 1.360 11.465 2.005 ;
        RECT 11.165 0.785 11.465 2.895 ;
        RECT 12.205 0.760 12.505 2.895 ;
        RECT 4.990 1.360 13.480 1.980 ;
        RECT 13.300 0.720 13.480 2.965 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.635 0.925 3.990 ;
        RECT 1.665 2.635 1.965 3.990 ;
        RECT 5.445 2.295 5.745 3.990 ;
        RECT 6.485 2.295 6.785 3.990 ;
        RECT 7.525 2.295 7.825 3.990 ;
        RECT 8.565 2.295 8.865 3.990 ;
        RECT 9.605 2.295 9.905 3.990 ;
        RECT 10.645 2.295 10.945 3.990 ;
        RECT 11.685 2.295 11.985 3.990 ;
        RECT 12.725 2.295 13.025 3.990 ;
        RECT 13.985 2.570 14.285 3.990 ;
        RECT 15.025 2.295 15.325 3.990 ;
        RECT 16.065 2.295 16.365 3.990 ;
        RECT 17.105 2.295 17.405 3.990 ;
        RECT 0.000 3.390 17.630 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.160 0.610 0.350 1.495 ;
        RECT 0.160 2.225 0.350 3.205 ;
        RECT 0.160 1.305 1.015 1.495 ;
        RECT 0.825 1.305 1.015 2.415 ;
        RECT 0.160 2.225 1.015 2.415 ;
        RECT 2.325 1.495 2.625 1.985 ;
        RECT 0.825 1.815 3.460 1.985 ;
        RECT 1.210 0.660 1.380 1.300 ;
        RECT 2.325 0.725 2.625 1.300 ;
        RECT 2.705 2.185 3.005 2.695 ;
        RECT 3.570 1.020 3.740 1.445 ;
        RECT 1.210 1.130 3.740 1.300 ;
        RECT 3.745 2.185 4.045 2.695 ;
        RECT 3.570 1.275 4.440 1.445 ;
        RECT 4.270 1.275 4.440 2.355 ;
        RECT 2.705 2.185 4.440 2.355 ;
        RECT 1.205 2.165 1.385 3.145 ;
        RECT 1.205 2.165 2.435 2.365 ;
        RECT 2.235 2.165 2.435 3.095 ;
        RECT 3.225 2.685 3.525 3.095 ;
        RECT 2.985 0.585 4.325 0.755 ;
        RECT 4.025 0.585 4.325 1.095 ;
        RECT 4.025 0.915 4.790 1.095 ;
        RECT 4.620 0.915 4.790 3.095 ;
        RECT 2.235 2.895 4.790 3.095 ;
        RECT 13.675 1.180 13.855 1.570 ;
        RECT 14.570 0.720 14.740 1.360 ;
        RECT 15.610 0.720 15.780 1.360 ;
        RECT 16.640 0.720 16.820 1.360 ;
        RECT 13.675 1.180 16.820 1.360 ;
        RECT 13.675 1.770 13.855 2.105 ;
        RECT 14.550 1.925 14.750 2.960 ;
        RECT 15.595 1.925 15.795 2.960 ;
        RECT 13.675 1.925 16.825 2.105 ;
        RECT 16.645 1.925 16.825 2.960 ;
  END 
END BUFTSHD16XHT

MACRO BUFCLKHD6XHT
  CLASS  CORE ;
  FOREIGN BUFCLKHD6XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.510 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.420 1.625 1.245 1.950 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.245 -0.300 0.545 1.225 ;
        RECT 1.365 -0.300 1.665 1.085 ;
        RECT 2.405 -0.300 2.705 1.085 ;
        RECT 3.445 -0.300 3.745 1.085 ;
        RECT 0.000 -0.300 4.510 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.950 0.980 2.120 1.435 ;
        RECT 1.950 1.965 2.120 2.960 ;
        RECT 2.925 1.045 3.225 1.435 ;
        RECT 2.925 1.965 3.225 2.960 ;
        RECT 1.950 1.265 4.265 1.435 ;
        RECT 3.550 1.265 4.265 2.270 ;
        RECT 1.950 1.965 4.265 2.270 ;
        RECT 3.965 1.045 4.265 2.960 ;
        RECT 3.960 1.265 4.265 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.245 2.325 0.545 3.990 ;
        RECT 1.285 2.665 1.585 3.990 ;
        RECT 2.405 2.485 2.705 3.990 ;
        RECT 3.445 2.485 3.745 3.990 ;
        RECT 0.000 3.390 4.510 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.830 1.060 1.000 1.445 ;
        RECT 0.830 2.145 1.000 2.790 ;
        RECT 0.830 1.275 1.695 1.445 ;
        RECT 1.525 1.275 1.695 2.365 ;
        RECT 0.830 2.145 1.695 2.365 ;
        RECT 1.525 1.615 3.360 1.785 ;
  END 
END BUFCLKHD6XHT

MACRO BUFCLKHD4XHT
  CLASS  CORE ;
  FOREIGN BUFCLKHD4XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.625 0.585 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.705 -0.300 1.005 1.055 ;
        RECT 1.750 -0.300 2.050 1.055 ;
        RECT 2.790 -0.300 3.090 1.045 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.295 1.265 2.770 1.405 ;
        RECT 1.295 1.050 1.465 1.405 ;
        RECT 1.230 1.935 1.530 2.960 ;
        RECT 2.225 1.235 2.505 2.115 ;
        RECT 1.230 1.935 2.570 2.115 ;
        RECT 2.335 1.050 2.505 2.960 ;
        RECT 1.295 1.235 2.505 1.405 ;
        RECT 2.270 1.265 2.570 2.960 ;
        RECT 2.225 1.265 2.770 2.100 ;
        RECT 1.230 1.935 2.770 2.100 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.705 2.635 1.005 3.990 ;
        RECT 1.750 2.295 2.050 3.990 ;
        RECT 2.790 2.295 3.090 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 1.445 ;
        RECT 0.170 2.195 0.340 3.175 ;
        RECT 0.170 1.275 1.040 1.445 ;
        RECT 0.870 1.275 1.040 2.365 ;
        RECT 0.170 2.195 1.040 2.365 ;
        RECT 0.870 1.585 2.030 1.755 ;
  END 
END BUFCLKHD4XHT

MACRO BUFCLKHD12XHT
  CLASS  CORE ;
  FOREIGN BUFCLKHD12XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.560 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.360 1.595 1.195 1.950 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.790 -0.300 1.090 1.065 ;
        RECT 1.830 -0.300 2.130 1.065 ;
        RECT 2.870 -0.300 3.170 1.065 ;
        RECT 3.910 -0.300 4.210 1.065 ;
        RECT 4.950 -0.300 5.250 1.055 ;
        RECT 5.990 -0.300 6.290 1.055 ;
        RECT 0.000 -0.300 6.560 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.350 1.115 2.650 1.450 ;
        RECT 2.350 1.980 2.650 2.895 ;
        RECT 3.390 1.115 3.690 1.450 ;
        RECT 3.390 1.980 3.690 2.895 ;
        RECT 4.430 1.115 4.730 1.450 ;
        RECT 4.430 1.980 4.730 2.895 ;
        RECT 4.430 1.235 6.195 1.450 ;
        RECT 2.350 1.245 6.195 1.450 ;
        RECT 5.470 1.125 5.770 2.895 ;
        RECT 5.175 1.235 6.195 2.315 ;
        RECT 2.350 1.980 6.195 2.315 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.790 2.635 1.090 3.990 ;
        RECT 1.830 2.295 2.130 3.990 ;
        RECT 2.870 2.635 3.170 3.990 ;
        RECT 3.910 2.635 4.210 3.990 ;
        RECT 4.950 2.615 5.250 3.990 ;
        RECT 5.990 2.615 6.290 3.990 ;
        RECT 0.000 3.390 6.560 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.335 1.060 0.505 1.415 ;
        RECT 0.335 2.170 0.505 3.150 ;
        RECT 0.335 1.245 1.545 1.415 ;
        RECT 0.335 2.170 1.545 2.340 ;
        RECT 1.375 1.060 1.545 2.960 ;
        RECT 1.375 1.630 4.945 1.800 ;
  END 
END BUFCLKHD12XHT

MACRO AOI22B2HD2XHT
  CLASS  CORE ;
  FOREIGN AOI22B2HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.515 0.310 2.425 ;
        RECT 0.100 1.515 0.535 1.820 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.770 1.585 3.180 2.050 ;
        RECT 4.395 1.520 4.565 2.050 ;
        RECT 2.770 1.880 4.565 2.050 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.500 1.330 4.065 1.700 ;
    END
  END D
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.845 2.670 1.190 3.180 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.275 ;
        RECT 1.255 -0.300 1.555 1.295 ;
        RECT 2.520 -0.300 2.820 1.055 ;
        RECT 4.510 -0.300 4.810 1.055 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 0.845 2.145 1.205 ;
        RECT 1.975 0.720 2.145 1.405 ;
        RECT 1.975 1.935 2.145 2.620 ;
        RECT 2.240 1.235 2.410 2.105 ;
        RECT 1.975 1.935 2.410 2.105 ;
        RECT 3.110 0.940 3.285 1.405 ;
        RECT 1.975 1.235 3.285 1.405 ;
        RECT 3.535 0.480 3.705 1.120 ;
        RECT 3.110 0.940 3.705 1.120 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.905 0.405 3.990 ;
        RECT 2.950 2.635 3.250 3.990 ;
        RECT 3.990 2.635 4.290 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.730 1.060 0.900 1.755 ;
        RECT 1.025 1.585 1.195 2.280 ;
        RECT 0.730 1.585 2.030 1.755 ;
        RECT 1.455 2.570 1.625 3.210 ;
        RECT 1.455 2.815 2.665 2.985 ;
        RECT 2.495 2.295 2.665 3.210 ;
        RECT 2.430 2.295 2.730 2.465 ;
        RECT 3.535 2.230 3.705 3.210 ;
        RECT 2.575 2.230 4.745 2.400 ;
        RECT 4.575 2.230 4.745 3.210 ;
  END 
END AOI22B2HD2XHT

MACRO AOI222HDMXHT
  CLASS  CORE ;
  FOREIGN AOI222HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.740 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.540 0.520 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.825 1.615 1.285 1.955 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.085 1.595 2.665 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.640 0.510 2.125 0.925 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.035 0.510 3.655 0.940 ;
    END
  END E
  PIN F
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.665 1.530 4.000 2.020 ;
    END
  END F
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.295 ;
        RECT 2.555 -0.300 2.855 0.945 ;
        RECT 4.870 -0.300 5.040 1.210 ;
        RECT 0.000 -0.300 5.740 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.020 2.045 5.230 2.425 ;
        RECT 5.390 1.060 5.585 1.360 ;
        RECT 5.415 1.060 5.585 2.215 ;
        RECT 5.020 2.045 5.585 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.355 0.405 3.990 ;
        RECT 1.175 2.830 1.475 3.990 ;
        RECT 4.705 2.715 5.005 3.990 ;
        RECT 0.000 3.390 5.740 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 2.210 0.860 2.850 ;
        RECT 0.690 2.480 2.505 2.650 ;
        RECT 1.685 2.130 2.960 2.300 ;
        RECT 2.790 2.130 2.960 2.970 ;
        RECT 3.830 2.290 4.000 2.970 ;
        RECT 2.790 2.800 4.000 2.970 ;
        RECT 3.310 1.125 3.480 2.620 ;
        RECT 3.840 0.705 4.010 1.295 ;
        RECT 1.200 1.125 4.010 1.295 ;
        RECT 3.840 0.705 4.665 0.875 ;
        RECT 4.290 1.060 4.510 1.360 ;
        RECT 4.340 1.060 4.510 2.280 ;
        RECT 4.340 1.585 5.235 1.755 ;
  END 
END AOI222HDMXHT

MACRO AND2CLKHD4XHT
  CLASS  CORE ;
  FOREIGN AND2CLKHD4XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.040 1.260 1.540 1.730 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.510 2.220 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.145 -0.300 1.445 0.865 ;
        RECT 2.225 -0.300 2.525 1.095 ;
        RECT 3.265 -0.300 3.565 1.095 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.720 1.060 2.005 1.445 ;
        RECT 1.705 2.285 2.005 2.925 ;
        RECT 1.720 1.275 3.180 1.445 ;
        RECT 2.745 1.060 3.045 2.960 ;
        RECT 2.560 1.275 3.180 2.455 ;
        RECT 1.705 2.285 3.180 2.455 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.635 0.405 3.990 ;
        RECT 1.185 2.635 1.485 3.990 ;
        RECT 2.225 2.635 2.525 3.990 ;
        RECT 3.265 2.635 3.565 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.785 0.405 1.295 ;
        RECT 0.105 1.125 0.860 1.295 ;
        RECT 0.690 1.125 0.860 2.960 ;
        RECT 1.720 1.625 1.895 2.105 ;
        RECT 0.690 1.935 1.895 2.105 ;
        RECT 1.720 1.625 2.360 1.795 ;
  END 
END AND2CLKHD4XHT

MACRO AND2CLKHD3XHT
  CLASS  CORE ;
  FOREIGN AND2CLKHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.170 1.235 1.540 1.730 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.640 2.120 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.275 -0.300 1.575 0.875 ;
        RECT 2.355 -0.300 2.655 1.095 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.835 1.060 2.135 1.445 ;
        RECT 1.835 2.285 2.135 2.920 ;
        RECT 1.835 1.275 3.180 1.445 ;
        RECT 1.835 2.285 3.180 2.455 ;
        RECT 2.835 1.060 3.180 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.235 2.605 0.535 3.990 ;
        RECT 1.315 2.635 1.615 3.990 ;
        RECT 2.355 2.635 2.655 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.235 1.125 0.990 1.295 ;
        RECT 0.820 1.125 0.990 2.960 ;
        RECT 1.720 1.625 1.890 2.105 ;
        RECT 0.820 1.935 1.890 2.105 ;
        RECT 1.720 1.625 2.360 1.795 ;
  END 
END AND2CLKHD3XHT

MACRO AND2CLKHD2XHT
  CLASS  CORE ;
  FOREIGN AND2CLKHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.715 2.800 1.235 3.185 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.640 2.065 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.325 -0.300 1.625 1.095 ;
        RECT 2.390 -0.300 2.690 1.095 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.935 1.060 2.170 2.960 ;
        RECT 1.935 1.330 2.425 2.115 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.235 2.545 0.535 3.990 ;
        RECT 1.415 2.230 1.585 3.990 ;
        RECT 2.390 2.295 2.690 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.235 1.125 1.055 1.295 ;
        RECT 0.885 1.125 1.055 2.620 ;
        RECT 0.820 1.980 1.055 2.620 ;
        RECT 0.885 1.520 1.755 1.820 ;
  END 
END AND2CLKHD2XHT

MACRO AND2CLKHD1XHT
  CLASS  CORE ;
  FOREIGN AND2CLKHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.710 2.395 1.330 2.825 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.475 0.445 2.065 ;
        RECT 0.100 1.475 0.570 1.755 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.105 -0.300 1.405 1.125 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.690 1.060 1.950 1.360 ;
        RECT 1.740 1.060 1.950 2.960 ;
        RECT 1.700 1.980 1.950 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.245 0.405 3.990 ;
        RECT 1.085 3.070 1.385 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 0.920 1.295 ;
        RECT 0.750 1.125 0.920 2.215 ;
        RECT 0.750 1.520 0.925 2.215 ;
        RECT 0.625 2.045 0.925 2.215 ;
        RECT 0.750 1.520 1.550 1.820 ;
  END 
END AND2CLKHD1XHT

MACRO XOR3HDMXHT
  CLASS  CORE ;
  FOREIGN XOR3HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.380 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.180 1.260 4.455 1.820 ;
        RECT 4.475 2.810 6.090 2.980 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.780 1.520 7.280 2.020 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.490 0.475 2.840 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.580 -0.300 0.880 0.605 ;
        RECT 3.115 -0.300 3.285 1.280 ;
        RECT 3.995 -0.300 4.295 0.595 ;
        RECT 6.530 -0.300 6.830 0.745 ;
        RECT 0.000 -0.300 7.380 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.705 0.850 3.875 2.215 ;
        RECT 3.570 2.045 3.875 2.215 ;
        RECT 3.535 0.850 4.000 1.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.715 0.955 3.990 ;
        RECT 3.080 3.095 3.380 3.990 ;
        RECT 3.995 2.875 4.295 3.990 ;
        RECT 6.410 2.715 6.710 3.990 ;
        RECT 0.000 3.390 7.380 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.890 0.985 1.060 2.215 ;
        RECT 0.105 2.045 1.060 2.215 ;
        RECT 1.215 0.570 1.385 1.155 ;
        RECT 0.105 0.985 1.385 1.155 ;
        RECT 1.215 0.570 2.255 0.740 ;
        RECT 2.085 0.570 2.255 2.215 ;
        RECT 2.020 2.045 2.320 2.215 ;
        RECT 2.435 1.370 2.765 1.670 ;
        RECT 2.595 0.980 2.765 2.215 ;
        RECT 2.530 2.045 2.830 2.215 ;
        RECT 1.565 0.920 1.735 2.565 ;
        RECT 3.065 1.520 3.235 2.565 ;
        RECT 1.565 2.395 3.235 2.565 ;
        RECT 3.065 1.520 3.465 1.820 ;
        RECT 4.645 1.060 4.975 1.360 ;
        RECT 4.805 1.060 4.975 2.215 ;
        RECT 4.580 2.045 4.975 2.215 ;
        RECT 3.540 2.460 3.710 2.915 ;
        RECT 1.840 2.745 3.710 2.915 ;
        RECT 5.675 0.955 5.845 2.630 ;
        RECT 3.540 2.460 5.845 2.630 ;
        RECT 5.155 0.605 5.325 2.280 ;
        RECT 5.155 0.605 6.195 0.775 ;
        RECT 6.025 0.605 6.195 1.295 ;
        RECT 6.335 1.125 6.505 2.370 ;
        RECT 6.025 1.125 7.270 1.295 ;
        RECT 6.335 2.200 7.270 2.370 ;
  END 
END XOR3HDMXHT

MACRO XOR3HDLXHT
  CLASS  CORE ;
  FOREIGN XOR3HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.380 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.180 1.260 4.455 1.820 ;
        RECT 4.475 2.810 6.090 2.980 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.780 1.520 7.280 2.020 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.490 0.475 2.840 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.580 -0.300 0.880 0.605 ;
        RECT 3.115 -0.300 3.285 1.280 ;
        RECT 3.995 -0.300 4.295 0.595 ;
        RECT 6.530 -0.300 6.830 0.745 ;
        RECT 0.000 -0.300 7.380 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.535 0.850 3.875 1.280 ;
        RECT 3.705 0.850 3.875 2.215 ;
        RECT 3.570 2.045 3.875 2.215 ;
        RECT 3.535 0.850 4.000 1.200 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.715 0.955 3.990 ;
        RECT 3.080 3.095 3.380 3.990 ;
        RECT 3.995 2.810 4.295 3.990 ;
        RECT 6.410 2.715 6.710 3.990 ;
        RECT 0.000 3.390 7.380 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.890 0.985 1.060 2.215 ;
        RECT 0.105 2.045 1.060 2.215 ;
        RECT 1.215 0.570 1.385 1.155 ;
        RECT 0.105 0.985 1.385 1.155 ;
        RECT 1.215 0.570 2.255 0.740 ;
        RECT 2.085 0.570 2.255 2.215 ;
        RECT 2.020 2.045 2.320 2.215 ;
        RECT 2.435 1.350 2.765 1.650 ;
        RECT 2.595 0.980 2.765 2.215 ;
        RECT 2.530 2.045 2.830 2.215 ;
        RECT 1.565 0.920 1.735 2.565 ;
        RECT 3.065 1.520 3.235 2.565 ;
        RECT 1.565 2.395 3.235 2.565 ;
        RECT 3.065 1.520 3.465 1.820 ;
        RECT 4.645 1.060 4.975 1.360 ;
        RECT 4.805 1.060 4.975 2.215 ;
        RECT 4.580 2.045 4.975 2.215 ;
        RECT 3.540 2.460 3.710 2.915 ;
        RECT 1.840 2.745 3.710 2.915 ;
        RECT 5.675 0.955 5.845 2.630 ;
        RECT 3.540 2.460 5.845 2.630 ;
        RECT 5.155 0.605 5.325 2.280 ;
        RECT 5.155 0.605 6.195 0.775 ;
        RECT 6.025 0.605 6.195 1.295 ;
        RECT 6.335 1.125 6.505 2.370 ;
        RECT 6.025 1.125 7.270 1.295 ;
        RECT 6.335 2.200 7.270 2.370 ;
  END 
END XOR3HDLXHT

MACRO XOR3HD3XHT
  CLASS  CORE ;
  FOREIGN XOR3HD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.610 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.330 1.325 5.760 1.755 ;
        RECT 5.860 2.810 7.320 2.980 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 8.025 1.585 8.515 2.010 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.575 0.585 2.020 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.795 ;
        RECT 3.230 -0.300 3.400 1.120 ;
        RECT 4.240 -0.300 4.540 1.055 ;
        RECT 5.270 -0.300 5.570 1.145 ;
        RECT 7.775 -0.300 8.075 0.790 ;
        RECT 0.000 -0.300 8.610 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.785 0.720 4.005 1.405 ;
        RECT 3.785 1.235 4.995 1.405 ;
        RECT 3.720 2.045 4.995 2.215 ;
        RECT 4.825 0.720 4.995 2.280 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.860 0.925 3.990 ;
        RECT 3.170 3.095 3.470 3.990 ;
        RECT 4.305 2.910 4.475 3.990 ;
        RECT 5.300 2.810 5.600 3.990 ;
        RECT 7.655 2.655 7.955 3.990 ;
        RECT 0.000 3.390 8.610 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.700 0.340 1.345 ;
        RECT 0.170 2.200 0.340 2.865 ;
        RECT 0.870 1.175 1.040 2.370 ;
        RECT 0.170 2.200 1.040 2.370 ;
        RECT 1.165 0.710 1.335 1.345 ;
        RECT 0.170 1.175 1.335 1.345 ;
        RECT 1.165 0.710 2.275 0.880 ;
        RECT 2.105 0.710 2.275 2.215 ;
        RECT 2.070 2.045 2.370 2.215 ;
        RECT 2.455 1.480 2.815 1.780 ;
        RECT 2.645 1.060 2.815 2.215 ;
        RECT 2.580 2.045 2.880 2.215 ;
        RECT 1.585 1.060 1.755 2.565 ;
        RECT 3.090 1.585 3.260 2.565 ;
        RECT 1.585 2.395 3.260 2.565 ;
        RECT 3.090 1.585 4.520 1.755 ;
        RECT 5.810 0.975 6.205 1.145 ;
        RECT 6.035 0.975 6.205 2.215 ;
        RECT 5.810 2.045 6.205 2.215 ;
        RECT 1.925 2.745 2.095 3.075 ;
        RECT 3.720 2.460 3.910 2.915 ;
        RECT 1.925 2.745 3.910 2.915 ;
        RECT 6.905 0.955 7.075 2.630 ;
        RECT 3.720 2.460 7.075 2.630 ;
        RECT 6.385 0.605 6.555 2.280 ;
        RECT 6.385 0.605 7.500 0.775 ;
        RECT 7.330 0.605 7.500 1.215 ;
        RECT 7.565 1.045 7.735 2.390 ;
        RECT 7.330 1.045 8.440 1.215 ;
        RECT 8.270 1.045 8.440 1.360 ;
        RECT 7.565 2.220 8.505 2.390 ;
  END 
END XOR3HD3XHT

MACRO XOR3HD2XHT
  CLASS  CORE ;
  FOREIGN XOR3HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.790 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.200 1.265 4.410 1.755 ;
        RECT 4.200 1.585 4.745 1.755 ;
        RECT 4.770 2.810 6.295 2.980 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.005 1.585 7.560 1.950 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 1.575 0.720 1.755 ;
        RECT 0.510 1.575 0.720 2.020 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.995 ;
        RECT 3.135 -0.300 3.435 1.055 ;
        RECT 4.235 -0.300 4.535 1.055 ;
        RECT 6.735 -0.300 7.035 0.760 ;
        RECT 0.000 -0.300 7.790 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.780 0.720 4.005 1.360 ;
        RECT 3.790 0.720 4.005 2.280 ;
        RECT 3.780 1.980 4.005 2.280 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.630 0.925 3.990 ;
        RECT 3.135 3.095 3.435 3.990 ;
        RECT 4.235 2.975 4.535 3.990 ;
        RECT 6.735 2.485 7.035 3.990 ;
        RECT 0.000 3.390 7.790 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 2.200 0.340 2.865 ;
        RECT 0.105 1.125 0.405 1.345 ;
        RECT 0.915 1.175 1.085 2.370 ;
        RECT 0.170 2.200 1.085 2.370 ;
        RECT 1.240 0.710 1.410 1.345 ;
        RECT 0.105 1.175 1.410 1.345 ;
        RECT 1.240 0.710 2.280 0.880 ;
        RECT 2.110 0.710 2.280 2.215 ;
        RECT 2.075 2.045 2.375 2.215 ;
        RECT 2.460 1.480 2.820 1.780 ;
        RECT 2.650 1.060 2.820 2.215 ;
        RECT 2.585 2.045 2.885 2.215 ;
        RECT 1.590 1.060 1.760 3.145 ;
        RECT 3.120 1.520 3.290 2.565 ;
        RECT 1.590 2.395 3.290 2.565 ;
        RECT 3.120 1.520 3.610 1.820 ;
        RECT 4.850 1.060 5.180 1.360 ;
        RECT 5.010 1.060 5.180 2.280 ;
        RECT 4.850 1.980 5.180 2.280 ;
        RECT 3.685 2.460 3.855 2.915 ;
        RECT 1.940 2.745 3.855 2.915 ;
        RECT 5.880 0.955 6.050 2.630 ;
        RECT 3.685 2.460 6.050 2.630 ;
        RECT 5.360 0.605 5.530 2.280 ;
        RECT 5.360 0.605 6.400 0.775 ;
        RECT 6.230 0.605 6.400 1.110 ;
        RECT 6.540 0.940 6.710 2.305 ;
        RECT 6.230 0.940 7.525 1.110 ;
        RECT 7.355 0.940 7.525 1.360 ;
        RECT 6.540 2.135 7.585 2.305 ;
  END 
END XOR3HD2XHT

MACRO XOR3HD1XHT
  CLASS  CORE ;
  FOREIGN XOR3HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.790 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.200 1.265 4.410 1.755 ;
        RECT 4.200 1.585 4.740 1.755 ;
        RECT 4.610 2.810 6.290 2.980 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.005 1.585 7.580 1.950 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.280 1.585 0.720 1.755 ;
        RECT 0.510 1.585 0.720 2.015 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 -0.300 0.905 0.655 ;
        RECT 3.105 -0.300 3.405 1.055 ;
        RECT 4.195 -0.300 4.495 1.085 ;
        RECT 6.730 -0.300 7.030 0.920 ;
        RECT 0.000 -0.300 7.790 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.745 0.720 4.000 1.360 ;
        RECT 3.820 0.720 4.000 2.215 ;
        RECT 3.685 2.045 4.000 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 2.785 0.905 3.990 ;
        RECT 3.105 3.095 3.465 3.990 ;
        RECT 4.260 2.810 4.430 3.990 ;
        RECT 6.730 2.480 7.030 3.990 ;
        RECT 0.000 3.390 7.790 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.915 1.085 1.085 2.365 ;
        RECT 0.105 2.195 1.085 2.365 ;
        RECT 1.240 0.570 1.410 1.255 ;
        RECT 0.105 1.085 1.410 1.255 ;
        RECT 1.240 0.570 2.280 0.740 ;
        RECT 2.110 0.570 2.280 2.215 ;
        RECT 2.045 2.045 2.345 2.215 ;
        RECT 2.460 1.370 2.790 1.670 ;
        RECT 2.620 0.980 2.790 2.215 ;
        RECT 2.555 2.045 2.855 2.215 ;
        RECT 1.590 0.920 1.760 2.565 ;
        RECT 3.090 1.585 3.260 2.565 ;
        RECT 1.590 2.395 3.260 2.565 ;
        RECT 3.090 1.585 3.640 1.755 ;
        RECT 4.845 1.060 5.175 1.360 ;
        RECT 5.005 1.060 5.175 2.215 ;
        RECT 4.780 2.045 5.175 2.215 ;
        RECT 3.655 2.460 3.825 2.915 ;
        RECT 1.865 2.745 3.825 2.915 ;
        RECT 5.875 0.955 6.045 2.630 ;
        RECT 3.655 2.460 6.045 2.630 ;
        RECT 5.355 0.605 5.530 2.280 ;
        RECT 5.355 0.605 6.395 0.775 ;
        RECT 6.225 0.605 6.395 1.295 ;
        RECT 6.535 1.125 6.705 2.300 ;
        RECT 6.535 2.130 7.580 2.300 ;
        RECT 6.225 1.125 7.585 1.295 ;
  END 
END XOR3HD1XHT

MACRO XOR2HDMXHT
  CLASS  CORE ;
  FOREIGN XOR2HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.395 2.745 2.870 3.180 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 1.585 0.720 1.755 ;
        RECT 0.510 1.585 0.720 2.015 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 -0.300 0.905 0.640 ;
        RECT 3.135 -0.300 3.435 1.300 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.720 0.855 4.000 1.360 ;
        RECT 3.790 0.855 4.000 2.280 ;
        RECT 3.720 1.980 4.000 2.280 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 2.715 0.905 3.990 ;
        RECT 3.170 2.745 3.340 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.165 0.405 2.400 ;
        RECT 0.915 1.020 1.085 2.400 ;
        RECT 0.105 2.195 1.085 2.400 ;
        RECT 1.240 0.585 1.410 1.190 ;
        RECT 0.105 1.020 1.410 1.190 ;
        RECT 1.240 0.585 2.280 0.755 ;
        RECT 2.110 0.585 2.280 2.215 ;
        RECT 2.045 2.045 2.345 2.215 ;
        RECT 2.460 1.430 2.695 1.730 ;
        RECT 2.525 1.125 2.695 2.215 ;
        RECT 2.525 1.125 2.855 1.295 ;
        RECT 2.525 2.045 2.855 2.215 ;
        RECT 1.590 0.955 1.760 2.565 ;
        RECT 3.350 1.520 3.520 2.565 ;
        RECT 1.590 2.395 3.520 2.565 ;
        RECT 3.350 1.520 3.550 1.820 ;
  END 
END XOR2HDMXHT

MACRO XOR2HDLXHT
  CLASS  CORE ;
  FOREIGN XOR2HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.395 2.745 2.870 3.180 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 1.585 0.720 1.755 ;
        RECT 0.510 1.585 0.720 2.015 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 -0.300 0.905 0.640 ;
        RECT 3.100 -0.300 3.400 1.295 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.720 0.855 4.000 1.360 ;
        RECT 3.790 0.855 4.000 2.280 ;
        RECT 3.720 1.980 4.000 2.280 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 2.715 0.905 3.990 ;
        RECT 3.170 2.745 3.340 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.165 0.405 2.400 ;
        RECT 0.915 1.020 1.085 2.400 ;
        RECT 0.105 2.195 1.085 2.400 ;
        RECT 1.240 0.585 1.410 1.190 ;
        RECT 0.105 1.020 1.410 1.190 ;
        RECT 1.240 0.585 2.280 0.755 ;
        RECT 2.110 0.585 2.280 2.215 ;
        RECT 2.045 2.045 2.345 2.215 ;
        RECT 2.460 1.430 2.695 1.730 ;
        RECT 2.525 1.125 2.695 2.215 ;
        RECT 2.525 1.125 2.855 1.295 ;
        RECT 2.525 2.045 2.855 2.215 ;
        RECT 1.590 0.955 1.760 2.565 ;
        RECT 3.350 1.520 3.520 2.565 ;
        RECT 1.590 2.395 3.520 2.565 ;
        RECT 3.350 1.520 3.550 1.820 ;
  END 
END XOR2HDLXHT

MACRO XOR2HD3XHT
  CLASS  CORE ;
  FOREIGN XOR2HD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.910 1.580 3.380 1.955 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.585 0.585 2.015 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.795 ;
        RECT 3.430 -0.300 3.600 1.360 ;
        RECT 4.470 -0.300 4.640 0.780 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.950 0.700 4.120 1.340 ;
        RECT 3.950 1.980 4.120 2.960 ;
        RECT 3.950 1.130 5.230 1.340 ;
        RECT 4.980 1.130 5.230 2.150 ;
        RECT 3.950 1.980 5.230 2.150 ;
        RECT 4.990 0.690 5.230 2.965 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.635 0.925 3.990 ;
        RECT 3.365 2.975 3.665 3.990 ;
        RECT 4.470 2.340 4.640 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.715 0.340 1.395 ;
        RECT 0.170 2.225 0.340 2.910 ;
        RECT 0.870 1.225 1.040 2.395 ;
        RECT 0.170 2.225 1.040 2.395 ;
        RECT 1.125 0.710 1.345 1.395 ;
        RECT 0.170 1.225 1.345 1.395 ;
        RECT 1.125 0.710 2.205 0.880 ;
        RECT 2.035 0.710 2.205 2.320 ;
        RECT 2.035 0.945 2.335 1.115 ;
        RECT 2.035 2.150 2.335 2.320 ;
        RECT 2.385 1.480 2.730 1.780 ;
        RECT 2.560 1.125 2.730 2.305 ;
        RECT 2.560 1.125 3.145 1.295 ;
        RECT 2.560 2.135 3.145 2.305 ;
        RECT 1.580 1.060 1.750 2.675 ;
        RECT 3.570 1.580 3.740 2.675 ;
        RECT 1.580 2.505 3.740 2.675 ;
        RECT 3.570 1.580 4.685 1.755 ;
  END 
END XOR2HD3XHT

MACRO XOR2HD2XHT
  CLASS  CORE ;
  FOREIGN XOR2HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.510 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.995 2.855 2.555 3.180 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 1.585 0.720 1.755 ;
        RECT 0.510 1.585 0.720 2.015 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.995 ;
        RECT 3.030 -0.300 3.330 0.715 ;
        RECT 4.070 -0.300 4.370 1.055 ;
        RECT 0.000 -0.300 4.510 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.615 1.330 4.060 1.360 ;
        RECT 3.695 0.720 3.865 2.960 ;
        RECT 3.615 0.720 3.865 1.360 ;
        RECT 3.695 1.330 3.900 2.960 ;
        RECT 3.615 1.980 3.900 2.960 ;
        RECT 3.695 1.330 4.060 1.540 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.635 0.925 3.990 ;
        RECT 3.030 2.975 3.330 3.990 ;
        RECT 4.100 2.295 4.400 3.990 ;
        RECT 0.000 3.390 4.510 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 1.395 ;
        RECT 0.170 2.195 0.340 2.870 ;
        RECT 0.915 1.225 1.085 2.365 ;
        RECT 0.170 2.195 1.085 2.365 ;
        RECT 1.150 0.710 1.320 1.395 ;
        RECT 0.170 1.225 1.320 1.395 ;
        RECT 1.150 0.710 2.215 0.880 ;
        RECT 2.045 0.710 2.215 2.320 ;
        RECT 2.045 0.945 2.345 1.115 ;
        RECT 2.045 2.150 2.345 2.320 ;
        RECT 2.395 1.480 2.725 1.780 ;
        RECT 2.555 1.125 2.725 2.215 ;
        RECT 2.555 1.125 2.855 1.295 ;
        RECT 2.555 2.045 2.855 2.215 ;
        RECT 1.590 1.060 1.760 2.675 ;
        RECT 3.235 1.520 3.405 2.675 ;
        RECT 1.590 2.505 3.405 2.675 ;
        RECT 3.235 1.520 3.450 1.820 ;
  END 
END XOR2HD2XHT

MACRO XOR2HD1XHT
  CLASS  CORE ;
  FOREIGN XOR2HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.615 2.745 2.165 3.180 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 1.585 0.720 1.755 ;
        RECT 0.510 1.585 0.720 2.015 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 -0.300 0.905 0.695 ;
        RECT 3.135 -0.300 3.435 1.055 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.720 0.720 4.000 1.360 ;
        RECT 3.790 0.720 4.000 2.960 ;
        RECT 3.720 1.980 4.000 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 2.785 0.905 3.990 ;
        RECT 3.105 2.975 3.405 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.915 1.125 1.085 2.365 ;
        RECT 0.105 2.195 1.085 2.365 ;
        RECT 1.240 0.585 1.410 1.295 ;
        RECT 0.105 1.125 1.410 1.295 ;
        RECT 1.240 0.585 2.280 0.755 ;
        RECT 2.110 0.585 2.280 2.215 ;
        RECT 2.045 2.045 2.345 2.215 ;
        RECT 2.460 1.430 2.700 1.730 ;
        RECT 2.530 1.125 2.700 2.215 ;
        RECT 2.530 1.125 2.855 1.295 ;
        RECT 2.530 2.045 2.855 2.215 ;
        RECT 1.590 0.955 1.760 2.565 ;
        RECT 3.350 1.520 3.520 2.565 ;
        RECT 1.590 2.395 3.520 2.565 ;
        RECT 3.350 1.520 3.550 1.820 ;
  END 
END XOR2HD1XHT

MACRO XOR2CLKHD4XHT
  CLASS  CORE ;
  FOREIGN XOR2CLKHD4XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.380 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.125 0.655 4.280 0.660 ;
        RECT 4.035 0.490 4.115 0.670 ;
        RECT 4.035 0.665 4.290 0.670 ;
        RECT 4.045 0.490 4.115 0.680 ;
        RECT 4.045 0.675 4.300 0.680 ;
        RECT 4.055 0.490 4.115 0.690 ;
        RECT 4.055 0.685 4.310 0.690 ;
        RECT 4.065 0.490 4.115 0.700 ;
        RECT 4.065 0.695 4.745 0.700 ;
        RECT 4.075 0.490 4.115 0.710 ;
        RECT 4.075 0.695 4.745 0.710 ;
        RECT 4.085 0.490 4.115 0.720 ;
        RECT 4.085 0.695 4.745 0.720 ;
        RECT 4.095 0.490 4.115 0.730 ;
        RECT 4.095 0.695 4.745 0.730 ;
        RECT 4.105 0.490 4.115 0.740 ;
        RECT 4.105 0.695 4.745 0.740 ;
        RECT 3.125 0.490 4.115 0.660 ;
        RECT 4.115 0.500 4.125 0.750 ;
        RECT 4.115 0.695 4.745 0.750 ;
        RECT 3.125 0.500 4.125 0.660 ;
        RECT 4.125 0.510 4.135 0.760 ;
        RECT 4.125 0.695 4.745 0.760 ;
        RECT 3.125 0.510 4.135 0.660 ;
        RECT 4.135 0.520 4.145 0.770 ;
        RECT 4.135 0.695 4.745 0.770 ;
        RECT 3.125 0.520 4.145 0.660 ;
        RECT 4.145 0.530 4.155 0.780 ;
        RECT 4.145 0.695 4.745 0.780 ;
        RECT 3.125 0.530 4.155 0.660 ;
        RECT 4.155 0.540 4.165 0.790 ;
        RECT 4.155 0.695 4.745 0.790 ;
        RECT 3.125 0.540 4.165 0.660 ;
        RECT 4.165 0.550 4.175 0.800 ;
        RECT 4.165 0.695 4.745 0.800 ;
        RECT 3.125 0.550 4.175 0.660 ;
        RECT 4.175 0.560 4.185 0.810 ;
        RECT 4.175 0.695 4.745 0.810 ;
        RECT 3.125 0.560 4.185 0.660 ;
        RECT 4.185 0.570 4.195 0.820 ;
        RECT 4.185 0.695 4.745 0.820 ;
        RECT 3.125 0.570 4.195 0.660 ;
        RECT 4.195 0.580 4.205 0.830 ;
        RECT 4.195 0.695 4.745 0.830 ;
        RECT 3.125 0.580 4.205 0.660 ;
        RECT 4.205 0.590 4.215 0.840 ;
        RECT 4.205 0.695 4.745 0.840 ;
        RECT 3.125 0.590 4.215 0.660 ;
        RECT 4.215 0.600 4.225 0.850 ;
        RECT 4.215 0.695 4.745 0.850 ;
        RECT 3.125 0.600 4.225 0.660 ;
        RECT 4.225 0.605 4.231 0.859 ;
        RECT 4.225 0.695 4.745 0.859 ;
        RECT 4.230 0.605 4.231 0.865 ;
        RECT 3.125 0.605 4.231 0.660 ;
        RECT 4.230 0.615 4.240 0.865 ;
        RECT 3.125 0.615 4.240 0.660 ;
        RECT 4.230 0.625 4.250 0.865 ;
        RECT 3.125 0.625 4.250 0.660 ;
        RECT 4.230 0.635 4.260 0.865 ;
        RECT 3.125 0.635 4.260 0.660 ;
        RECT 4.230 0.645 4.270 0.865 ;
        RECT 3.125 0.645 4.270 0.660 ;
        RECT 4.230 0.655 4.280 0.865 ;
        RECT 4.035 0.655 4.280 0.670 ;
        RECT 4.230 0.665 4.290 0.865 ;
        RECT 4.045 0.665 4.290 0.680 ;
        RECT 4.230 0.675 4.300 0.865 ;
        RECT 4.055 0.675 4.300 0.690 ;
        RECT 4.230 0.685 4.310 0.865 ;
        RECT 4.065 0.685 4.310 0.700 ;
        RECT 4.230 0.695 4.745 0.865 ;
        RECT 4.850 1.265 5.235 1.755 ;
        RECT 4.755 1.530 5.235 1.755 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.420 1.320 0.970 1.835 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.630 -0.300 0.800 1.110 ;
        RECT 2.485 -0.300 2.785 1.295 ;
        RECT 4.930 -0.300 5.100 0.725 ;
        RECT 5.935 -0.300 6.235 1.080 ;
        RECT 7.040 -0.300 7.210 1.110 ;
        RECT 0.000 -0.300 7.380 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.430 1.350 7.030 1.430 ;
        RECT 5.430 1.060 5.715 1.430 ;
        RECT 5.415 2.295 5.715 2.990 ;
        RECT 5.415 2.295 6.765 2.465 ;
        RECT 6.455 1.055 6.830 1.430 ;
        RECT 6.455 2.045 6.765 2.960 ;
        RECT 6.595 1.055 6.765 2.960 ;
        RECT 6.450 2.295 6.765 2.960 ;
        RECT 6.595 1.055 6.830 2.250 ;
        RECT 5.430 1.260 6.830 1.430 ;
        RECT 6.595 1.350 7.030 2.250 ;
        RECT 6.455 2.045 7.030 2.250 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.600 3.070 0.900 3.990 ;
        RECT 2.485 2.345 2.785 3.990 ;
        RECT 4.820 3.185 5.120 3.990 ;
        RECT 5.935 2.910 6.235 3.990 ;
        RECT 7.040 2.570 7.210 3.990 ;
        RECT 0.000 3.390 7.380 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 2.030 0.340 2.670 ;
        RECT 0.170 2.130 1.320 2.300 ;
        RECT 1.150 0.585 1.320 2.670 ;
        RECT 1.150 0.585 2.295 0.755 ;
        RECT 2.125 0.585 2.295 1.755 ;
        RECT 2.985 0.840 3.165 1.755 ;
        RECT 2.125 1.585 3.165 1.755 ;
        RECT 2.985 0.840 3.860 1.010 ;
        RECT 3.990 0.895 4.000 2.459 ;
        RECT 4.000 0.905 4.010 2.459 ;
        RECT 4.010 0.915 4.020 2.459 ;
        RECT 4.020 0.925 4.030 2.459 ;
        RECT 4.030 0.935 4.040 2.459 ;
        RECT 4.040 0.945 4.050 2.459 ;
        RECT 4.050 0.955 4.060 2.459 ;
        RECT 4.060 0.965 4.070 2.459 ;
        RECT 4.070 0.975 4.080 2.459 ;
        RECT 4.080 0.985 4.090 2.459 ;
        RECT 4.090 0.995 4.100 2.459 ;
        RECT 4.100 1.005 4.110 2.459 ;
        RECT 4.110 1.015 4.120 2.459 ;
        RECT 4.120 1.025 4.130 2.459 ;
        RECT 4.130 1.035 4.140 2.459 ;
        RECT 4.140 1.045 4.150 2.459 ;
        RECT 4.150 1.055 4.160 2.459 ;
        RECT 3.945 0.850 3.955 1.094 ;
        RECT 3.955 0.860 3.965 1.104 ;
        RECT 3.965 0.870 3.975 1.114 ;
        RECT 3.975 0.880 3.985 1.124 ;
        RECT 3.985 0.885 3.991 1.135 ;
        RECT 3.860 0.840 3.870 1.010 ;
        RECT 3.870 0.840 3.880 1.020 ;
        RECT 3.880 0.840 3.890 1.030 ;
        RECT 3.890 0.840 3.900 1.040 ;
        RECT 3.900 0.840 3.910 1.050 ;
        RECT 3.910 0.840 3.920 1.060 ;
        RECT 3.920 0.840 3.930 1.070 ;
        RECT 3.930 0.840 3.940 1.080 ;
        RECT 3.940 0.840 3.946 1.090 ;
        RECT 4.340 1.060 4.510 2.280 ;
        RECT 4.340 1.060 4.670 1.360 ;
        RECT 4.340 2.110 4.735 2.280 ;
        RECT 1.660 1.060 1.830 2.685 ;
        RECT 1.660 1.995 3.610 2.165 ;
        RECT 3.440 1.190 3.610 2.825 ;
        RECT 3.405 1.190 3.705 1.360 ;
        RECT 4.985 1.935 5.175 2.825 ;
        RECT 3.440 2.655 5.175 2.825 ;
        RECT 5.415 1.665 5.650 2.115 ;
        RECT 4.985 1.935 5.650 2.115 ;
        RECT 5.415 1.665 6.395 1.835 ;
  END 
END XOR2CLKHD4XHT

MACRO XOR2CLKHD3XHT
  CLASS  CORE ;
  FOREIGN XOR2CLKHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.170 1.265 3.595 1.755 ;
        RECT 3.075 1.530 3.595 1.755 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.675 0.585 2.015 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.135 ;
        RECT 3.305 -0.300 3.605 1.060 ;
        RECT 4.345 -0.300 4.645 1.070 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.890 1.055 4.060 1.430 ;
        RECT 3.825 2.295 4.125 2.935 ;
        RECT 3.825 2.295 5.230 2.465 ;
        RECT 4.930 1.060 5.230 1.430 ;
        RECT 3.890 1.260 5.230 1.430 ;
        RECT 4.995 1.060 5.230 2.960 ;
        RECT 4.865 2.045 5.230 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.570 0.860 3.990 ;
        RECT 3.305 2.975 3.605 3.990 ;
        RECT 4.345 2.910 4.645 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 1.495 ;
        RECT 0.105 2.200 0.405 3.145 ;
        RECT 0.870 1.325 1.040 2.370 ;
        RECT 0.105 2.200 1.040 2.370 ;
        RECT 1.265 0.655 1.435 1.495 ;
        RECT 0.170 1.325 1.435 1.495 ;
        RECT 1.265 0.655 2.480 0.825 ;
        RECT 2.310 0.655 2.480 2.395 ;
        RECT 2.660 1.060 2.830 2.215 ;
        RECT 2.660 1.060 2.990 1.360 ;
        RECT 2.660 2.045 3.055 2.215 ;
        RECT 1.760 1.060 1.930 2.960 ;
        RECT 3.390 1.935 3.585 2.745 ;
        RECT 1.760 2.575 3.585 2.745 ;
        RECT 3.775 1.665 3.955 2.115 ;
        RECT 3.390 1.935 3.955 2.115 ;
        RECT 3.775 1.665 4.755 1.835 ;
  END 
END XOR2CLKHD3XHT

MACRO XOR2CLKHD1XHT
  CLASS  CORE ;
  FOREIGN XOR2CLKHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.895 1.530 3.215 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.680 0.585 2.015 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.800 ;
        RECT 3.205 -0.300 3.375 1.295 ;
        RECT 3.140 1.125 3.440 1.295 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.760 1.060 4.000 1.360 ;
        RECT 3.790 1.060 4.000 3.055 ;
        RECT 3.760 2.075 4.000 3.055 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.545 0.925 3.990 ;
        RECT 3.175 2.975 3.475 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 1.485 ;
        RECT 0.870 1.315 1.040 2.365 ;
        RECT 0.105 2.195 1.040 2.365 ;
        RECT 1.230 0.680 1.400 1.485 ;
        RECT 0.170 1.315 1.400 1.485 ;
        RECT 1.230 0.680 2.300 0.850 ;
        RECT 2.130 0.680 2.300 2.395 ;
        RECT 2.480 1.060 2.650 2.375 ;
        RECT 2.480 1.060 2.810 1.360 ;
        RECT 2.480 2.205 2.875 2.375 ;
        RECT 1.580 1.060 1.750 2.780 ;
        RECT 3.405 1.540 3.580 2.780 ;
        RECT 1.580 2.610 3.580 2.780 ;
        RECT 3.405 1.540 3.610 1.840 ;
  END 
END XOR2CLKHD1XHT

MACRO XNOR3HDMXHT
  CLASS  CORE ;
  FOREIGN XNOR3HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.790 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.200 1.585 4.410 2.015 ;
        RECT 4.200 1.585 4.685 1.755 ;
        RECT 4.590 2.810 5.715 2.980 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.920 1.540 7.440 1.950 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 1.585 0.720 1.755 ;
        RECT 0.510 1.585 0.720 2.015 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 -0.300 0.905 0.670 ;
        RECT 3.100 -0.300 3.400 1.295 ;
        RECT 4.205 -0.300 4.505 1.295 ;
        RECT 6.675 -0.300 6.975 0.745 ;
        RECT 0.000 -0.300 7.790 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.730 0.860 3.900 2.280 ;
        RECT 3.730 0.860 4.000 1.240 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 2.715 0.905 3.990 ;
        RECT 3.105 3.095 3.405 3.990 ;
        RECT 4.240 2.810 4.410 3.990 ;
        RECT 6.675 2.715 6.975 3.990 ;
        RECT 0.000 3.390 7.790 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.165 0.405 2.365 ;
        RECT 0.915 1.050 1.085 2.365 ;
        RECT 0.105 2.195 1.085 2.365 ;
        RECT 1.240 0.585 1.410 1.220 ;
        RECT 0.105 1.050 1.410 1.220 ;
        RECT 1.240 0.585 2.280 0.755 ;
        RECT 2.110 0.585 2.280 2.215 ;
        RECT 2.045 2.005 2.345 2.215 ;
        RECT 2.460 1.430 2.725 1.730 ;
        RECT 2.555 1.125 2.725 2.215 ;
        RECT 2.555 1.125 2.855 1.295 ;
        RECT 2.555 2.045 2.855 2.215 ;
        RECT 1.590 0.955 1.760 2.565 ;
        RECT 3.350 1.540 3.520 2.565 ;
        RECT 1.590 2.395 3.520 2.565 ;
        RECT 3.350 1.540 3.550 1.840 ;
        RECT 4.725 1.125 5.120 1.295 ;
        RECT 4.950 1.125 5.120 2.215 ;
        RECT 4.725 2.045 5.120 2.215 ;
        RECT 3.765 2.460 3.935 2.915 ;
        RECT 1.865 2.745 3.935 2.915 ;
        RECT 5.820 0.955 5.990 2.630 ;
        RECT 3.765 2.460 5.990 2.630 ;
        RECT 5.300 0.585 5.470 2.280 ;
        RECT 5.300 0.585 6.340 0.755 ;
        RECT 6.170 0.585 6.340 1.295 ;
        RECT 6.495 1.125 6.665 2.300 ;
        RECT 6.170 1.125 7.475 1.295 ;
        RECT 6.495 2.130 7.475 2.300 ;
  END 
END XNOR3HDMXHT

MACRO XNOR3HDLXHT
  CLASS  CORE ;
  FOREIGN XNOR3HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.790 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.200 1.585 4.410 2.015 ;
        RECT 4.200 1.585 4.685 1.755 ;
        RECT 4.590 2.810 5.715 2.980 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.920 1.540 7.440 1.950 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 1.585 0.720 1.755 ;
        RECT 0.510 1.585 0.720 2.015 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 -0.300 0.905 0.670 ;
        RECT 3.110 -0.300 3.410 1.295 ;
        RECT 4.205 -0.300 4.505 1.295 ;
        RECT 6.675 -0.300 6.975 0.745 ;
        RECT 0.000 -0.300 7.790 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.730 0.860 3.900 2.280 ;
        RECT 3.730 0.860 4.000 1.240 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 2.715 0.905 3.990 ;
        RECT 3.105 3.095 3.405 3.990 ;
        RECT 4.240 2.810 4.410 3.990 ;
        RECT 6.675 2.715 6.975 3.990 ;
        RECT 0.000 3.390 7.790 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.165 0.405 2.365 ;
        RECT 0.915 1.050 1.085 2.365 ;
        RECT 0.105 2.195 1.085 2.365 ;
        RECT 1.240 0.585 1.410 1.220 ;
        RECT 0.105 1.050 1.410 1.220 ;
        RECT 1.240 0.585 2.280 0.755 ;
        RECT 2.110 0.585 2.280 2.215 ;
        RECT 2.045 2.040 2.345 2.215 ;
        RECT 2.460 1.430 2.725 1.730 ;
        RECT 2.555 1.125 2.725 2.215 ;
        RECT 2.555 1.125 2.855 1.295 ;
        RECT 2.555 2.045 2.855 2.215 ;
        RECT 1.590 0.955 1.760 2.565 ;
        RECT 3.350 1.540 3.520 2.565 ;
        RECT 1.590 2.395 3.520 2.565 ;
        RECT 3.350 1.540 3.550 1.840 ;
        RECT 4.725 1.125 5.120 1.295 ;
        RECT 4.950 1.125 5.120 2.215 ;
        RECT 4.725 2.045 5.120 2.215 ;
        RECT 3.765 2.460 3.935 2.915 ;
        RECT 1.865 2.745 3.935 2.915 ;
        RECT 5.820 0.955 5.990 2.630 ;
        RECT 3.765 2.460 5.990 2.630 ;
        RECT 5.300 0.585 5.470 2.280 ;
        RECT 5.300 0.585 6.340 0.755 ;
        RECT 6.170 0.585 6.340 1.295 ;
        RECT 6.495 1.125 6.665 2.300 ;
        RECT 6.170 1.125 7.475 1.295 ;
        RECT 6.495 2.130 7.475 2.300 ;
  END 
END XNOR3HDLXHT

MACRO XNOR3HD3XHT
  CLASS  CORE ;
  FOREIGN XNOR3HD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.610 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.285 1.520 5.640 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.830 1.585 8.340 1.950 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 1.580 0.720 2.010 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.935 ;
        RECT 3.155 -0.300 3.455 1.055 ;
        RECT 4.195 -0.300 4.495 1.055 ;
        RECT 5.290 -0.300 5.460 0.780 ;
        RECT 7.625 -0.300 7.925 1.055 ;
        RECT 0.000 -0.300 8.610 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.735 0.715 4.005 1.405 ;
        RECT 3.735 1.235 4.950 1.405 ;
        RECT 4.780 0.715 4.950 2.280 ;
        RECT 3.675 2.110 4.950 2.280 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.635 0.925 3.990 ;
        RECT 3.125 3.095 3.425 3.990 ;
        RECT 4.195 2.975 4.495 3.990 ;
        RECT 5.225 2.975 5.525 3.990 ;
        RECT 7.650 2.480 7.950 3.990 ;
        RECT 0.000 3.390 8.610 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.645 0.340 1.285 ;
        RECT 0.105 2.190 0.405 2.765 ;
        RECT 0.920 1.115 1.090 2.360 ;
        RECT 0.105 2.190 1.090 2.360 ;
        RECT 1.230 0.690 1.400 1.285 ;
        RECT 0.170 1.115 1.400 1.285 ;
        RECT 1.230 0.690 2.300 0.860 ;
        RECT 2.130 0.690 2.300 2.215 ;
        RECT 2.065 2.045 2.365 2.215 ;
        RECT 2.480 1.430 2.745 1.730 ;
        RECT 2.575 1.125 2.745 2.215 ;
        RECT 2.575 1.125 2.875 1.295 ;
        RECT 2.575 2.045 2.875 2.215 ;
        RECT 1.580 1.060 1.750 2.565 ;
        RECT 3.190 1.585 3.360 2.565 ;
        RECT 1.580 2.395 3.360 2.565 ;
        RECT 3.190 1.585 4.475 1.755 ;
        RECT 5.655 1.125 6.050 1.300 ;
        RECT 5.880 1.125 6.050 2.380 ;
        RECT 5.655 2.210 6.050 2.380 ;
        RECT 1.920 2.745 2.090 3.095 ;
        RECT 3.785 2.560 3.955 2.915 ;
        RECT 1.920 2.745 3.955 2.915 ;
        RECT 6.750 0.925 6.920 2.730 ;
        RECT 3.785 2.560 6.920 2.730 ;
        RECT 6.230 0.575 6.400 2.280 ;
        RECT 6.230 0.575 7.270 0.745 ;
        RECT 7.100 0.575 7.270 1.405 ;
        RECT 7.420 1.235 7.590 2.300 ;
        RECT 8.200 1.020 8.500 1.405 ;
        RECT 7.100 1.235 8.500 1.405 ;
        RECT 7.420 2.130 8.505 2.300 ;
  END 
END XNOR3HD3XHT

MACRO XNOR3HD2XHT
  CLASS  CORE ;
  FOREIGN XNOR3HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.790 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.135 1.520 4.475 1.950 ;
        RECT 4.135 1.520 4.700 1.820 ;
        RECT 4.640 2.810 5.955 2.980 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.005 1.585 7.490 1.950 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 1.580 0.720 2.020 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.935 ;
        RECT 3.185 -0.300 3.485 1.055 ;
        RECT 4.225 -0.300 4.525 1.055 ;
        RECT 6.755 -0.300 7.055 0.715 ;
        RECT 0.000 -0.300 7.790 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.770 0.720 3.940 2.280 ;
        RECT 3.770 0.720 4.025 1.195 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.865 0.955 3.990 ;
        RECT 3.155 3.095 3.455 3.990 ;
        RECT 4.290 2.910 4.460 3.990 ;
        RECT 6.755 2.755 7.055 3.990 ;
        RECT 0.000 3.390 7.790 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.065 0.405 1.285 ;
        RECT 0.105 2.205 0.405 2.755 ;
        RECT 0.950 1.115 1.120 2.375 ;
        RECT 0.105 2.205 1.120 2.375 ;
        RECT 1.260 0.585 1.430 1.285 ;
        RECT 0.105 1.115 1.430 1.285 ;
        RECT 1.260 0.585 2.330 0.755 ;
        RECT 2.160 0.585 2.330 2.215 ;
        RECT 2.095 2.045 2.395 2.215 ;
        RECT 2.510 1.430 2.775 1.730 ;
        RECT 2.605 1.125 2.775 2.215 ;
        RECT 2.605 1.125 2.905 1.295 ;
        RECT 2.605 2.045 2.905 2.215 ;
        RECT 1.610 0.955 1.780 2.565 ;
        RECT 3.400 1.520 3.570 2.565 ;
        RECT 1.610 2.395 3.570 2.565 ;
        RECT 3.400 1.520 3.590 1.820 ;
        RECT 4.805 1.125 5.200 1.300 ;
        RECT 5.030 1.125 5.200 2.215 ;
        RECT 4.805 2.045 5.200 2.215 ;
        RECT 3.815 2.460 3.985 2.915 ;
        RECT 1.885 2.745 3.985 2.915 ;
        RECT 5.900 0.925 6.070 2.630 ;
        RECT 3.815 2.460 6.070 2.630 ;
        RECT 5.380 0.575 5.550 2.280 ;
        RECT 5.380 0.575 6.420 0.745 ;
        RECT 6.250 0.575 6.420 1.295 ;
        RECT 6.610 1.125 6.780 2.300 ;
        RECT 6.250 1.125 7.555 1.295 ;
        RECT 6.610 2.130 7.560 2.300 ;
  END 
END XNOR3HD2XHT

MACRO XNOR3HD1XHT
  CLASS  CORE ;
  FOREIGN XNOR3HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.790 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.200 1.520 4.600 2.015 ;
        RECT 4.200 1.520 4.685 1.790 ;
        RECT 4.590 2.810 5.715 2.980 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.970 1.540 7.490 1.950 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.205 1.585 0.720 2.015 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 -0.300 0.905 0.670 ;
        RECT 3.135 -0.300 3.435 1.055 ;
        RECT 4.205 -0.300 4.505 1.295 ;
        RECT 6.675 -0.300 6.975 0.945 ;
        RECT 0.000 -0.300 7.790 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.730 0.720 4.005 2.280 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 2.785 0.905 3.990 ;
        RECT 3.105 3.095 3.405 3.990 ;
        RECT 4.240 2.810 4.410 3.990 ;
        RECT 6.675 2.500 6.975 3.990 ;
        RECT 0.000 3.390 7.790 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.915 1.050 1.085 2.365 ;
        RECT 0.105 2.195 1.085 2.365 ;
        RECT 1.240 0.585 1.410 1.220 ;
        RECT 0.105 1.050 1.410 1.220 ;
        RECT 1.240 0.585 2.280 0.755 ;
        RECT 2.110 0.585 2.280 2.215 ;
        RECT 2.045 2.045 2.345 2.215 ;
        RECT 2.460 1.430 2.725 1.730 ;
        RECT 2.555 1.125 2.725 2.215 ;
        RECT 2.555 1.125 2.855 1.295 ;
        RECT 2.555 2.045 2.855 2.215 ;
        RECT 1.590 0.955 1.760 2.565 ;
        RECT 3.350 1.520 3.520 2.565 ;
        RECT 1.590 2.395 3.520 2.565 ;
        RECT 3.350 1.520 3.550 1.820 ;
        RECT 4.790 1.060 5.120 1.360 ;
        RECT 4.950 1.060 5.120 2.280 ;
        RECT 4.790 1.980 5.120 2.280 ;
        RECT 3.765 2.460 3.935 2.915 ;
        RECT 1.865 2.745 3.935 2.915 ;
        RECT 5.820 0.955 5.990 2.630 ;
        RECT 3.765 2.460 5.990 2.630 ;
        RECT 5.300 0.605 5.470 2.280 ;
        RECT 5.300 0.605 6.340 0.775 ;
        RECT 6.170 0.605 6.340 1.295 ;
        RECT 6.495 1.125 6.665 2.320 ;
        RECT 6.170 1.125 7.525 1.295 ;
        RECT 6.495 2.150 7.525 2.320 ;
  END 
END XNOR3HD1XHT

MACRO XNOR2HDMXHT
  CLASS  CORE ;
  FOREIGN XNOR2HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.345 2.810 2.990 2.980 ;
        RECT 2.475 2.810 2.990 3.180 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 1.585 0.720 1.945 ;
        RECT 0.510 1.585 0.720 2.015 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 -0.300 0.905 0.745 ;
        RECT 3.075 -0.300 3.375 1.295 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.675 1.125 4.000 1.295 ;
        RECT 3.830 1.125 4.000 2.440 ;
        RECT 3.740 2.000 4.000 2.440 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 2.715 0.905 3.990 ;
        RECT 3.170 2.810 3.340 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.165 0.405 2.365 ;
        RECT 0.915 1.125 1.085 2.365 ;
        RECT 0.105 2.195 1.085 2.365 ;
        RECT 1.240 0.605 1.410 1.295 ;
        RECT 0.105 1.125 1.410 1.295 ;
        RECT 1.240 0.605 2.280 0.775 ;
        RECT 2.110 0.605 2.280 2.280 ;
        RECT 2.460 1.125 2.630 2.215 ;
        RECT 2.460 1.125 2.855 1.295 ;
        RECT 2.460 2.045 2.855 2.215 ;
        RECT 1.590 0.955 1.760 2.630 ;
        RECT 3.360 1.540 3.530 2.630 ;
        RECT 1.590 2.460 3.530 2.630 ;
        RECT 3.360 1.540 3.610 1.840 ;
  END 
END XNOR2HDMXHT

MACRO XNOR2HDLXHT
  CLASS  CORE ;
  FOREIGN XNOR2HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.345 2.810 2.990 2.980 ;
        RECT 2.475 2.810 2.990 3.180 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 1.585 0.720 1.945 ;
        RECT 0.510 1.585 0.720 2.015 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 -0.300 0.905 0.695 ;
        RECT 3.075 -0.300 3.375 1.295 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.675 1.125 4.000 1.295 ;
        RECT 3.830 1.125 4.000 2.440 ;
        RECT 3.740 2.000 4.000 2.440 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 2.715 0.905 3.990 ;
        RECT 3.170 2.810 3.340 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.165 0.405 2.365 ;
        RECT 0.915 1.125 1.085 2.365 ;
        RECT 0.105 2.195 1.085 2.365 ;
        RECT 1.240 0.605 1.410 1.295 ;
        RECT 0.105 1.125 1.410 1.295 ;
        RECT 1.240 0.605 2.280 0.775 ;
        RECT 2.110 0.605 2.280 2.280 ;
        RECT 2.460 1.125 2.630 2.215 ;
        RECT 2.460 1.125 2.855 1.295 ;
        RECT 2.460 2.045 2.855 2.215 ;
        RECT 1.590 0.955 1.760 2.630 ;
        RECT 3.360 1.540 3.530 2.630 ;
        RECT 1.590 2.460 3.530 2.630 ;
        RECT 3.360 1.540 3.610 1.840 ;
  END 
END XNOR2HDLXHT

MACRO XNOR2HD3XHT
  CLASS  CORE ;
  FOREIGN XNOR2HD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.315 1.265 3.590 1.755 ;
        RECT 3.125 1.530 3.590 1.755 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.585 2.015 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.940 ;
        RECT 3.335 -0.300 3.635 1.055 ;
        RECT 4.405 -0.300 4.705 1.055 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.950 0.700 4.120 1.405 ;
        RECT 4.120 2.030 4.290 2.990 ;
        RECT 3.950 2.350 4.290 2.990 ;
        RECT 4.120 2.030 5.230 2.230 ;
        RECT 4.990 0.695 5.230 1.405 ;
        RECT 3.950 1.235 5.230 1.405 ;
        RECT 5.020 0.695 5.230 3.010 ;
        RECT 4.990 2.030 5.230 3.010 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.635 0.925 3.990 ;
        RECT 3.365 2.950 3.665 3.990 ;
        RECT 4.470 2.570 4.640 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.710 0.340 1.350 ;
        RECT 0.105 2.195 0.405 2.765 ;
        RECT 0.870 1.180 1.040 2.365 ;
        RECT 0.105 2.195 1.040 2.365 ;
        RECT 1.340 0.605 1.510 1.350 ;
        RECT 0.170 1.180 1.510 1.350 ;
        RECT 1.340 0.605 2.380 0.775 ;
        RECT 2.210 0.605 2.380 2.280 ;
        RECT 2.690 1.060 2.860 2.215 ;
        RECT 2.690 1.060 3.020 1.360 ;
        RECT 2.690 2.045 3.085 2.215 ;
        RECT 1.660 1.980 1.830 2.960 ;
        RECT 1.690 0.955 1.860 2.630 ;
        RECT 1.660 1.980 1.860 2.630 ;
        RECT 3.405 1.935 3.575 2.630 ;
        RECT 1.660 2.460 3.575 2.630 ;
        RECT 3.770 1.585 3.940 2.115 ;
        RECT 3.405 1.935 3.940 2.115 ;
        RECT 3.770 1.585 4.750 1.755 ;
  END 
END XNOR2HD3XHT

MACRO XNOR2HD2XHT
  CLASS  CORE ;
  FOREIGN XNOR2HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.510 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.970 1.265 3.180 1.755 ;
        RECT 2.875 1.530 3.180 1.755 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.585 2.015 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.940 ;
        RECT 3.060 -0.300 3.360 0.715 ;
        RECT 4.100 -0.300 4.400 1.055 ;
        RECT 0.000 -0.300 4.510 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.645 1.175 3.940 1.340 ;
        RECT 3.770 0.700 3.815 2.990 ;
        RECT 3.645 0.700 3.815 1.340 ;
        RECT 3.770 1.175 3.940 2.990 ;
        RECT 3.645 2.350 3.940 2.990 ;
        RECT 3.770 1.675 4.000 2.015 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.585 0.925 3.990 ;
        RECT 3.060 2.975 3.360 3.990 ;
        RECT 4.170 2.230 4.340 3.990 ;
        RECT 0.000 3.390 4.510 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.005 0.340 1.350 ;
        RECT 0.105 2.200 0.405 2.755 ;
        RECT 0.870 1.180 1.040 2.370 ;
        RECT 0.105 2.200 1.040 2.370 ;
        RECT 1.240 0.575 1.410 1.350 ;
        RECT 0.170 1.180 1.410 1.350 ;
        RECT 1.240 0.575 2.280 0.745 ;
        RECT 2.110 0.575 2.280 2.280 ;
        RECT 2.460 1.060 2.630 2.215 ;
        RECT 2.460 1.060 2.790 1.360 ;
        RECT 2.460 2.045 2.855 2.215 ;
        RECT 1.590 0.955 1.760 3.100 ;
        RECT 3.295 1.935 3.465 2.630 ;
        RECT 1.590 2.460 3.465 2.630 ;
        RECT 3.395 1.520 3.590 2.115 ;
        RECT 3.295 1.935 3.590 2.115 ;
  END 
END XNOR2HD2XHT

MACRO XNOR2HD1XHT
  CLASS  CORE ;
  FOREIGN XNOR2HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.345 2.810 2.990 2.980 ;
        RECT 2.970 1.270 3.195 1.820 ;
        RECT 2.825 1.540 3.195 1.820 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 1.585 0.720 2.015 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 -0.300 0.905 0.605 ;
        RECT 3.135 -0.300 3.435 1.055 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.720 0.720 4.000 1.360 ;
        RECT 3.805 0.720 4.000 2.980 ;
        RECT 3.740 2.000 4.000 2.980 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 2.785 0.905 3.990 ;
        RECT 3.170 2.910 3.340 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.915 1.085 1.085 2.365 ;
        RECT 0.105 2.195 1.085 2.365 ;
        RECT 1.240 0.570 1.410 1.255 ;
        RECT 0.105 1.085 1.410 1.255 ;
        RECT 1.240 0.570 2.280 0.740 ;
        RECT 2.110 0.570 2.280 2.280 ;
        RECT 2.460 1.060 2.630 2.215 ;
        RECT 2.460 1.060 2.790 1.360 ;
        RECT 2.460 2.045 2.855 2.215 ;
        RECT 1.590 0.920 1.760 2.630 ;
        RECT 3.375 1.520 3.545 2.630 ;
        RECT 1.590 2.460 3.545 2.630 ;
        RECT 3.375 1.520 3.615 1.820 ;
  END 
END XNOR2HD1XHT

MACRO TIEHHDHT
  CLASS  CORE ;
  FOREIGN TIEHHDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.230 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.165 -0.300 0.465 1.295 ;
        RECT 0.000 -0.300 1.230 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.820 1.980 1.130 2.425 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.165 2.045 0.465 3.990 ;
        RECT 0.000 3.390 1.230 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.830 1.060 1.000 1.755 ;
        RECT 0.385 1.585 1.000 1.755 ;
  END 
END TIEHHDHT

MACRO RSLATNHDMXHT
  CLASS  CORE ;
  FOREIGN RSLATNHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.875 1.125 3.045 2.360 ;
        RECT 2.875 1.125 3.175 1.295 ;
        RECT 2.875 2.150 3.340 2.360 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.090 1.235 2.260 2.280 ;
        RECT 2.365 1.125 2.665 1.625 ;
        RECT 2.090 1.235 2.665 1.625 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.485 2.900 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.680 -0.300 0.875 1.360 ;
        RECT 1.805 -0.300 2.105 0.595 ;
        RECT 3.435 -0.300 3.735 0.595 ;
        RECT 4.590 -0.300 4.785 1.295 ;
        RECT 4.405 1.125 4.785 1.295 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.380 1.940 4.820 2.430 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.100 0.860 3.990 ;
        RECT 2.575 2.940 2.875 3.990 ;
        RECT 4.470 2.610 4.640 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.605 1.105 1.775 ;
        RECT 1.400 2.590 1.570 2.940 ;
        RECT 3.290 1.570 3.390 1.870 ;
        RECT 3.565 1.125 3.630 2.760 ;
        RECT 1.400 2.590 3.630 2.760 ;
        RECT 3.580 1.125 3.630 2.835 ;
        RECT 3.565 1.125 4.185 1.295 ;
        RECT 3.630 1.865 3.640 2.835 ;
        RECT 3.640 1.875 3.650 2.835 ;
        RECT 3.650 1.885 3.660 2.835 ;
        RECT 3.660 1.895 3.670 2.835 ;
        RECT 3.670 1.905 3.680 2.835 ;
        RECT 3.680 1.915 3.690 2.835 ;
        RECT 3.690 1.925 3.700 2.835 ;
        RECT 3.700 1.935 3.710 2.835 ;
        RECT 3.710 1.945 3.720 2.835 ;
        RECT 3.720 1.955 3.730 2.835 ;
        RECT 3.730 1.965 3.740 2.835 ;
        RECT 3.740 1.975 3.750 2.835 ;
        RECT 3.460 1.125 3.470 1.939 ;
        RECT 3.470 1.125 3.480 1.949 ;
        RECT 3.480 1.125 3.490 1.959 ;
        RECT 3.490 1.125 3.500 1.969 ;
        RECT 3.500 1.125 3.510 1.979 ;
        RECT 3.510 1.125 3.520 1.989 ;
        RECT 3.520 1.125 3.530 1.999 ;
        RECT 3.530 1.125 3.540 2.009 ;
        RECT 3.540 1.125 3.550 2.019 ;
        RECT 3.550 1.125 3.560 2.029 ;
        RECT 3.560 1.125 3.566 2.039 ;
        RECT 3.390 1.570 3.400 1.870 ;
        RECT 3.400 1.570 3.410 1.880 ;
        RECT 3.410 1.570 3.420 1.890 ;
        RECT 3.420 1.570 3.430 1.900 ;
        RECT 3.430 1.570 3.440 1.910 ;
        RECT 3.440 1.570 3.450 1.920 ;
        RECT 3.450 1.570 3.460 1.930 ;
        RECT 1.145 1.125 1.500 1.295 ;
        RECT 1.330 0.775 1.500 2.215 ;
        RECT 1.330 2.045 1.815 2.215 ;
        RECT 2.285 0.605 2.585 0.945 ;
        RECT 4.240 0.640 4.410 0.945 ;
        RECT 1.330 0.775 4.410 0.945 ;
        RECT 3.810 1.475 3.980 1.775 ;
        RECT 4.990 1.060 5.170 1.645 ;
        RECT 3.810 1.475 5.170 1.645 ;
        RECT 5.000 1.060 5.170 2.910 ;
        RECT 4.990 2.610 5.170 2.910 ;
  END 
END RSLATNHDMXHT

MACRO RSLATNHDLXHT
  CLASS  CORE ;
  FOREIGN RSLATNHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.875 1.125 3.045 2.360 ;
        RECT 2.875 1.125 3.175 1.295 ;
        RECT 2.875 2.150 3.340 2.360 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.090 1.125 2.260 2.280 ;
        RECT 2.090 1.125 2.665 1.540 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.485 2.900 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 1.805 -0.300 2.105 0.595 ;
        RECT 3.435 -0.300 3.735 0.595 ;
        RECT 4.590 -0.300 4.785 1.295 ;
        RECT 4.405 1.125 4.785 1.295 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.380 1.925 4.820 2.430 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.100 0.860 3.990 ;
        RECT 2.575 2.900 2.875 3.990 ;
        RECT 4.470 2.610 4.640 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.605 1.105 1.775 ;
        RECT 1.400 2.540 1.570 2.940 ;
        RECT 3.290 1.570 3.400 1.870 ;
        RECT 1.400 2.540 3.630 2.720 ;
        RECT 3.580 1.125 3.630 2.835 ;
        RECT 3.580 1.125 4.185 1.295 ;
        RECT 3.630 1.865 3.640 2.835 ;
        RECT 3.640 1.875 3.650 2.835 ;
        RECT 3.650 1.885 3.660 2.835 ;
        RECT 3.660 1.895 3.670 2.835 ;
        RECT 3.670 1.905 3.680 2.835 ;
        RECT 3.680 1.915 3.690 2.835 ;
        RECT 3.690 1.925 3.700 2.835 ;
        RECT 3.700 1.935 3.710 2.835 ;
        RECT 3.710 1.945 3.720 2.835 ;
        RECT 3.720 1.955 3.730 2.835 ;
        RECT 3.730 1.965 3.740 2.835 ;
        RECT 3.740 1.975 3.750 2.835 ;
        RECT 3.460 1.125 3.470 1.929 ;
        RECT 3.470 1.125 3.480 1.939 ;
        RECT 3.480 1.125 3.490 1.949 ;
        RECT 3.490 1.125 3.500 1.959 ;
        RECT 3.500 1.125 3.510 1.969 ;
        RECT 3.510 1.125 3.520 1.979 ;
        RECT 3.520 1.125 3.530 1.989 ;
        RECT 3.530 1.125 3.540 1.999 ;
        RECT 3.540 1.125 3.550 2.009 ;
        RECT 3.550 1.125 3.560 2.019 ;
        RECT 3.560 1.125 3.570 2.029 ;
        RECT 3.570 1.125 3.580 2.039 ;
        RECT 3.400 1.570 3.410 1.870 ;
        RECT 3.410 1.570 3.420 1.880 ;
        RECT 3.420 1.570 3.430 1.890 ;
        RECT 3.430 1.570 3.440 1.900 ;
        RECT 3.440 1.570 3.450 1.910 ;
        RECT 3.450 1.570 3.460 1.920 ;
        RECT 1.145 1.125 1.500 1.295 ;
        RECT 1.330 0.775 1.500 2.215 ;
        RECT 1.330 2.045 1.815 2.215 ;
        RECT 2.285 0.755 2.585 0.945 ;
        RECT 4.175 0.640 4.410 0.945 ;
        RECT 1.330 0.775 4.410 0.945 ;
        RECT 3.810 1.475 3.980 1.775 ;
        RECT 4.985 1.060 5.170 1.660 ;
        RECT 3.810 1.475 5.170 1.660 ;
        RECT 5.000 1.060 5.170 2.910 ;
        RECT 4.990 2.595 5.170 2.910 ;
  END 
END RSLATNHDLXHT

MACRO RSLATNHD2XHT
  CLASS  CORE ;
  FOREIGN RSLATNHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.560 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.620 1.125 3.790 2.360 ;
        RECT 3.620 1.125 3.920 1.295 ;
        RECT 3.620 2.045 4.090 2.360 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.310 0.720 2.480 1.475 ;
        RECT 2.310 1.230 2.770 1.475 ;
        RECT 2.560 1.230 2.770 2.255 ;
        RECT 2.560 2.085 2.975 2.255 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.900 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.295 ;
        RECT 1.725 -0.300 2.025 1.055 ;
        RECT 2.920 -0.300 3.090 1.120 ;
        RECT 4.180 -0.300 4.480 0.595 ;
        RECT 5.585 -0.300 5.885 0.995 ;
        RECT 0.000 -0.300 6.560 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.040 2.420 6.460 2.840 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 2.140 0.890 3.990 ;
        RECT 2.155 2.975 2.455 3.990 ;
        RECT 3.195 2.975 3.495 3.990 ;
        RECT 4.235 2.975 4.535 3.990 ;
        RECT 5.545 2.545 5.845 3.990 ;
        RECT 0.000 3.390 6.560 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.605 1.030 1.775 ;
        RECT 0.860 1.540 1.030 1.840 ;
        RECT 1.175 1.125 1.500 1.295 ;
        RECT 1.330 1.125 1.500 1.825 ;
        RECT 1.660 1.655 1.830 2.280 ;
        RECT 1.330 1.655 2.365 1.825 ;
        RECT 3.970 1.535 4.655 1.835 ;
        RECT 4.485 1.125 4.655 2.775 ;
        RECT 4.485 1.980 4.890 2.775 ;
        RECT 1.875 2.605 4.890 2.775 ;
        RECT 4.485 1.125 5.030 1.295 ;
        RECT 3.270 0.775 3.440 1.890 ;
        RECT 2.950 1.590 3.440 1.890 ;
        RECT 3.270 0.775 5.405 0.945 ;
        RECT 5.235 0.775 5.405 1.345 ;
        RECT 5.235 1.175 5.600 1.345 ;
        RECT 5.430 1.175 5.600 1.730 ;
        RECT 4.835 1.540 5.240 1.710 ;
        RECT 5.070 1.540 5.240 2.215 ;
        RECT 6.220 1.060 6.390 2.215 ;
        RECT 5.070 2.045 6.455 2.215 ;
  END 
END RSLATNHD2XHT

MACRO RSLATHDMXHT
  CLASS  CORE ;
  FOREIGN RSLATHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.980 1.125 2.360 1.295 ;
        RECT 2.150 1.125 2.360 2.215 ;
        RECT 2.150 2.045 2.595 2.215 ;
    END
  END Q
  PIN R
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.485 2.900 ;
    END
  END R
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.820 2.470 5.230 2.885 ;
    END
  END S
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.870 1.125 3.050 2.430 ;
        RECT 2.870 2.050 3.220 2.430 ;
        RECT 2.870 1.125 3.305 1.295 ;
    END
  END QN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.580 -0.300 0.880 1.295 ;
        RECT 2.530 -0.300 2.830 0.595 ;
        RECT 4.590 -0.300 4.785 1.295 ;
        RECT 4.405 1.125 4.785 1.295 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.035 0.860 3.990 ;
        RECT 1.695 2.745 1.995 3.990 ;
        RECT 3.420 2.630 3.590 3.990 ;
        RECT 4.470 2.040 4.640 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.510 0.340 2.280 ;
        RECT 0.170 1.605 1.030 1.775 ;
        RECT 0.860 1.540 1.030 1.840 ;
        RECT 1.565 1.520 1.735 2.565 ;
        RECT 1.565 2.395 2.610 2.565 ;
        RECT 2.440 2.395 2.610 2.915 ;
        RECT 2.440 2.745 3.240 2.915 ;
        RECT 3.230 1.570 3.290 1.870 ;
        RECT 3.515 1.125 3.630 2.260 ;
        RECT 3.515 2.090 4.185 2.260 ;
        RECT 3.630 1.125 3.640 1.519 ;
        RECT 3.640 1.125 3.650 1.509 ;
        RECT 3.650 1.125 3.660 1.499 ;
        RECT 3.660 1.125 3.670 1.489 ;
        RECT 3.670 1.125 3.680 1.479 ;
        RECT 3.680 1.125 3.690 1.469 ;
        RECT 3.690 1.125 3.700 1.459 ;
        RECT 3.700 1.125 3.710 1.449 ;
        RECT 3.710 1.125 3.720 1.439 ;
        RECT 3.720 1.125 3.730 1.429 ;
        RECT 3.730 1.125 3.740 1.419 ;
        RECT 3.740 1.125 3.750 1.409 ;
        RECT 3.750 1.125 3.760 1.399 ;
        RECT 3.760 1.125 3.770 1.389 ;
        RECT 3.770 1.125 3.780 1.379 ;
        RECT 3.780 1.125 3.790 1.369 ;
        RECT 3.790 1.125 3.800 1.359 ;
        RECT 3.800 1.125 3.810 1.349 ;
        RECT 3.810 1.125 3.816 1.345 ;
        RECT 3.445 1.415 3.455 2.259 ;
        RECT 3.455 1.405 3.465 2.259 ;
        RECT 3.465 1.395 3.475 2.259 ;
        RECT 3.475 1.385 3.485 2.259 ;
        RECT 3.485 1.375 3.495 2.259 ;
        RECT 3.495 1.365 3.505 2.259 ;
        RECT 3.505 1.355 3.515 2.259 ;
        RECT 3.290 1.570 3.300 1.870 ;
        RECT 3.300 1.560 3.310 1.870 ;
        RECT 3.310 1.550 3.320 1.870 ;
        RECT 3.320 1.540 3.330 1.870 ;
        RECT 3.330 1.530 3.340 1.870 ;
        RECT 3.340 1.520 3.350 1.870 ;
        RECT 3.350 1.510 3.360 1.870 ;
        RECT 3.360 1.500 3.370 1.870 ;
        RECT 3.370 1.490 3.380 1.870 ;
        RECT 3.380 1.480 3.390 1.870 ;
        RECT 3.390 1.470 3.400 1.870 ;
        RECT 3.400 1.460 3.410 1.870 ;
        RECT 3.410 1.450 3.420 1.870 ;
        RECT 3.420 1.440 3.430 1.870 ;
        RECT 3.430 1.430 3.440 1.870 ;
        RECT 3.440 1.420 3.446 1.870 ;
        RECT 1.210 1.125 1.385 2.280 ;
        RECT 1.600 0.775 1.770 1.295 ;
        RECT 1.210 1.125 1.770 1.295 ;
        RECT 2.180 0.540 2.350 0.945 ;
        RECT 4.240 0.640 4.410 0.945 ;
        RECT 1.600 0.775 4.410 0.945 ;
        RECT 3.810 1.610 3.980 1.910 ;
        RECT 3.810 1.610 5.160 1.780 ;
        RECT 4.990 1.060 5.160 2.280 ;
  END 
END RSLATHDMXHT

MACRO TIELHDHT
  CLASS  CORE ;
  FOREIGN TIELHDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.230 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.165 -0.300 0.465 1.295 ;
        RECT 0.000 -0.300 1.230 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.795 0.855 1.130 1.295 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.165 2.045 0.465 3.990 ;
        RECT 0.000 3.390 1.230 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.385 1.585 1.000 1.755 ;
        RECT 0.830 1.585 1.000 2.280 ;
  END 
END TIELHDHT

MACRO RSLATHDLXHT
  CLASS  CORE ;
  FOREIGN RSLATHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.980 1.125 2.360 1.295 ;
        RECT 2.150 1.125 2.360 2.215 ;
        RECT 2.150 2.045 2.595 2.215 ;
    END
  END Q
  PIN R
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.485 2.900 ;
    END
  END R
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.820 2.470 5.230 2.885 ;
    END
  END S
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.870 1.125 3.050 2.430 ;
        RECT 2.870 2.050 3.220 2.430 ;
        RECT 2.870 1.125 3.305 1.295 ;
    END
  END QN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.580 -0.300 0.880 1.295 ;
        RECT 2.530 -0.300 2.830 0.595 ;
        RECT 4.590 -0.300 4.785 1.295 ;
        RECT 4.405 1.125 4.785 1.295 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.035 0.860 3.990 ;
        RECT 1.695 2.745 1.995 3.990 ;
        RECT 3.420 2.630 3.590 3.990 ;
        RECT 4.470 2.040 4.640 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.510 0.340 2.280 ;
        RECT 0.170 1.605 1.030 1.775 ;
        RECT 0.860 1.540 1.030 1.840 ;
        RECT 1.565 1.520 1.735 2.565 ;
        RECT 1.565 2.395 2.610 2.565 ;
        RECT 2.440 2.395 2.610 2.780 ;
        RECT 2.440 2.610 3.240 2.780 ;
        RECT 3.230 1.570 3.290 1.870 ;
        RECT 3.515 1.125 3.630 2.260 ;
        RECT 3.515 2.090 4.185 2.260 ;
        RECT 3.630 1.125 3.640 1.519 ;
        RECT 3.640 1.125 3.650 1.509 ;
        RECT 3.650 1.125 3.660 1.499 ;
        RECT 3.660 1.125 3.670 1.489 ;
        RECT 3.670 1.125 3.680 1.479 ;
        RECT 3.680 1.125 3.690 1.469 ;
        RECT 3.690 1.125 3.700 1.459 ;
        RECT 3.700 1.125 3.710 1.449 ;
        RECT 3.710 1.125 3.720 1.439 ;
        RECT 3.720 1.125 3.730 1.429 ;
        RECT 3.730 1.125 3.740 1.419 ;
        RECT 3.740 1.125 3.750 1.409 ;
        RECT 3.750 1.125 3.760 1.399 ;
        RECT 3.760 1.125 3.770 1.389 ;
        RECT 3.770 1.125 3.780 1.379 ;
        RECT 3.780 1.125 3.790 1.369 ;
        RECT 3.790 1.125 3.800 1.359 ;
        RECT 3.800 1.125 3.810 1.349 ;
        RECT 3.810 1.125 3.816 1.345 ;
        RECT 3.445 1.415 3.455 2.259 ;
        RECT 3.455 1.405 3.465 2.259 ;
        RECT 3.465 1.395 3.475 2.259 ;
        RECT 3.475 1.385 3.485 2.259 ;
        RECT 3.485 1.375 3.495 2.259 ;
        RECT 3.495 1.365 3.505 2.259 ;
        RECT 3.505 1.355 3.515 2.259 ;
        RECT 3.290 1.570 3.300 1.870 ;
        RECT 3.300 1.560 3.310 1.870 ;
        RECT 3.310 1.550 3.320 1.870 ;
        RECT 3.320 1.540 3.330 1.870 ;
        RECT 3.330 1.530 3.340 1.870 ;
        RECT 3.340 1.520 3.350 1.870 ;
        RECT 3.350 1.510 3.360 1.870 ;
        RECT 3.360 1.500 3.370 1.870 ;
        RECT 3.370 1.490 3.380 1.870 ;
        RECT 3.380 1.480 3.390 1.870 ;
        RECT 3.390 1.470 3.400 1.870 ;
        RECT 3.400 1.460 3.410 1.870 ;
        RECT 3.410 1.450 3.420 1.870 ;
        RECT 3.420 1.440 3.430 1.870 ;
        RECT 3.430 1.430 3.440 1.870 ;
        RECT 3.440 1.420 3.446 1.870 ;
        RECT 1.210 1.125 1.385 2.280 ;
        RECT 1.600 0.775 1.770 1.295 ;
        RECT 1.210 1.125 1.770 1.295 ;
        RECT 2.180 0.645 2.350 0.945 ;
        RECT 4.240 0.640 4.410 0.945 ;
        RECT 1.600 0.775 4.410 0.945 ;
        RECT 3.810 1.610 3.980 1.910 ;
        RECT 3.810 1.610 5.160 1.780 ;
        RECT 4.990 1.060 5.160 2.280 ;
  END 
END RSLATHDLXHT

MACRO RSLATHD2XHT
  CLASS  CORE ;
  FOREIGN RSLATHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.560 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.465 0.510 2.635 2.215 ;
        RECT 2.335 2.045 2.635 2.215 ;
        RECT 2.465 0.510 2.720 1.360 ;
        RECT 2.465 0.510 2.840 0.720 ;
    END
  END Q
  PIN R
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.485 2.900 ;
    END
  END R
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.035 2.470 6.460 2.885 ;
    END
  END S
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.585 1.125 3.885 1.295 ;
        RECT 3.715 1.125 3.770 2.960 ;
        RECT 3.600 1.980 3.770 2.960 ;
        RECT 3.715 1.125 3.885 2.430 ;
        RECT 3.600 1.980 3.885 2.430 ;
        RECT 3.600 2.050 4.000 2.430 ;
    END
  END QN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.235 ;
        RECT 2.030 -0.300 2.200 0.780 ;
        RECT 3.035 -0.300 3.335 0.595 ;
        RECT 4.135 -0.300 4.435 0.595 ;
        RECT 5.600 -0.300 5.900 1.235 ;
        RECT 0.000 -0.300 6.560 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 2.180 0.890 3.990 ;
        RECT 1.765 2.975 2.065 3.990 ;
        RECT 2.855 2.975 3.155 3.990 ;
        RECT 4.205 2.230 4.375 3.990 ;
        RECT 5.515 2.245 5.815 3.990 ;
        RECT 0.000 3.390 6.560 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.605 1.060 1.775 ;
        RECT 0.890 1.540 1.060 1.840 ;
        RECT 1.240 1.125 1.415 2.620 ;
        RECT 1.240 1.125 2.245 1.295 ;
        RECT 2.075 1.125 2.245 1.840 ;
        RECT 1.595 1.520 1.765 2.565 ;
        RECT 3.250 1.510 3.420 2.565 ;
        RECT 1.595 2.395 3.420 2.565 ;
        RECT 3.250 1.510 3.485 1.810 ;
        RECT 4.065 1.510 4.235 1.810 ;
        RECT 4.065 1.575 4.790 1.745 ;
        RECT 4.620 1.125 4.790 2.150 ;
        RECT 4.620 1.980 4.985 2.150 ;
        RECT 4.555 1.125 4.855 1.295 ;
        RECT 4.815 1.980 4.985 2.620 ;
        RECT 2.900 1.110 3.070 1.840 ;
        RECT 2.815 1.540 3.070 1.840 ;
        RECT 3.170 0.775 3.340 1.280 ;
        RECT 2.900 1.110 3.340 1.280 ;
        RECT 3.170 0.775 5.300 0.945 ;
        RECT 5.120 0.775 5.300 1.665 ;
        RECT 5.120 1.495 5.560 1.665 ;
        RECT 4.635 2.890 4.805 3.190 ;
        RECT 5.165 1.845 5.335 3.060 ;
        RECT 4.635 2.890 5.335 3.060 ;
        RECT 5.165 1.845 6.385 2.015 ;
        RECT 6.215 1.060 6.385 2.280 ;
  END 
END RSLATHD2XHT

MACRO RSLATHD1XHT
  CLASS  CORE ;
  FOREIGN RSLATHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.650 0.510 2.125 0.720 ;
        RECT 1.955 0.510 2.125 2.215 ;
        RECT 2.370 2.045 2.540 2.620 ;
        RECT 1.955 2.045 2.605 2.215 ;
    END
  END Q
  PIN R
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.485 2.900 ;
    END
  END R
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.820 2.470 5.230 2.885 ;
    END
  END S
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.880 1.125 3.050 2.620 ;
        RECT 2.880 2.050 3.180 2.620 ;
        RECT 2.880 1.125 3.305 1.295 ;
    END
  END QN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.580 -0.300 0.880 1.295 ;
        RECT 2.440 -0.300 2.740 0.595 ;
        RECT 4.590 -0.300 4.785 1.295 ;
        RECT 4.405 1.125 4.785 1.295 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.095 0.860 3.990 ;
        RECT 1.735 2.910 1.905 3.990 ;
        RECT 3.400 2.570 3.570 3.990 ;
        RECT 4.470 2.100 4.640 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.510 0.340 2.280 ;
        RECT 0.170 1.605 1.030 1.775 ;
        RECT 0.860 1.540 1.030 1.840 ;
        RECT 1.210 1.125 1.385 3.210 ;
        RECT 1.210 3.040 1.555 3.210 ;
        RECT 1.210 1.125 1.770 1.295 ;
        RECT 1.565 1.520 1.735 2.730 ;
        RECT 1.565 2.560 1.980 2.730 ;
        RECT 2.260 3.005 2.835 3.210 ;
        RECT 2.090 2.605 2.100 3.209 ;
        RECT 2.100 2.615 2.110 3.209 ;
        RECT 2.110 2.625 2.120 3.209 ;
        RECT 2.120 2.635 2.130 3.209 ;
        RECT 2.130 2.645 2.140 3.209 ;
        RECT 2.140 2.655 2.150 3.209 ;
        RECT 2.150 2.665 2.160 3.209 ;
        RECT 2.160 2.675 2.170 3.209 ;
        RECT 2.170 2.685 2.180 3.209 ;
        RECT 2.180 2.695 2.190 3.209 ;
        RECT 2.190 2.705 2.200 3.209 ;
        RECT 2.200 2.715 2.210 3.209 ;
        RECT 2.210 2.725 2.220 3.209 ;
        RECT 2.220 2.735 2.230 3.209 ;
        RECT 2.230 2.745 2.240 3.209 ;
        RECT 2.240 2.755 2.250 3.209 ;
        RECT 2.250 2.765 2.260 3.209 ;
        RECT 2.055 2.570 2.065 2.804 ;
        RECT 2.065 2.580 2.075 2.814 ;
        RECT 2.075 2.590 2.085 2.824 ;
        RECT 2.085 2.595 2.091 2.835 ;
        RECT 1.980 2.560 1.990 2.730 ;
        RECT 1.990 2.560 2.000 2.740 ;
        RECT 2.000 2.560 2.010 2.750 ;
        RECT 2.010 2.560 2.020 2.760 ;
        RECT 2.020 2.560 2.030 2.770 ;
        RECT 2.030 2.560 2.040 2.780 ;
        RECT 2.040 2.560 2.050 2.790 ;
        RECT 2.050 2.560 2.056 2.800 ;
        RECT 3.230 1.570 3.290 1.870 ;
        RECT 3.515 1.125 3.630 2.260 ;
        RECT 3.515 2.090 4.185 2.260 ;
        RECT 3.630 1.125 3.640 1.519 ;
        RECT 3.640 1.125 3.650 1.509 ;
        RECT 3.650 1.125 3.660 1.499 ;
        RECT 3.660 1.125 3.670 1.489 ;
        RECT 3.670 1.125 3.680 1.479 ;
        RECT 3.680 1.125 3.690 1.469 ;
        RECT 3.690 1.125 3.700 1.459 ;
        RECT 3.700 1.125 3.710 1.449 ;
        RECT 3.710 1.125 3.720 1.439 ;
        RECT 3.720 1.125 3.730 1.429 ;
        RECT 3.730 1.125 3.740 1.419 ;
        RECT 3.740 1.125 3.750 1.409 ;
        RECT 3.750 1.125 3.760 1.399 ;
        RECT 3.760 1.125 3.770 1.389 ;
        RECT 3.770 1.125 3.780 1.379 ;
        RECT 3.780 1.125 3.790 1.369 ;
        RECT 3.790 1.125 3.800 1.359 ;
        RECT 3.800 1.125 3.810 1.349 ;
        RECT 3.810 1.125 3.816 1.345 ;
        RECT 3.445 1.415 3.455 2.259 ;
        RECT 3.455 1.405 3.465 2.259 ;
        RECT 3.465 1.395 3.475 2.259 ;
        RECT 3.475 1.385 3.485 2.259 ;
        RECT 3.485 1.375 3.495 2.259 ;
        RECT 3.495 1.365 3.505 2.259 ;
        RECT 3.505 1.355 3.515 2.259 ;
        RECT 3.290 1.570 3.300 1.870 ;
        RECT 3.300 1.560 3.310 1.870 ;
        RECT 3.310 1.550 3.320 1.870 ;
        RECT 3.320 1.540 3.330 1.870 ;
        RECT 3.330 1.530 3.340 1.870 ;
        RECT 3.340 1.520 3.350 1.870 ;
        RECT 3.350 1.510 3.360 1.870 ;
        RECT 3.360 1.500 3.370 1.870 ;
        RECT 3.370 1.490 3.380 1.870 ;
        RECT 3.380 1.480 3.390 1.870 ;
        RECT 3.390 1.470 3.400 1.870 ;
        RECT 3.400 1.460 3.410 1.870 ;
        RECT 3.410 1.450 3.420 1.870 ;
        RECT 3.420 1.440 3.430 1.870 ;
        RECT 3.430 1.430 3.440 1.870 ;
        RECT 3.440 1.420 3.446 1.870 ;
        RECT 2.350 0.775 2.520 1.810 ;
        RECT 4.240 0.640 4.410 0.945 ;
        RECT 2.350 0.775 4.410 0.945 ;
        RECT 3.810 1.610 3.980 1.910 ;
        RECT 3.810 1.675 5.160 1.845 ;
        RECT 4.990 1.060 5.160 2.280 ;
  END 
END RSLATHD1XHT

MACRO PULLUHDHT
  CLASS  CORE ;
  FOREIGN PULLUHDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.860 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.295 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.235 1.980 1.540 2.465 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 2.100 0.890 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.205 1.755 ;
  END 
END PULLUHDHT

MACRO OR4HDMXHT
  CLASS  CORE ;
  FOREIGN OR4HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.670 2.560 2.080 3.010 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.220 1.630 1.625 1.950 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 2.710 1.040 3.180 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.380 2.020 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.090 ;
        RECT 1.145 -0.300 1.445 1.090 ;
        RECT 2.215 -0.300 2.515 1.090 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.800 0.850 2.970 2.280 ;
        RECT 2.800 0.850 3.180 1.200 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.280 2.310 2.450 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.585 2.130 0.840 2.370 ;
        RECT 0.105 2.200 0.840 2.370 ;
        RECT 0.690 0.855 0.860 1.450 ;
        RECT 0.690 1.270 2.090 1.450 ;
        RECT 0.585 2.130 2.090 2.305 ;
        RECT 1.760 0.855 1.930 1.450 ;
        RECT 1.920 1.270 2.090 2.305 ;
        RECT 1.920 1.520 2.620 1.820 ;
  END 
END OR4HDMXHT

MACRO OR4HDLXHT
  CLASS  CORE ;
  FOREIGN OR4HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.670 2.560 2.080 3.045 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.220 1.630 1.625 1.950 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 2.710 1.040 3.180 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.400 2.020 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.090 ;
        RECT 1.145 -0.300 1.445 1.090 ;
        RECT 2.215 -0.300 2.515 1.090 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.800 0.850 2.970 2.280 ;
        RECT 2.800 0.850 3.180 1.200 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.280 2.100 2.450 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.585 2.130 0.760 2.370 ;
        RECT 0.105 2.200 0.760 2.370 ;
        RECT 0.690 0.855 0.860 1.450 ;
        RECT 0.690 1.270 2.090 1.450 ;
        RECT 0.585 2.130 2.090 2.305 ;
        RECT 1.760 0.855 1.930 1.450 ;
        RECT 1.920 1.270 2.090 2.305 ;
        RECT 1.920 1.520 2.620 1.820 ;
  END 
END OR4HDLXHT

MACRO OR4HD2XHT
  CLASS  CORE ;
  FOREIGN OR4HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.630 2.145 2.020 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 1.610 1.540 2.430 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.675 0.720 2.020 ;
        RECT 0.510 1.675 1.105 1.845 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.260 0.330 1.820 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.070 ;
        RECT 1.145 -0.300 1.445 1.070 ;
        RECT 2.215 -0.300 2.515 1.070 ;
        RECT 3.255 -0.300 3.555 1.055 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.800 0.720 2.970 2.960 ;
        RECT 2.800 1.260 3.180 1.610 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.280 2.570 2.450 3.990 ;
        RECT 3.255 2.295 3.555 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.185 0.405 3.035 ;
        RECT 0.690 1.025 0.860 1.430 ;
        RECT 1.760 1.025 1.930 1.430 ;
        RECT 1.870 2.200 2.050 2.780 ;
        RECT 0.105 2.610 2.050 2.780 ;
        RECT 0.690 1.260 2.620 1.430 ;
        RECT 2.450 1.260 2.620 2.380 ;
        RECT 1.870 2.200 2.620 2.380 ;
  END 
END OR4HD2XHT

MACRO OR4HD1XHT
  CLASS  CORE ;
  FOREIGN OR4HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.585 1.610 2.110 1.950 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.260 2.560 1.625 3.080 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 2.800 1.040 3.180 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.380 2.020 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.090 ;
        RECT 1.145 -0.300 1.445 1.080 ;
        RECT 2.215 -0.300 2.515 1.080 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.800 0.720 2.970 2.960 ;
        RECT 2.800 0.850 3.180 1.200 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.215 2.635 2.515 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 0.845 0.860 1.430 ;
        RECT 1.760 0.845 1.930 1.430 ;
        RECT 0.690 1.260 2.620 1.430 ;
        RECT 2.450 1.260 2.620 2.370 ;
        RECT 0.105 2.200 2.620 2.370 ;
  END 
END OR4HD1XHT

MACRO OR3HDLXHT
  CLASS  CORE ;
  FOREIGN OR3HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.850 2.710 1.400 3.180 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.530 0.720 2.020 ;
        RECT 0.510 1.530 1.070 1.755 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.255 0.330 1.820 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.555 -0.300 0.855 1.295 ;
        RECT 1.505 -0.300 1.805 0.715 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.120 1.060 2.360 1.360 ;
        RECT 2.170 1.060 2.360 2.840 ;
        RECT 2.120 2.100 2.360 2.840 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.600 2.100 1.770 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.060 0.510 1.230 1.295 ;
        RECT 1.060 1.125 1.420 1.295 ;
        RECT 1.250 1.125 1.420 2.370 ;
        RECT 0.105 2.200 1.420 2.370 ;
        RECT 1.250 1.610 1.990 1.910 ;
  END 
END OR3HDLXHT

MACRO OR3HD2XHT
  CLASS  CORE ;
  FOREIGN OR3HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.245 1.615 1.730 1.995 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.610 0.720 2.430 ;
        RECT 0.510 1.610 1.000 1.910 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.090 1.610 0.330 2.160 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.000 ;
        RECT 1.695 -0.300 1.995 1.055 ;
        RECT 2.735 -0.300 3.035 1.055 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.280 0.720 2.450 3.075 ;
        RECT 2.280 1.330 2.840 1.540 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.665 2.635 1.965 3.990 ;
        RECT 2.735 2.295 3.035 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.025 0.345 1.405 ;
        RECT 0.105 2.610 0.405 3.145 ;
        RECT 1.075 2.220 1.245 2.780 ;
        RECT 0.105 2.610 1.245 2.780 ;
        RECT 1.145 1.090 1.445 1.405 ;
        RECT 0.170 1.180 1.445 1.405 ;
        RECT 0.170 1.235 2.080 1.405 ;
        RECT 1.910 1.235 2.080 2.390 ;
        RECT 1.075 2.220 2.080 2.390 ;
  END 
END OR3HD2XHT

MACRO OR3HD1XHT
  CLASS  CORE ;
  FOREIGN OR3HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.850 2.910 1.400 3.210 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.530 0.720 2.020 ;
        RECT 0.510 1.530 1.070 1.755 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.260 0.325 1.820 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 1.295 ;
        RECT 1.535 -0.300 1.835 0.715 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.120 0.720 2.360 1.405 ;
        RECT 2.170 0.720 2.360 3.010 ;
        RECT 2.055 2.095 2.360 3.010 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.600 2.230 1.770 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.055 0.510 1.225 1.295 ;
        RECT 1.055 1.125 1.420 1.295 ;
        RECT 1.250 1.125 1.420 2.370 ;
        RECT 0.105 2.200 1.420 2.370 ;
        RECT 1.250 1.610 1.990 1.910 ;
  END 
END OR3HD1XHT

MACRO OR2ODHDHT
  CLASS  CORE ;
  FOREIGN OR2ODHDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 1.585 1.130 2.020 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.510 2.020 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.195 ;
        RECT 1.175 -0.300 1.475 1.055 ;
        RECT 2.215 -0.300 2.515 1.055 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 1.760 0.720 1.930 1.415 ;
        RECT 2.090 1.235 2.420 1.540 ;
        RECT 2.800 0.720 2.970 1.415 ;
        RECT 1.760 1.235 2.970 1.415 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.175 2.550 1.475 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 1.060 0.860 1.405 ;
        RECT 0.690 1.235 1.475 1.405 ;
        RECT 1.310 1.270 1.480 2.370 ;
        RECT 0.105 2.200 1.480 2.370 ;
        RECT 1.310 1.720 2.495 1.890 ;
  END 
END OR2ODHDHT

MACRO OR2HDUXHT
  CLASS  CORE ;
  FOREIGN OR2HDUXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.090 1.705 0.495 2.490 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.675 1.270 1.130 1.835 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.215 -0.300 0.515 0.510 ;
        RECT 0.775 -0.300 1.075 0.660 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.255 0.480 1.830 0.735 ;
        RECT 1.660 0.480 1.830 2.900 ;
        RECT 1.105 2.600 1.830 2.900 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.145 2.795 0.445 3.990 ;
        RECT 1.060 3.180 1.380 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.710 2.155 0.880 3.210 ;
        RECT 0.315 0.915 1.480 1.090 ;
        RECT 1.310 0.915 1.480 2.325 ;
        RECT 0.710 2.155 1.480 2.325 ;
  END 
END OR2HDUXHT

MACRO OR2HDMXHT
  CLASS  CORE ;
  FOREIGN OR2HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.375 2.910 0.890 3.210 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.510 2.020 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.295 ;
        RECT 1.055 -0.300 1.355 0.720 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.605 1.125 1.950 1.295 ;
        RECT 1.740 1.125 1.950 2.215 ;
        RECT 1.545 1.980 1.950 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.090 2.310 1.260 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 1.060 0.860 2.370 ;
        RECT 0.105 2.200 0.860 2.370 ;
        RECT 0.690 1.495 1.520 1.795 ;
  END 
END OR2HDMXHT

MACRO OR2HDLXHT
  CLASS  CORE ;
  FOREIGN OR2HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 2.870 0.890 3.210 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.510 2.020 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.295 ;
        RECT 1.145 -0.300 1.445 0.745 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.710 1.060 1.950 1.360 ;
        RECT 1.740 1.060 1.950 2.215 ;
        RECT 1.545 2.045 1.950 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.090 2.100 1.260 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 1.060 0.860 2.370 ;
        RECT 0.105 2.200 0.860 2.370 ;
        RECT 0.690 1.495 1.540 1.795 ;
  END 
END OR2HDLXHT

MACRO OR2HD2XHT
  CLASS  CORE ;
  FOREIGN OR2HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.815 1.590 1.130 2.020 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.260 0.310 1.820 ;
        RECT 0.100 1.520 0.510 1.820 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 0.995 ;
        RECT 1.175 -0.300 1.475 1.055 ;
        RECT 2.215 -0.300 2.515 1.055 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.760 1.945 1.930 2.960 ;
        RECT 1.740 0.720 1.950 1.415 ;
        RECT 1.740 1.235 2.165 1.415 ;
        RECT 1.995 1.235 2.165 2.115 ;
        RECT 1.760 1.945 2.165 2.115 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.175 2.635 1.475 3.990 ;
        RECT 2.215 2.295 2.515 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.200 0.405 3.055 ;
        RECT 0.690 1.060 0.860 1.405 ;
        RECT 0.690 1.235 1.475 1.405 ;
        RECT 1.310 1.270 1.480 2.370 ;
        RECT 0.105 2.200 1.480 2.370 ;
        RECT 1.310 1.595 1.815 1.765 ;
  END 
END OR2HD2XHT

MACRO OR2HD2XSPGHT
  CLASS  CORE ;
  FOREIGN OR2HD2XSPGHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 2.805 0.425 3.345 3.070 ;
      LAYER V7 ;
        RECT 2.895 2.485 3.255 2.845 ;
      LAYER M7 ;
        RECT 0.405 2.475 3.345 2.855 ;
      LAYER V6 ;
        RECT 2.980 2.570 3.170 2.760 ;
      LAYER M4 ;
        RECT 0.515 1.925 0.715 2.945 ;
      LAYER V3 ;
        RECT 0.520 2.160 0.710 2.350 ;
      LAYER M3 ;
        RECT 0.385 2.155 1.635 2.355 ;
      LAYER V2 ;
        RECT 1.340 2.160 1.530 2.350 ;
      LAYER M2 ;
        RECT 1.335 1.540 1.535 2.460 ;
      LAYER V1 ;
        RECT 1.340 1.750 1.530 1.940 ;
      LAYER M1 ;
        RECT 1.330 1.590 1.675 2.020 ;
      LAYER M6 ;
        RECT 2.975 0.750 3.175 3.070 ;
      LAYER V5 ;
        RECT 2.980 2.570 3.170 2.760 ;
      LAYER M5 ;
        RECT 0.405 2.565 3.345 2.765 ;
      LAYER V4 ;
        RECT 0.520 2.570 0.710 2.760 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 0.345 0.425 0.885 3.085 ;
      LAYER V7 ;
        RECT 0.435 0.845 0.795 1.205 ;
      LAYER M7 ;
        RECT 0.310 0.835 1.105 1.215 ;
      LAYER V6 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M4 ;
        RECT 0.515 0.760 0.715 1.490 ;
      LAYER V3 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M3 ;
        RECT 0.105 0.860 0.835 1.190 ;
      LAYER V2 ;
        RECT 0.110 0.930 0.300 1.120 ;
      LAYER M2 ;
        RECT 0.105 0.860 0.305 1.920 ;
      LAYER V1 ;
        RECT 0.110 1.575 0.300 1.765 ;
      LAYER M1 ;
        RECT 0.100 1.260 0.310 1.840 ;
        RECT 0.100 1.520 1.055 1.840 ;
      LAYER M6 ;
        RECT 0.515 0.425 0.715 1.690 ;
      LAYER V5 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M5 ;
        RECT 0.310 0.925 1.105 1.125 ;
      LAYER V4 ;
        RECT 0.520 0.930 0.710 1.120 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.650 -0.300 0.950 0.995 ;
        RECT 1.720 -0.300 2.020 1.055 ;
        RECT 2.760 -0.300 3.060 0.780 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 1.575 0.425 2.115 3.070 ;
      LAYER V7 ;
        RECT 1.665 0.845 2.025 1.205 ;
      LAYER M7 ;
        RECT 1.510 0.835 2.525 1.215 ;
      LAYER V6 ;
        RECT 1.750 0.930 1.940 1.120 ;
      LAYER M4 ;
        RECT 2.155 0.790 2.355 1.670 ;
      LAYER V3 ;
        RECT 2.160 1.340 2.350 1.530 ;
      LAYER M3 ;
        RECT 1.975 1.335 2.905 1.535 ;
      LAYER V2 ;
        RECT 2.570 1.340 2.760 1.530 ;
      LAYER M2 ;
        RECT 2.565 1.230 2.765 2.050 ;
      LAYER V1 ;
        RECT 2.570 1.750 2.760 1.940 ;
      LAYER M1 ;
        RECT 2.280 0.480 2.490 1.330 ;
        RECT 2.240 2.045 2.540 2.960 ;
        RECT 2.280 1.120 2.770 1.330 ;
        RECT 2.560 1.120 2.770 2.260 ;
        RECT 2.240 2.045 2.770 2.260 ;
      LAYER M6 ;
        RECT 1.745 0.425 1.945 1.690 ;
      LAYER V5 ;
        RECT 1.750 0.930 1.940 1.120 ;
      LAYER M5 ;
        RECT 1.510 0.925 2.525 1.125 ;
      LAYER V4 ;
        RECT 2.160 0.930 2.350 1.120 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.720 2.635 2.020 3.990 ;
        RECT 2.760 2.475 3.060 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.650 2.200 0.950 3.055 ;
        RECT 1.235 1.060 1.405 1.405 ;
        RECT 1.235 1.235 2.020 1.405 ;
        RECT 1.855 1.270 2.025 2.370 ;
        RECT 0.650 2.200 2.025 2.370 ;
        RECT 1.855 1.530 2.360 1.830 ;
  END 
END OR2HD2XSPGHT

MACRO OAI22B2HD1XHT
  CLASS  CORE ;
  FOREIGN OAI22B2HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.650 1.300 2.015 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.480 1.650 1.780 2.360 ;
        RECT 1.480 2.150 2.010 2.360 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.000 1.675 2.500 1.950 ;
    END
  END D
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.570 0.390 2.010 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.140 -0.300 1.440 1.055 ;
        RECT 2.180 -0.300 2.480 0.715 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.405 2.130 2.575 3.045 ;
        RECT 3.325 0.720 3.495 2.300 ;
        RECT 2.340 2.130 3.495 2.300 ;
        RECT 3.325 1.220 3.590 1.635 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.195 2.190 0.365 3.990 ;
        RECT 1.230 2.635 1.530 3.990 ;
        RECT 2.890 2.635 3.530 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.130 1.050 0.740 1.220 ;
        RECT 0.570 1.050 0.740 2.365 ;
        RECT 0.570 2.195 0.950 2.365 ;
        RECT 0.570 1.300 2.945 1.470 ;
        RECT 2.775 1.300 2.945 1.920 ;
        RECT 1.725 0.480 1.895 1.120 ;
        RECT 2.805 0.480 2.975 1.120 ;
        RECT 1.725 0.950 2.975 1.120 ;
  END 
END OAI22B2HD1XHT

MACRO OAI222HDLXHT
  CLASS  CORE ;
  FOREIGN OAI222HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.635 0.310 2.015 ;
        RECT 0.100 1.635 0.615 1.870 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.860 1.805 1.030 2.360 ;
        RECT 0.445 2.150 1.030 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.875 1.650 2.175 1.950 ;
        RECT 1.875 1.740 2.425 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.215 1.635 1.625 1.950 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.560 1.220 2.790 1.620 ;
        RECT 2.605 1.220 2.790 1.800 ;
    END
  END E
  PIN F
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.970 1.245 3.185 1.950 ;
        RECT 2.970 1.245 3.230 1.865 ;
    END
  END F
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 -0.300 0.895 0.745 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.735 0.895 3.590 1.040 ;
        RECT 1.210 2.130 1.380 2.605 ;
        RECT 2.895 0.870 3.065 1.065 ;
        RECT 2.735 0.870 3.065 1.040 ;
        RECT 1.210 2.130 3.590 2.300 ;
        RECT 2.895 0.895 3.590 1.065 ;
        RECT 3.380 2.065 3.490 2.715 ;
        RECT 3.380 2.065 3.590 2.450 ;
        RECT 3.410 0.895 3.490 2.715 ;
        RECT 3.320 2.130 3.490 2.715 ;
        RECT 3.410 0.895 3.590 2.450 ;
        RECT 3.320 2.130 3.590 2.450 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.540 0.405 3.990 ;
        RECT 2.215 2.480 2.515 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 1.455 ;
        RECT 1.210 1.060 1.380 1.455 ;
        RECT 2.210 1.060 2.380 1.455 ;
        RECT 0.170 1.285 2.380 1.455 ;
        RECT 2.250 0.520 2.485 0.715 ;
        RECT 1.695 0.545 2.485 0.715 ;
        RECT 3.285 0.520 3.455 0.715 ;
        RECT 2.250 0.520 3.455 0.690 ;
        RECT 3.285 0.545 3.585 0.715 ;
  END 
END OAI222HDLXHT

MACRO OAI222HD2XHT
  CLASS  CORE ;
  FOREIGN OAI222HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.740 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.645 0.310 2.015 ;
        RECT 0.100 1.645 0.615 1.815 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.795 2.545 1.375 2.830 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.875 1.635 2.175 1.950 ;
        RECT 1.875 1.740 2.425 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.215 1.635 1.655 1.950 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.560 1.220 2.790 1.620 ;
        RECT 2.605 1.220 2.790 1.800 ;
    END
  END E
  PIN F
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.320 0.920 3.810 1.260 ;
    END
  END F
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.570 -0.300 0.870 0.745 ;
        RECT 4.360 -0.300 4.530 0.780 ;
        RECT 5.335 -0.300 5.635 1.055 ;
        RECT 0.000 -0.300 5.740 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.880 0.720 5.050 2.960 ;
        RECT 4.880 1.235 5.230 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.195 0.405 3.990 ;
        RECT 2.215 2.480 2.515 3.990 ;
        RECT 4.295 2.295 4.595 3.990 ;
        RECT 5.335 2.295 5.635 3.990 ;
        RECT 0.000 3.390 5.740 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 1.455 ;
        RECT 1.185 1.060 1.355 1.455 ;
        RECT 2.200 1.060 2.370 1.455 ;
        RECT 0.170 1.285 2.370 1.455 ;
        RECT 2.230 0.520 2.465 0.715 ;
        RECT 1.670 0.545 2.465 0.715 ;
        RECT 3.265 0.520 3.435 0.715 ;
        RECT 2.230 0.520 3.435 0.690 ;
        RECT 3.265 0.545 3.565 0.715 ;
        RECT 2.890 0.870 3.060 1.065 ;
        RECT 2.890 0.895 3.140 1.065 ;
        RECT 2.715 0.870 3.060 1.040 ;
        RECT 2.970 0.895 3.140 2.300 ;
        RECT 1.145 2.130 3.535 2.300 ;
        RECT 2.970 1.595 4.255 1.765 ;
        RECT 3.810 1.945 3.980 2.280 ;
        RECT 3.775 0.545 4.160 0.715 ;
        RECT 3.990 0.545 4.160 1.130 ;
        RECT 3.990 0.960 4.670 1.130 ;
        RECT 4.500 0.960 4.670 2.115 ;
        RECT 3.810 1.945 4.670 2.115 ;
  END 
END OAI222HD2XHT

MACRO OAI222HD1XHT
  CLASS  CORE ;
  FOREIGN OAI222HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.630 0.310 2.015 ;
        RECT 0.100 1.630 0.585 1.845 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.830 1.610 1.000 2.360 ;
        RECT 0.445 2.150 1.000 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.835 1.635 2.430 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.215 1.635 1.655 1.950 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.650 1.450 2.820 1.880 ;
        RECT 2.650 1.710 3.180 1.880 ;
        RECT 2.970 1.710 3.180 2.420 ;
    END
  END E
  PIN F
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.715 1.250 4.000 1.910 ;
    END
  END F
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.055 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.345 1.320 3.530 1.490 ;
        RECT 1.210 2.200 1.380 3.180 ;
        RECT 0.860 2.970 1.380 3.180 ;
        RECT 1.210 2.200 2.790 2.370 ;
        RECT 2.620 2.200 2.790 2.960 ;
        RECT 3.175 1.005 3.515 1.175 ;
        RECT 3.360 1.005 3.515 2.960 ;
        RECT 3.345 1.005 3.515 1.490 ;
        RECT 3.360 1.320 3.530 2.960 ;
        RECT 2.620 2.790 3.530 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.635 0.405 3.990 ;
        RECT 2.140 2.635 2.440 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.690 0.340 1.430 ;
        RECT 1.210 0.690 1.380 1.430 ;
        RECT 2.250 1.030 2.420 1.430 ;
        RECT 0.170 1.260 2.420 1.430 ;
        RECT 1.665 0.545 1.965 1.055 ;
        RECT 1.665 0.545 3.995 0.715 ;
        RECT 3.695 0.545 3.995 1.055 ;
  END 
END OAI222HD1XHT

MACRO OAI221HDMXHT
  CLASS  CORE ;
  FOREIGN OAI221HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.640 0.310 2.015 ;
        RECT 0.100 1.640 0.585 1.810 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.830 1.575 1.000 2.360 ;
        RECT 0.445 2.150 1.000 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.835 1.630 2.430 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.215 1.575 1.610 1.950 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.785 1.330 3.240 1.865 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.045 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.210 2.130 1.380 2.775 ;
        RECT 3.105 2.060 3.590 2.300 ;
        RECT 1.210 2.130 3.590 2.300 ;
        RECT 3.245 0.875 3.590 1.045 ;
        RECT 3.380 2.030 3.590 2.430 ;
        RECT 3.420 0.875 3.590 2.430 ;
        RECT 3.375 2.060 3.590 2.430 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.540 0.405 3.990 ;
        RECT 2.215 2.540 2.855 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 1.395 ;
        RECT 1.210 1.060 1.380 1.395 ;
        RECT 2.280 1.060 2.450 1.395 ;
        RECT 0.170 1.225 2.450 1.395 ;
        RECT 1.910 0.710 2.080 1.045 ;
        RECT 1.695 0.875 2.080 1.045 ;
        RECT 2.725 0.710 2.895 1.045 ;
        RECT 1.910 0.710 2.895 0.880 ;
        RECT 2.725 0.875 3.025 1.045 ;
  END 
END OAI221HDMXHT

MACRO OAI221HDLXHT
  CLASS  CORE ;
  FOREIGN OAI221HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.640 0.310 2.015 ;
        RECT 0.100 1.640 0.585 1.810 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.815 2.665 1.215 3.180 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.835 1.630 2.430 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.215 1.575 1.610 1.950 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.790 1.265 3.180 1.815 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.045 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.310 0.810 3.530 1.110 ;
        RECT 3.105 2.045 3.590 2.300 ;
        RECT 1.145 2.130 3.590 2.300 ;
        RECT 3.380 0.810 3.530 2.455 ;
        RECT 3.360 0.810 3.530 2.300 ;
        RECT 3.380 2.045 3.590 2.455 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 2.215 2.480 2.855 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.900 0.340 1.395 ;
        RECT 1.210 0.900 1.380 1.395 ;
        RECT 2.280 0.900 2.450 1.395 ;
        RECT 0.170 1.225 2.450 1.395 ;
        RECT 1.910 0.550 2.080 1.045 ;
        RECT 1.695 0.875 2.080 1.045 ;
        RECT 1.910 0.550 2.895 0.720 ;
        RECT 2.725 0.550 2.895 1.045 ;
        RECT 2.725 0.875 3.025 1.045 ;
  END 
END OAI221HDLXHT

MACRO OR2HD1XHT
  CLASS  CORE ;
  FOREIGN OR2HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 2.910 0.890 3.210 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.510 2.020 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.295 ;
        RECT 1.085 -0.300 1.385 0.720 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.670 1.190 1.950 1.360 ;
        RECT 1.700 0.720 1.840 2.895 ;
        RECT 1.670 0.720 1.840 1.360 ;
        RECT 1.700 1.190 1.870 2.895 ;
        RECT 1.545 1.980 1.870 2.895 ;
        RECT 1.700 1.190 1.950 1.650 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.090 2.230 1.260 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 1.060 0.860 2.370 ;
        RECT 0.105 2.200 0.860 2.370 ;
        RECT 0.690 1.495 1.520 1.795 ;
  END 
END OR2HD1XHT

MACRO OAI21B2HD1XHT
  CLASS  CORE ;
  FOREIGN OAI21B2HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.270 1.150 2.055 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 1.530 1.605 2.020 ;
    END
  END C
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.570 0.390 2.020 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.200 -0.300 1.500 0.715 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.785 2.060 2.020 3.040 ;
        RECT 1.740 2.490 2.020 3.040 ;
        RECT 2.305 0.720 2.475 2.230 ;
        RECT 1.785 2.060 2.475 2.230 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.195 2.200 0.365 3.990 ;
        RECT 1.200 2.465 1.500 3.990 ;
        RECT 2.240 2.465 2.540 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.130 1.050 0.740 1.220 ;
        RECT 0.570 0.920 0.740 2.435 ;
        RECT 0.570 2.265 0.950 2.435 ;
        RECT 0.570 0.920 2.125 1.090 ;
        RECT 1.955 0.920 2.125 1.865 ;
  END 
END OAI21B2HD1XHT

MACRO OAI211HDMXHT
  CLASS  CORE ;
  FOREIGN OAI211HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.575 0.310 2.015 ;
        RECT 0.100 1.575 0.570 1.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.880 1.575 1.050 2.360 ;
        RECT 0.445 2.150 1.050 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.265 1.575 1.655 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.560 1.265 2.770 1.865 ;
        RECT 2.185 1.565 2.770 1.865 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.675 -0.300 0.975 1.045 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.260 2.130 1.430 2.775 ;
        RECT 1.740 0.855 2.005 1.210 ;
        RECT 1.835 0.855 2.005 2.300 ;
        RECT 1.260 2.130 2.500 2.300 ;
        RECT 2.330 2.130 2.500 2.645 ;
        RECT 1.740 0.855 2.565 1.045 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.540 0.455 3.990 ;
        RECT 1.745 2.540 2.045 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.220 1.060 0.390 1.395 ;
        RECT 1.260 1.060 1.430 1.395 ;
        RECT 0.220 1.225 1.430 1.395 ;
  END 
END OAI211HDMXHT

MACRO OAI211HDLXHT
  CLASS  CORE ;
  FOREIGN OAI211HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.575 0.310 2.015 ;
        RECT 0.100 1.575 0.570 1.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.880 1.575 1.050 2.360 ;
        RECT 0.445 2.150 1.050 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.265 1.575 1.655 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.185 1.265 2.770 1.800 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.675 -0.300 0.975 1.045 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.260 2.130 1.430 2.525 ;
        RECT 1.740 0.855 2.005 1.200 ;
        RECT 1.835 0.855 2.005 2.300 ;
        RECT 1.260 2.130 2.500 2.300 ;
        RECT 2.330 2.130 2.500 2.775 ;
        RECT 1.740 0.855 2.565 1.045 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.540 0.455 3.990 ;
        RECT 1.745 2.540 2.045 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.220 0.900 0.390 1.395 ;
        RECT 1.260 0.900 1.430 1.395 ;
        RECT 0.220 1.225 1.430 1.395 ;
  END 
END OAI211HDLXHT

MACRO OR2HD1XSPGHT
  CLASS  CORE ;
  FOREIGN OR2HD1XSPGHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 2.805 0.425 3.345 3.380 ;
      LAYER V7 ;
        RECT 2.895 2.895 3.255 3.255 ;
      LAYER M7 ;
        RECT 1.305 2.885 3.345 3.265 ;
      LAYER V6 ;
        RECT 2.980 2.980 3.170 3.170 ;
      LAYER M4 ;
        RECT 1.745 2.375 1.945 3.290 ;
      LAYER V3 ;
        RECT 1.750 2.565 1.940 2.755 ;
      LAYER M3 ;
        RECT 1.190 2.560 2.075 2.760 ;
      LAYER V2 ;
        RECT 1.340 2.565 1.530 2.755 ;
      LAYER M2 ;
        RECT 1.335 2.405 1.535 3.300 ;
      LAYER V1 ;
        RECT 1.340 2.980 1.530 3.170 ;
      LAYER M1 ;
        RECT 1.200 2.865 1.720 3.210 ;
      LAYER M6 ;
        RECT 2.975 0.830 3.175 3.340 ;
      LAYER V5 ;
        RECT 2.980 2.980 3.170 3.170 ;
      LAYER M5 ;
        RECT 1.575 2.975 3.345 3.175 ;
      LAYER V4 ;
        RECT 1.750 2.980 1.940 3.170 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 0.345 0.425 0.885 3.075 ;
      LAYER V7 ;
        RECT 0.435 1.665 0.795 2.025 ;
      LAYER M7 ;
        RECT 0.205 1.595 0.885 2.095 ;
      LAYER V6 ;
        RECT 0.520 1.750 0.710 1.940 ;
      LAYER M4 ;
        RECT 0.515 1.180 0.715 2.095 ;
      LAYER V3 ;
        RECT 0.520 1.340 0.710 1.530 ;
      LAYER M3 ;
        RECT 0.105 1.265 0.750 1.605 ;
      LAYER V2 ;
        RECT 0.110 1.340 0.300 1.530 ;
      LAYER M2 ;
        RECT 0.105 1.165 0.305 2.060 ;
      LAYER V1 ;
        RECT 0.110 1.750 0.300 1.940 ;
      LAYER M1 ;
        RECT 0.100 1.520 0.310 2.020 ;
        RECT 0.100 1.520 1.340 1.820 ;
      LAYER M6 ;
        RECT 0.515 0.830 0.715 2.495 ;
      LAYER V5 ;
        RECT 0.520 1.750 0.710 1.940 ;
      LAYER M5 ;
        RECT 0.205 1.745 1.265 1.945 ;
      LAYER V4 ;
        RECT 0.520 1.750 0.710 1.940 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.935 -0.300 1.235 1.295 ;
        RECT 1.915 -0.300 2.215 0.720 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 1.575 0.425 2.115 3.075 ;
      LAYER V7 ;
        RECT 1.665 1.255 2.025 1.615 ;
      LAYER M7 ;
        RECT 1.205 1.185 2.115 1.685 ;
      LAYER V6 ;
        RECT 1.750 1.340 1.940 1.530 ;
      LAYER M4 ;
        RECT 1.335 0.720 1.535 1.675 ;
      LAYER V3 ;
        RECT 1.340 0.930 1.530 1.120 ;
      LAYER M3 ;
        RECT 1.205 0.925 2.925 1.125 ;
      LAYER V2 ;
        RECT 2.570 0.930 2.760 1.120 ;
      LAYER M2 ;
        RECT 2.565 0.845 2.765 1.670 ;
      LAYER V1 ;
        RECT 2.570 1.340 2.760 1.530 ;
      LAYER M1 ;
        RECT 2.500 1.190 2.780 1.360 ;
        RECT 2.530 0.720 2.670 2.960 ;
        RECT 2.500 0.720 2.670 1.360 ;
        RECT 2.530 1.190 2.780 2.960 ;
        RECT 2.375 1.980 2.780 2.960 ;
      LAYER M6 ;
        RECT 1.745 0.830 1.945 2.495 ;
      LAYER V5 ;
        RECT 1.750 1.340 1.940 1.530 ;
      LAYER M5 ;
        RECT 1.060 1.335 2.435 1.535 ;
      LAYER V4 ;
        RECT 1.340 1.340 1.530 1.530 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.920 2.230 2.090 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.520 1.060 1.690 2.370 ;
        RECT 0.935 2.200 1.690 2.370 ;
        RECT 1.520 1.495 2.350 1.795 ;
  END 
END OR2HD1XSPGHT

MACRO OAI33HDMXHT
  CLASS  CORE ;
  FOREIGN OAI33HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.270 0.325 1.880 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.505 1.595 0.720 2.020 ;
        RECT 0.505 1.595 1.040 1.895 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.350 1.595 1.520 2.360 ;
        RECT 0.860 2.150 1.520 2.360 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.625 1.950 2.030 ;
        RECT 1.740 1.625 2.245 1.795 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.460 1.610 2.630 2.360 ;
        RECT 2.090 2.150 2.630 2.360 ;
    END
  END E
  PIN F
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.880 1.595 3.180 2.020 ;
    END
  END F
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.065 ;
        RECT 1.145 -0.300 1.445 1.065 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.700 2.230 1.870 3.210 ;
        RECT 2.250 0.920 2.420 1.415 ;
        RECT 2.875 2.200 3.045 2.770 ;
        RECT 1.700 2.560 3.045 2.770 ;
        RECT 3.290 0.920 3.530 1.415 ;
        RECT 2.250 1.245 3.530 1.415 ;
        RECT 3.360 0.920 3.530 2.370 ;
        RECT 2.875 2.200 3.530 2.370 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 3.225 2.635 3.525 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 0.920 0.860 1.415 ;
        RECT 1.730 0.570 1.900 1.415 ;
        RECT 0.690 1.245 1.900 1.415 ;
        RECT 1.730 0.570 3.005 0.740 ;
        RECT 2.705 0.570 3.005 1.065 ;
  END 
END OAI33HDMXHT

MACRO OAI33HDLXHT
  CLASS  CORE ;
  FOREIGN OAI33HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.270 0.330 2.115 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.595 1.040 2.020 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.350 1.685 1.520 2.770 ;
        RECT 0.860 2.560 1.520 2.770 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.610 1.950 2.030 ;
        RECT 1.740 1.610 2.105 1.910 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.430 1.610 2.600 2.360 ;
        RECT 2.090 2.150 2.600 2.360 ;
    END
  END E
  PIN F
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.880 1.595 3.180 2.020 ;
    END
  END F
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.065 ;
        RECT 1.145 -0.300 1.445 1.065 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.700 2.485 1.870 3.125 ;
        RECT 2.185 0.895 2.485 1.065 ;
        RECT 2.315 0.895 2.485 1.415 ;
        RECT 2.875 2.200 3.045 2.770 ;
        RECT 1.700 2.560 3.045 2.770 ;
        RECT 3.290 0.830 3.530 1.415 ;
        RECT 2.315 1.245 3.530 1.415 ;
        RECT 3.360 0.830 3.530 2.370 ;
        RECT 2.875 2.200 3.530 2.370 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.550 0.405 3.990 ;
        RECT 3.225 2.550 3.525 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 0.830 0.860 1.415 ;
        RECT 1.730 0.520 1.900 1.415 ;
        RECT 0.690 1.245 1.900 1.415 ;
        RECT 1.730 0.520 3.005 0.690 ;
        RECT 2.705 0.520 3.005 1.065 ;
  END 
END OAI33HDLXHT

MACRO OAI33HD2XHT
  CLASS  CORE ;
  FOREIGN OAI33HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.740 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.270 0.310 1.810 ;
        RECT 0.100 1.640 0.585 1.810 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.870 1.595 1.040 2.360 ;
        RECT 0.450 2.150 1.040 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.350 1.685 1.520 2.770 ;
        RECT 0.860 2.560 1.520 2.770 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.700 1.610 2.040 2.010 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.570 1.610 2.740 2.770 ;
        RECT 2.500 2.560 2.830 2.770 ;
    END
  END E
  PIN F
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.950 1.595 3.250 2.020 ;
    END
  END F
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.065 ;
        RECT 1.145 -0.300 1.445 1.065 ;
        RECT 4.285 -0.300 4.585 1.055 ;
        RECT 5.325 -0.300 5.625 1.055 ;
        RECT 0.000 -0.300 5.740 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.870 0.720 5.040 2.960 ;
        RECT 4.870 1.235 5.230 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.550 0.405 3.990 ;
        RECT 3.225 2.550 3.525 3.990 ;
        RECT 4.285 2.635 4.585 3.990 ;
        RECT 5.325 2.295 5.625 3.990 ;
        RECT 0.000 3.390 5.740 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 0.830 0.860 1.415 ;
        RECT 1.730 0.520 1.900 1.415 ;
        RECT 0.690 1.245 1.900 1.415 ;
        RECT 1.730 0.520 3.005 0.690 ;
        RECT 2.705 0.520 3.005 1.065 ;
        RECT 1.700 2.200 1.870 2.840 ;
        RECT 2.220 0.895 2.390 2.370 ;
        RECT 1.700 2.200 2.390 2.370 ;
        RECT 2.220 0.895 2.420 1.415 ;
        RECT 2.185 0.895 2.485 1.065 ;
        RECT 2.220 1.245 3.630 1.415 ;
        RECT 3.290 0.830 3.460 1.415 ;
        RECT 3.460 1.245 3.630 1.835 ;
        RECT 3.460 1.630 4.215 1.835 ;
        RECT 3.735 0.860 4.075 1.030 ;
        RECT 3.905 0.860 4.075 1.445 ;
        RECT 3.905 1.275 4.690 1.445 ;
        RECT 4.520 1.275 4.690 2.215 ;
        RECT 3.735 2.045 4.690 2.215 ;
  END 
END OAI33HD2XHT

MACRO OAI33HD1XHT
  CLASS  CORE ;
  FOREIGN OAI33HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.090 1.270 0.325 1.880 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.505 1.660 0.800 2.020 ;
        RECT 0.505 1.660 1.105 1.830 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.285 1.685 1.520 2.770 ;
        RECT 0.860 2.560 1.520 2.770 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.720 1.610 1.950 2.010 ;
        RECT 1.720 1.610 2.110 1.910 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.430 1.610 2.600 2.360 ;
        RECT 2.090 2.150 2.600 2.360 ;
    END
  END E
  PIN F
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.885 1.595 3.250 1.950 ;
    END
  END F
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.065 ;
        RECT 1.145 -0.300 1.445 1.065 ;
        RECT 4.285 -0.300 4.585 1.055 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.870 0.720 5.040 2.960 ;
        RECT 4.870 1.235 5.230 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.480 0.405 3.990 ;
        RECT 3.225 2.480 3.525 3.990 ;
        RECT 4.285 2.635 4.585 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 0.830 0.860 1.415 ;
        RECT 1.730 0.520 1.900 1.415 ;
        RECT 0.690 1.245 1.900 1.415 ;
        RECT 1.730 0.520 3.005 0.690 ;
        RECT 2.705 0.520 3.005 1.065 ;
        RECT 1.700 2.415 1.870 3.055 ;
        RECT 2.185 0.895 2.485 1.065 ;
        RECT 2.315 0.895 2.485 1.415 ;
        RECT 2.875 2.130 3.045 2.710 ;
        RECT 1.700 2.540 3.045 2.710 ;
        RECT 2.315 1.245 3.600 1.415 ;
        RECT 3.290 0.830 3.460 1.415 ;
        RECT 3.430 1.245 3.600 2.300 ;
        RECT 2.875 2.130 3.600 2.300 ;
        RECT 3.430 1.625 4.215 1.795 ;
        RECT 3.735 0.860 4.090 1.030 ;
        RECT 3.800 1.980 3.970 2.280 ;
        RECT 3.920 0.860 4.090 1.445 ;
        RECT 3.920 1.275 4.690 1.445 ;
        RECT 4.520 1.275 4.690 2.150 ;
        RECT 3.800 1.980 4.690 2.150 ;
  END 
END OAI33HD1XHT

MACRO OAI32HDMXHT
  CLASS  CORE ;
  FOREIGN OAI32HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.270 0.330 1.880 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.595 0.720 2.020 ;
        RECT 0.510 1.595 1.065 1.895 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.310 1.595 1.500 2.830 ;
        RECT 1.310 2.500 1.540 2.830 ;
        RECT 1.310 1.595 1.585 1.895 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.625 1.610 3.180 2.020 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.925 1.610 2.095 2.360 ;
        RECT 1.680 2.150 2.095 2.360 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 -0.300 0.430 1.065 ;
        RECT 1.170 -0.300 1.470 1.065 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.725 2.560 1.895 3.200 ;
        RECT 2.275 0.920 2.445 2.770 ;
        RECT 1.725 2.560 2.445 2.770 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 2.295 0.430 3.990 ;
        RECT 2.730 2.550 3.030 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.715 0.920 0.885 1.415 ;
        RECT 1.755 0.570 1.925 1.415 ;
        RECT 0.715 1.245 1.925 1.415 ;
        RECT 1.755 0.570 2.965 0.740 ;
        RECT 2.795 0.570 2.965 1.130 ;
  END 
END OAI32HDMXHT

MACRO OAI32HDLXHT
  CLASS  CORE ;
  FOREIGN OAI32HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.270 0.330 1.815 ;
        RECT 0.100 1.645 0.610 1.815 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.895 1.595 1.130 2.420 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.310 1.595 1.545 2.830 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.625 1.270 3.180 1.740 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.610 2.065 2.020 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 -0.300 0.430 1.065 ;
        RECT 1.170 -0.300 1.470 1.065 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.725 2.200 1.895 2.940 ;
        RECT 1.725 2.770 2.420 2.940 ;
        RECT 2.090 2.770 2.420 3.180 ;
        RECT 2.275 0.895 2.445 2.370 ;
        RECT 1.725 2.200 2.445 2.370 ;
        RECT 2.210 0.895 2.510 1.065 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 2.365 0.430 3.990 ;
        RECT 2.730 2.345 3.030 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.715 0.830 0.885 1.415 ;
        RECT 1.755 0.520 1.925 1.415 ;
        RECT 0.715 1.245 1.925 1.415 ;
        RECT 1.755 0.520 2.900 0.690 ;
        RECT 2.730 0.520 2.900 1.065 ;
        RECT 2.730 0.895 3.030 1.065 ;
  END 
END OAI32HDLXHT

MACRO OAI32HD2XHT
  CLASS  CORE ;
  FOREIGN OAI32HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.270 0.330 1.815 ;
        RECT 0.100 1.645 0.610 1.815 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.895 1.595 1.130 2.420 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.310 1.595 1.545 2.830 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.625 1.310 3.245 1.545 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.610 2.065 2.020 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 -0.300 0.430 1.065 ;
        RECT 1.170 -0.300 1.470 1.065 ;
        RECT 3.790 -0.300 4.090 1.055 ;
        RECT 4.830 -0.300 5.130 1.055 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.375 0.720 4.545 2.960 ;
        RECT 4.375 1.555 4.820 2.045 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 2.365 0.430 3.990 ;
        RECT 2.730 2.345 3.030 3.990 ;
        RECT 3.790 2.635 4.090 3.990 ;
        RECT 4.830 2.295 5.130 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.715 0.830 0.885 1.415 ;
        RECT 1.755 0.520 1.925 1.415 ;
        RECT 0.715 1.245 1.925 1.415 ;
        RECT 1.755 0.520 2.965 0.690 ;
        RECT 2.795 0.520 2.965 1.130 ;
        RECT 1.725 2.200 1.895 2.940 ;
        RECT 2.275 0.895 2.445 2.370 ;
        RECT 1.725 2.200 2.445 2.370 ;
        RECT 2.210 0.895 2.510 1.065 ;
        RECT 3.425 1.690 3.725 1.895 ;
        RECT 2.275 1.725 3.725 1.895 ;
        RECT 3.240 0.955 3.595 1.125 ;
        RECT 3.425 0.955 3.595 1.445 ;
        RECT 3.425 1.275 4.195 1.445 ;
        RECT 4.025 1.275 4.195 2.245 ;
        RECT 3.240 2.075 4.195 2.245 ;
  END 
END OAI32HD2XHT

MACRO OAI32HD1XHT
  CLASS  CORE ;
  FOREIGN OAI32HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.270 0.330 1.815 ;
        RECT 0.100 1.645 0.610 1.815 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.895 1.595 1.130 2.420 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.310 1.595 1.545 2.830 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.625 1.310 3.245 1.545 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.610 2.065 2.020 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 -0.300 0.430 1.065 ;
        RECT 1.170 -0.300 1.470 1.065 ;
        RECT 3.790 -0.300 4.090 1.055 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.375 0.720 4.545 2.960 ;
        RECT 4.375 2.500 4.820 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 2.365 0.430 3.990 ;
        RECT 2.730 2.345 3.030 3.990 ;
        RECT 3.790 2.635 4.090 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.715 0.830 0.885 1.415 ;
        RECT 1.755 0.520 1.925 1.415 ;
        RECT 0.715 1.245 1.925 1.415 ;
        RECT 1.755 0.520 2.965 0.690 ;
        RECT 2.795 0.520 2.965 1.130 ;
        RECT 1.725 2.200 1.895 2.940 ;
        RECT 2.275 0.895 2.445 2.370 ;
        RECT 1.725 2.200 2.445 2.370 ;
        RECT 2.210 0.895 2.510 1.065 ;
        RECT 3.425 1.690 3.725 1.895 ;
        RECT 2.275 1.725 3.725 1.895 ;
        RECT 3.240 0.960 3.595 1.130 ;
        RECT 3.425 0.960 3.595 1.405 ;
        RECT 3.425 1.235 4.195 1.405 ;
        RECT 4.025 1.235 4.195 2.245 ;
        RECT 3.240 2.075 4.195 2.245 ;
  END 
END OAI32HD1XHT

MACRO OAI31HDMXHT
  CLASS  CORE ;
  FOREIGN OAI31HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.270 0.310 1.815 ;
        RECT 0.100 1.645 0.610 1.815 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.895 1.595 1.130 2.420 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.310 1.595 1.545 2.830 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.610 2.065 2.020 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 -0.300 0.430 1.065 ;
        RECT 1.170 -0.300 1.470 1.065 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.725 2.200 1.895 3.210 ;
        RECT 2.275 0.860 2.445 2.370 ;
        RECT 1.725 2.200 2.445 2.370 ;
        RECT 2.275 0.860 2.770 1.220 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 2.295 0.430 3.990 ;
        RECT 2.210 2.550 2.510 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.715 0.920 0.885 1.415 ;
        RECT 1.755 0.920 1.925 1.415 ;
        RECT 0.715 1.245 1.925 1.415 ;
  END 
END OAI31HDMXHT

MACRO OAI31HDLXHT
  CLASS  CORE ;
  FOREIGN OAI31HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.270 0.335 1.815 ;
        RECT 0.100 1.645 0.610 1.815 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.895 1.595 1.130 2.420 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.310 1.595 1.545 2.830 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.610 2.065 2.020 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 -0.300 0.430 1.065 ;
        RECT 1.170 -0.300 1.470 1.065 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.725 2.200 1.895 2.940 ;
        RECT 2.275 0.830 2.445 2.370 ;
        RECT 1.725 2.200 2.445 2.370 ;
        RECT 2.275 0.830 2.770 1.230 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 2.365 0.430 3.990 ;
        RECT 2.210 2.550 2.510 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.715 0.830 0.885 1.415 ;
        RECT 1.755 0.830 1.925 1.415 ;
        RECT 0.715 1.245 1.925 1.415 ;
  END 
END OAI31HDLXHT

MACRO OAI31HD2XHT
  CLASS  CORE ;
  FOREIGN OAI31HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.270 0.330 1.880 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.660 0.720 2.020 ;
        RECT 0.510 1.660 1.105 1.830 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.290 1.595 1.460 2.360 ;
        RECT 0.860 2.150 1.460 2.360 ;
        RECT 1.290 1.595 1.560 1.895 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.610 2.065 2.020 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.065 ;
        RECT 1.145 -0.300 1.445 1.065 ;
        RECT 3.245 -0.300 3.545 1.055 ;
        RECT 4.285 -0.300 4.585 1.055 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.830 0.720 4.000 2.960 ;
        RECT 3.790 2.470 4.000 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.365 0.405 3.990 ;
        RECT 2.185 2.550 2.485 3.990 ;
        RECT 3.245 2.295 3.545 3.990 ;
        RECT 4.285 2.295 4.585 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 0.830 0.860 1.415 ;
        RECT 1.730 0.830 1.900 1.415 ;
        RECT 0.690 1.245 1.900 1.415 ;
        RECT 1.695 2.200 1.865 2.940 ;
        RECT 2.245 1.485 2.420 1.765 ;
        RECT 2.250 0.830 2.420 2.370 ;
        RECT 1.695 2.200 2.420 2.370 ;
        RECT 2.245 1.595 3.175 1.765 ;
        RECT 2.760 1.060 2.930 1.415 ;
        RECT 2.760 1.945 2.930 2.280 ;
        RECT 2.760 1.245 3.615 1.415 ;
        RECT 3.445 1.245 3.615 2.115 ;
        RECT 2.760 1.945 3.615 2.115 ;
  END 
END OAI31HD2XHT

MACRO OAI31HD1XHT
  CLASS  CORE ;
  FOREIGN OAI31HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.270 0.335 1.815 ;
        RECT 0.100 1.645 0.610 1.815 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.895 1.595 1.130 1.895 ;
        RECT 0.920 1.595 1.130 2.420 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 1.595 1.545 2.830 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.610 2.065 2.020 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 -0.300 0.430 1.065 ;
        RECT 1.170 -0.300 1.470 1.065 ;
        RECT 3.150 -0.300 3.450 1.055 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.735 0.720 3.905 2.960 ;
        RECT 3.735 2.470 4.000 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 2.365 0.430 3.990 ;
        RECT 2.210 2.705 2.510 3.990 ;
        RECT 3.150 2.295 3.450 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.715 0.830 0.885 1.415 ;
        RECT 1.755 0.830 1.925 1.415 ;
        RECT 0.715 1.245 1.925 1.415 ;
        RECT 1.725 2.200 1.895 2.840 ;
        RECT 2.305 1.060 2.475 2.370 ;
        RECT 1.725 2.200 2.475 2.370 ;
        RECT 2.305 1.595 3.080 1.765 ;
        RECT 2.600 0.545 2.945 0.715 ;
        RECT 2.665 1.945 2.835 2.280 ;
        RECT 2.775 0.545 2.945 1.415 ;
        RECT 2.775 1.245 3.555 1.415 ;
        RECT 3.385 1.245 3.555 2.115 ;
        RECT 2.665 1.945 3.555 2.115 ;
  END 
END OAI31HD1XHT

MACRO OAI22HDUXHT
  CLASS  CORE ;
  FOREIGN OAI22HDUXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.560 0.520 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.750 1.585 0.920 2.770 ;
        RECT 0.750 1.585 1.000 1.885 ;
        RECT 0.750 2.560 1.195 2.770 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.070 1.270 2.360 1.870 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.255 1.520 1.540 2.015 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.785 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.655 0.510 1.890 1.360 ;
        RECT 1.720 0.510 1.890 2.365 ;
        RECT 1.100 2.195 1.890 2.365 ;
        RECT 1.655 0.510 2.060 0.720 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.195 0.405 3.990 ;
        RECT 2.115 2.130 2.285 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.550 0.340 1.335 ;
        RECT 1.200 0.550 1.370 1.335 ;
        RECT 0.170 1.165 1.370 1.335 ;
  END 
END OAI22HDUXHT

MACRO OAI22HDMXHT
  CLASS  CORE ;
  FOREIGN OAI22HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.560 0.520 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.750 1.585 0.920 2.770 ;
        RECT 0.750 1.585 1.000 1.885 ;
        RECT 0.750 2.560 1.195 2.770 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.070 1.270 2.360 1.870 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.255 1.520 1.540 2.015 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.580 -0.300 0.880 1.145 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.670 0.510 1.890 1.360 ;
        RECT 1.720 0.510 1.890 2.365 ;
        RECT 1.100 2.195 1.890 2.365 ;
        RECT 1.670 0.510 2.060 0.720 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.395 0.405 3.990 ;
        RECT 2.115 2.330 2.285 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
END OAI22HDMXHT

MACRO OAI22HDLXHT
  CLASS  CORE ;
  FOREIGN OAI22HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.560 0.520 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.750 1.585 0.920 2.770 ;
        RECT 0.750 1.585 1.000 1.885 ;
        RECT 0.750 2.560 1.195 2.770 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.070 1.270 2.360 1.870 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.255 1.520 1.540 2.015 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.580 -0.300 0.880 1.295 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.670 0.510 1.890 1.360 ;
        RECT 1.720 0.510 1.890 2.365 ;
        RECT 1.100 2.195 1.890 2.365 ;
        RECT 1.670 0.510 2.060 0.720 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.195 0.405 3.990 ;
        RECT 2.115 2.130 2.285 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
END OAI22HDLXHT

MACRO OAI22HD2XHT
  CLASS  CORE ;
  FOREIGN OAI22HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.595 0.545 2.095 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.780 2.560 1.280 2.875 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.130 1.675 2.390 2.150 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.210 1.600 1.600 1.950 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.650 -0.300 0.950 1.065 ;
        RECT 3.290 -0.300 3.590 1.055 ;
        RECT 4.330 -0.300 4.630 1.055 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.790 0.720 4.045 1.210 ;
        RECT 3.875 0.720 4.045 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 2.330 0.430 3.990 ;
        RECT 2.210 2.330 2.510 3.990 ;
        RECT 3.290 2.295 3.590 3.990 ;
        RECT 4.330 2.295 4.630 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.195 0.830 0.365 1.415 ;
        RECT 1.235 0.520 1.405 1.415 ;
        RECT 0.195 1.245 1.405 1.415 ;
        RECT 1.235 0.520 2.445 0.690 ;
        RECT 2.275 0.520 2.445 1.130 ;
        RECT 1.780 0.895 1.950 2.350 ;
        RECT 1.170 2.180 1.950 2.350 ;
        RECT 1.690 0.895 1.990 1.065 ;
        RECT 1.780 1.315 2.740 1.485 ;
        RECT 2.570 1.315 2.740 1.765 ;
        RECT 2.570 1.595 3.220 1.765 ;
        RECT 2.740 0.965 3.090 1.135 ;
        RECT 2.805 1.945 2.975 2.280 ;
        RECT 2.920 0.965 3.090 1.415 ;
        RECT 2.920 1.245 3.375 1.415 ;
        RECT 2.805 1.945 3.525 2.115 ;
        RECT 3.525 1.320 3.535 2.114 ;
        RECT 3.535 1.330 3.545 2.114 ;
        RECT 3.545 1.340 3.555 2.114 ;
        RECT 3.555 1.350 3.565 2.114 ;
        RECT 3.565 1.360 3.575 2.114 ;
        RECT 3.575 1.370 3.585 2.114 ;
        RECT 3.585 1.380 3.595 2.114 ;
        RECT 3.595 1.390 3.605 2.114 ;
        RECT 3.605 1.400 3.615 2.114 ;
        RECT 3.615 1.410 3.625 2.114 ;
        RECT 3.625 1.420 3.635 2.114 ;
        RECT 3.635 1.430 3.645 2.114 ;
        RECT 3.645 1.440 3.655 2.114 ;
        RECT 3.655 1.450 3.665 2.114 ;
        RECT 3.665 1.460 3.675 2.114 ;
        RECT 3.675 1.470 3.685 2.114 ;
        RECT 3.685 1.480 3.695 2.114 ;
        RECT 3.460 1.255 3.470 1.499 ;
        RECT 3.470 1.265 3.480 1.509 ;
        RECT 3.480 1.275 3.490 1.519 ;
        RECT 3.490 1.285 3.500 1.529 ;
        RECT 3.500 1.295 3.510 1.539 ;
        RECT 3.510 1.305 3.520 1.549 ;
        RECT 3.520 1.310 3.526 1.560 ;
        RECT 3.375 1.245 3.385 1.415 ;
        RECT 3.385 1.245 3.395 1.425 ;
        RECT 3.395 1.245 3.405 1.435 ;
        RECT 3.405 1.245 3.415 1.445 ;
        RECT 3.415 1.245 3.425 1.455 ;
        RECT 3.425 1.245 3.435 1.465 ;
        RECT 3.435 1.245 3.445 1.475 ;
        RECT 3.445 1.245 3.455 1.485 ;
        RECT 3.455 1.245 3.461 1.495 ;
  END 
END OAI22HD2XHT

MACRO OAI22HD1XHT
  CLASS  CORE ;
  FOREIGN OAI22HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.585 0.545 2.115 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.895 1.595 1.065 2.830 ;
        RECT 0.895 2.500 1.130 2.830 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.270 2.460 1.870 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.245 1.600 1.600 1.950 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.650 -0.300 0.950 1.055 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.310 2.130 1.480 3.110 ;
        RECT 1.755 1.060 1.950 1.360 ;
        RECT 1.740 2.085 1.950 2.440 ;
        RECT 1.780 1.060 1.950 2.440 ;
        RECT 1.310 2.130 1.950 2.440 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 2.295 0.430 3.990 ;
        RECT 2.210 2.295 2.510 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.195 0.720 0.365 1.405 ;
        RECT 1.235 0.580 1.405 1.405 ;
        RECT 0.195 1.235 1.405 1.405 ;
        RECT 1.235 0.580 2.510 0.750 ;
        RECT 2.210 0.580 2.510 1.090 ;
  END 
END OAI22HD1XHT

MACRO OAI22B2HDMXHT
  CLASS  CORE ;
  FOREIGN OAI22B2HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.700 2.480 1.280 2.770 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.265 1.535 1.660 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.875 2.775 2.425 3.180 ;
    END
  END D
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.550 0.425 2.010 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.860 -0.300 1.160 0.745 ;
        RECT 1.960 -0.300 2.260 0.565 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.385 1.685 2.555 2.215 ;
        RECT 2.215 2.045 2.555 2.215 ;
        RECT 2.870 1.125 3.180 1.295 ;
        RECT 2.970 1.125 3.180 1.855 ;
        RECT 2.385 1.685 3.180 1.855 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.655 0.405 3.990 ;
        RECT 1.145 2.950 1.445 3.990 ;
        RECT 2.735 2.045 3.145 2.215 ;
        RECT 2.975 2.045 3.145 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.410 1.125 2.650 1.295 ;
        RECT 0.170 0.510 0.340 1.295 ;
        RECT 0.170 1.125 0.775 1.295 ;
        RECT 0.605 1.125 0.775 2.215 ;
        RECT 0.915 2.045 1.085 2.300 ;
        RECT 0.605 2.045 1.085 2.215 ;
        RECT 0.915 2.130 1.990 2.300 ;
        RECT 1.820 2.130 1.990 2.595 ;
        RECT 1.820 2.425 2.790 2.595 ;
        RECT 2.620 2.425 2.790 2.980 ;
  END 
END OAI22B2HDMXHT

MACRO OAI22B2HDLXHT
  CLASS  CORE ;
  FOREIGN OAI22B2HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.700 2.480 1.280 2.770 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.265 1.535 1.660 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.875 2.775 2.460 3.180 ;
    END
  END D
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.550 0.425 2.010 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.110 -0.300 2.090 0.745 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.385 1.685 2.555 2.215 ;
        RECT 2.215 2.045 2.555 2.215 ;
        RECT 2.865 0.575 3.180 0.745 ;
        RECT 2.970 0.575 3.180 1.855 ;
        RECT 2.385 1.685 3.180 1.855 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.655 0.405 3.990 ;
        RECT 1.175 2.950 1.475 3.990 ;
        RECT 2.735 2.055 3.145 2.225 ;
        RECT 2.975 2.055 3.145 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.455 1.125 2.695 1.295 ;
        RECT 0.105 1.125 0.775 1.295 ;
        RECT 0.605 1.125 0.775 2.215 ;
        RECT 0.915 2.045 1.085 2.300 ;
        RECT 0.605 2.045 1.085 2.215 ;
        RECT 0.915 2.130 1.990 2.300 ;
        RECT 1.820 2.130 1.990 2.595 ;
        RECT 1.820 2.425 2.795 2.595 ;
  END 
END OAI22B2HDLXHT

MACRO OAI221HD1XHT
  CLASS  CORE ;
  FOREIGN OAI221HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.640 0.310 2.015 ;
        RECT 0.100 1.640 0.585 1.810 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.830 1.585 1.000 2.360 ;
        RECT 0.445 2.150 1.000 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.835 1.630 2.430 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.215 1.585 1.610 1.950 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.655 1.330 3.240 1.820 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.055 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.210 2.130 1.380 3.110 ;
        RECT 1.210 2.130 3.590 2.300 ;
        RECT 3.310 0.510 3.590 1.150 ;
        RECT 3.420 0.510 3.590 2.455 ;
        RECT 3.380 2.050 3.590 2.455 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.635 0.405 3.990 ;
        RECT 2.185 2.635 2.485 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.690 0.340 1.405 ;
        RECT 1.210 0.690 1.380 1.405 ;
        RECT 2.280 1.030 2.450 1.405 ;
        RECT 0.170 1.235 2.450 1.405 ;
        RECT 1.695 0.520 1.995 1.055 ;
        RECT 1.695 0.520 3.025 0.690 ;
        RECT 2.725 0.520 3.025 1.055 ;
  END 
END OAI221HD1XHT

MACRO OAI21HDUXHT
  CLASS  CORE ;
  FOREIGN OAI21HDUXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.660 0.585 2.075 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.750 2.760 1.275 3.180 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.970 1.565 1.590 2.035 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 -0.300 0.905 0.745 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.665 0.500 1.950 1.195 ;
        RECT 1.770 0.500 1.950 2.430 ;
        RECT 1.095 2.255 1.950 2.430 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.335 0.405 3.990 ;
        RECT 1.645 2.815 1.945 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.105 1.485 1.275 ;
  END 
END OAI21HDUXHT

MACRO OAI21HDMXHT
  CLASS  CORE ;
  FOREIGN OAI21HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.310 2.010 ;
        RECT 0.100 1.520 0.520 1.820 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.700 1.580 0.870 2.360 ;
        RECT 0.450 2.150 0.870 2.360 ;
        RECT 0.700 1.580 1.065 1.765 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.245 1.610 1.610 1.950 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.575 -0.300 0.875 0.515 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.095 2.130 1.395 3.000 ;
        RECT 1.710 0.855 1.960 1.360 ;
        RECT 1.790 0.855 1.960 2.300 ;
        RECT 1.095 2.130 1.960 2.300 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.545 0.405 3.990 ;
        RECT 1.645 2.480 1.945 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 1.425 1.295 ;
  END 
END OAI21HDMXHT

MACRO OAI21HDLXHT
  CLASS  CORE ;
  FOREIGN OAI21HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.660 0.585 2.075 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.750 2.850 1.190 3.180 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.180 1.660 1.610 1.950 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.575 -0.300 0.875 0.745 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.095 2.130 1.395 2.640 ;
        RECT 1.710 0.850 1.960 1.385 ;
        RECT 1.790 0.850 1.960 2.300 ;
        RECT 1.095 2.130 1.960 2.300 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.480 0.405 3.990 ;
        RECT 1.645 2.480 1.945 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 1.425 1.295 ;
  END 
END OAI21HDLXHT

MACRO OAI21HD2XHT
  CLASS  CORE ;
  FOREIGN OAI21HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.660 0.320 2.010 ;
        RECT 0.100 1.660 0.585 1.835 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.830 1.660 1.000 2.360 ;
        RECT 0.450 2.150 1.000 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.180 1.660 1.600 1.960 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.130 ;
        RECT 2.655 -0.300 2.955 0.715 ;
        RECT 3.695 -0.300 3.995 1.055 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.240 0.720 3.410 2.960 ;
        RECT 3.240 1.270 3.590 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.545 0.405 3.990 ;
        RECT 1.695 2.905 1.995 3.990 ;
        RECT 2.655 2.295 2.955 3.990 ;
        RECT 3.695 2.295 3.995 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.895 0.340 1.480 ;
        RECT 1.210 0.895 1.380 1.480 ;
        RECT 0.170 1.310 1.380 1.480 ;
        RECT 1.760 1.305 1.950 1.475 ;
        RECT 1.210 2.140 1.380 3.120 ;
        RECT 1.760 1.060 1.930 1.475 ;
        RECT 1.780 1.305 1.950 2.310 ;
        RECT 1.210 2.140 1.950 2.310 ;
        RECT 1.780 1.530 2.585 1.700 ;
        RECT 2.170 0.480 2.340 1.285 ;
        RECT 2.170 1.945 2.340 2.280 ;
        RECT 2.170 1.115 3.060 1.285 ;
        RECT 2.890 1.115 3.060 2.115 ;
        RECT 2.170 1.945 3.060 2.115 ;
  END 
END OAI21HD2XHT

MACRO OAI21HD1XHT
  CLASS  CORE ;
  FOREIGN OAI21HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.090 1.590 0.520 2.065 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.585 1.130 2.455 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 1.585 1.670 2.015 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.660 -0.300 0.960 1.055 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.840 1.215 2.360 1.385 ;
        RECT 1.310 2.195 1.480 3.175 ;
        RECT 1.850 0.720 2.010 2.365 ;
        RECT 1.840 0.720 2.010 1.385 ;
        RECT 1.850 1.215 2.020 2.365 ;
        RECT 1.310 2.195 2.020 2.365 ;
        RECT 1.850 1.215 2.360 1.625 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 1.795 2.545 2.095 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.720 0.340 1.405 ;
        RECT 1.305 0.720 1.475 1.405 ;
        RECT 0.170 1.235 1.475 1.405 ;
  END 
END OAI21HD1XHT

MACRO OAI21B2HDMXHT
  CLASS  CORE ;
  FOREIGN OAI21B2HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.520 1.150 2.055 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 1.530 1.615 2.055 ;
    END
  END C
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.570 0.390 2.010 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.200 -0.300 1.500 0.990 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.785 2.130 1.955 2.430 ;
        RECT 2.305 0.985 2.475 2.300 ;
        RECT 1.785 2.130 2.475 2.300 ;
        RECT 2.305 1.225 2.770 1.645 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.195 2.190 0.365 3.990 ;
        RECT 1.200 2.525 1.500 3.990 ;
        RECT 2.240 2.525 2.540 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.570 1.050 0.740 2.405 ;
        RECT 0.570 1.050 0.745 1.340 ;
        RECT 0.130 1.050 0.745 1.220 ;
        RECT 0.570 2.235 0.950 2.405 ;
        RECT 0.570 1.170 2.125 1.340 ;
        RECT 1.955 1.170 2.125 1.865 ;
  END 
END OAI21B2HDMXHT

MACRO OAI21B2HDLXHT
  CLASS  CORE ;
  FOREIGN OAI21B2HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.910 1.520 1.150 2.050 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 1.530 1.660 2.050 ;
    END
  END C
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.270 0.380 1.900 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.210 -0.300 1.510 0.990 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.835 2.130 2.005 2.850 ;
        RECT 1.740 2.490 2.005 2.850 ;
        RECT 2.355 0.755 2.525 2.300 ;
        RECT 1.835 2.130 2.525 2.300 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.190 0.370 3.990 ;
        RECT 1.210 2.255 1.510 3.990 ;
        RECT 2.320 2.480 2.620 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.820 0.730 0.990 ;
        RECT 0.560 0.820 0.730 2.405 ;
        RECT 0.560 1.050 0.745 1.340 ;
        RECT 0.560 2.235 0.950 2.405 ;
        RECT 0.560 1.170 2.175 1.340 ;
        RECT 2.005 1.170 2.175 1.800 ;
  END 
END OAI21B2HDLXHT

MACRO OAI21B2HD2XHT
  CLASS  CORE ;
  FOREIGN OAI21B2HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.175 1.150 1.730 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.405 1.120 1.575 1.730 ;
        RECT 1.630 0.710 1.800 1.290 ;
        RECT 1.405 1.120 1.800 1.290 ;
        RECT 1.630 0.710 2.750 0.880 ;
        RECT 2.580 0.710 2.750 1.065 ;
        RECT 2.580 0.895 3.590 1.065 ;
        RECT 3.380 0.860 3.590 1.570 ;
        RECT 3.365 0.895 3.590 1.570 ;
    END
  END C
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.570 0.390 2.010 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.150 -0.300 1.450 0.715 ;
        RECT 2.950 -0.300 3.250 0.715 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.695 2.260 1.950 2.900 ;
        RECT 2.105 1.060 2.275 1.415 ;
        RECT 2.105 1.245 2.905 1.415 ;
        RECT 1.695 2.260 2.905 2.430 ;
        RECT 2.735 1.245 2.905 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 2.275 0.430 3.990 ;
        RECT 1.060 2.870 1.360 3.990 ;
        RECT 2.150 2.805 2.450 3.990 ;
        RECT 3.190 2.125 3.490 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.130 1.125 0.740 1.295 ;
        RECT 0.570 1.125 0.740 2.080 ;
        RECT 0.715 1.910 0.885 2.280 ;
        RECT 2.355 1.610 2.525 2.080 ;
        RECT 0.570 1.910 2.525 2.080 ;
  END 
END OAI21B2HD2XHT

MACRO OAI211HD1XHT
  CLASS  CORE ;
  FOREIGN OAI211HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.640 0.310 2.015 ;
        RECT 0.100 1.640 0.635 1.810 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.880 1.585 1.050 2.360 ;
        RECT 0.445 2.150 1.050 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.265 1.585 1.655 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.560 1.265 2.770 1.865 ;
        RECT 2.185 1.565 2.770 1.865 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.675 -0.300 0.975 1.055 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.260 2.130 1.430 3.180 ;
        RECT 0.860 2.970 1.430 3.180 ;
        RECT 1.835 0.885 2.005 2.300 ;
        RECT 2.265 0.545 2.565 1.055 ;
        RECT 1.835 0.885 2.565 1.055 ;
        RECT 1.260 2.130 2.565 2.300 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.635 0.455 3.990 ;
        RECT 1.745 2.480 2.045 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.220 0.690 0.390 1.405 ;
        RECT 1.260 0.690 1.430 1.405 ;
        RECT 0.220 1.235 1.430 1.405 ;
  END 
END OAI211HD1XHT

MACRO NOR4HDMXHT
  CLASS  CORE ;
  FOREIGN NOR4HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.255 0.615 1.800 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.800 1.585 1.150 2.020 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 1.585 1.540 2.430 ;
        RECT 1.330 1.585 1.755 1.885 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.155 1.585 2.325 2.770 ;
        RECT 1.670 2.560 2.325 2.770 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.175 -0.300 0.475 1.035 ;
        RECT 1.315 -0.300 1.615 1.035 ;
        RECT 2.455 -0.300 2.755 1.035 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.810 0.950 0.980 1.405 ;
        RECT 1.950 0.950 2.120 1.405 ;
        RECT 0.810 1.235 2.675 1.405 ;
        RECT 2.505 1.235 2.675 2.960 ;
        RECT 2.505 2.060 2.690 2.960 ;
        RECT 2.505 2.060 2.770 2.450 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.175 2.195 0.475 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
END NOR4HDMXHT

MACRO NOR4HDLXHT
  CLASS  CORE ;
  FOREIGN NOR4HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.260 0.615 1.800 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.800 1.585 1.150 2.020 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 1.585 1.540 2.840 ;
        RECT 1.330 1.585 1.755 1.885 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.155 1.585 2.325 2.430 ;
        RECT 1.740 2.080 2.325 2.430 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.175 -0.300 0.475 1.035 ;
        RECT 1.315 -0.300 1.615 1.035 ;
        RECT 2.455 -0.300 2.755 1.035 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.810 0.800 0.980 1.405 ;
        RECT 1.950 0.800 2.120 1.405 ;
        RECT 0.810 1.235 2.675 1.405 ;
        RECT 2.505 1.235 2.675 2.850 ;
        RECT 2.505 2.465 2.770 2.850 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.175 2.155 0.475 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
END NOR4HDLXHT

MACRO NOR4HD3XHT
  CLASS  CORE ;
  FOREIGN NOR4HD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.255 0.580 1.815 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 2.465 1.145 3.110 ;
        RECT 0.805 2.810 1.165 3.110 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.325 2.070 1.685 2.445 ;
        RECT 1.515 2.070 1.685 3.110 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.035 2.530 2.450 3.115 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.060 ;
        RECT 1.335 -0.300 1.505 1.360 ;
        RECT 2.375 -0.300 2.545 1.360 ;
        RECT 3.430 -0.300 3.600 0.910 ;
        RECT 4.405 -0.300 4.705 1.055 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.950 0.595 4.120 1.415 ;
        RECT 3.950 2.010 4.120 3.095 ;
        RECT 3.950 1.245 5.235 1.415 ;
        RECT 4.935 1.245 5.235 2.245 ;
        RECT 3.950 2.010 5.235 2.245 ;
        RECT 4.990 0.595 5.235 3.090 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.295 2.090 0.465 3.990 ;
        RECT 3.430 2.390 3.600 3.990 ;
        RECT 4.470 2.570 4.640 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.815 1.060 0.985 1.750 ;
        RECT 1.855 1.060 2.025 1.750 ;
        RECT 2.375 1.580 2.545 2.280 ;
        RECT 0.815 1.580 3.310 1.750 ;
        RECT 2.910 0.650 3.080 1.295 ;
        RECT 2.910 2.025 3.080 3.005 ;
        RECT 2.910 1.125 3.675 1.295 ;
        RECT 3.505 1.125 3.675 2.195 ;
        RECT 2.910 2.025 3.675 2.195 ;
        RECT 3.505 1.595 4.685 1.765 ;
  END 
END NOR4HD3XHT

MACRO NOR4HD2XHT
  CLASS  CORE ;
  FOREIGN NOR4HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.850 2.040 2.020 3.180 ;
        RECT 2.000 1.610 2.020 3.180 ;
        RECT 1.670 2.970 2.020 3.180 ;
        RECT 2.000 1.610 2.170 2.210 ;
        RECT 1.850 2.040 2.170 2.210 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.390 1.565 1.540 2.840 ;
        RECT 1.330 2.490 1.540 2.840 ;
        RECT 1.390 1.565 1.560 2.770 ;
        RECT 1.330 2.490 1.560 2.770 ;
        RECT 1.390 1.565 1.690 1.865 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.040 1.565 1.200 2.360 ;
        RECT 0.850 2.150 1.200 2.360 ;
        RECT 1.040 1.565 1.210 2.320 ;
        RECT 0.850 2.150 1.210 2.320 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.215 0.510 1.610 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.035 ;
        RECT 1.145 -0.300 1.445 1.035 ;
        RECT 2.120 -0.300 2.420 0.485 ;
        RECT 3.310 -0.300 3.610 0.455 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.715 1.125 3.055 1.295 ;
        RECT 2.885 1.125 3.055 2.360 ;
        RECT 2.715 2.090 3.055 2.360 ;
        RECT 2.715 2.150 3.250 2.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.230 2.980 2.400 3.990 ;
        RECT 3.310 3.115 3.610 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 3.345 1.520 3.660 1.690 ;
        RECT 0.170 1.790 0.340 2.620 ;
        RECT 0.690 0.800 0.860 1.960 ;
        RECT 0.170 1.790 0.860 1.960 ;
        RECT 1.730 0.775 1.900 1.385 ;
        RECT 0.690 1.215 1.900 1.385 ;
        RECT 1.730 0.775 3.515 0.945 ;
        RECT 3.345 0.775 3.515 1.690 ;
        RECT 3.490 1.520 3.660 1.845 ;
        RECT 2.365 1.670 2.535 2.710 ;
        RECT 2.520 1.540 2.690 1.840 ;
        RECT 2.365 1.670 2.690 1.840 ;
        RECT 3.695 1.125 4.010 1.295 ;
        RECT 3.760 2.055 3.930 2.710 ;
        RECT 2.365 2.540 3.930 2.710 ;
        RECT 3.840 1.125 4.010 2.225 ;
        RECT 3.760 2.055 4.010 2.225 ;
  END 
END NOR4HD2XHT

MACRO NOR4HD1XHT
  CLASS  CORE ;
  FOREIGN NOR4HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.000 2.090 2.360 2.260 ;
        RECT 2.150 1.610 2.170 2.420 ;
        RECT 2.000 1.610 2.170 2.260 ;
        RECT 2.150 2.090 2.360 2.420 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.430 1.610 1.600 3.180 ;
        RECT 1.270 2.970 1.600 3.180 ;
        RECT 1.430 1.610 1.660 1.910 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.010 1.610 1.180 2.770 ;
        RECT 0.850 2.560 1.210 2.770 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.260 0.470 1.800 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 0.745 ;
        RECT 1.135 -0.300 1.435 0.810 ;
        RECT 2.155 -0.300 2.455 0.745 ;
        RECT 3.145 -0.300 3.445 1.055 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.760 0.720 3.930 2.960 ;
        RECT 3.760 2.090 4.010 2.420 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.290 2.975 3.270 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.350 1.570 2.650 1.740 ;
        RECT 0.170 1.980 0.340 2.620 ;
        RECT 0.650 1.060 0.830 1.430 ;
        RECT 0.660 1.060 0.830 2.150 ;
        RECT 0.170 1.980 0.830 2.150 ;
        RECT 1.670 1.060 1.840 1.430 ;
        RECT 0.650 1.260 2.520 1.430 ;
        RECT 2.350 1.260 2.520 1.740 ;
        RECT 2.480 1.570 2.650 1.870 ;
        RECT 2.700 1.060 2.870 1.390 ;
        RECT 2.700 1.220 3.055 1.390 ;
        RECT 2.885 1.220 3.055 2.215 ;
        RECT 2.715 2.045 3.055 2.215 ;
        RECT 2.885 1.600 3.580 1.770 ;
  END 
END NOR4HD1XHT

MACRO NOR4B2HDMXHT
  CLASS  CORE ;
  FOREIGN NOR4B2HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.205 0.805 1.615 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.900 1.500 3.130 2.360 ;
        RECT 2.900 2.150 3.250 2.360 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.310 1.360 3.660 1.950 ;
    END
  END D
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.030 1.205 1.540 1.615 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.025 ;
        RECT 1.575 -0.300 1.875 0.485 ;
        RECT 2.595 -0.300 2.895 0.435 ;
        RECT 3.695 -0.300 3.995 0.685 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.125 0.865 4.010 1.035 ;
        RECT 3.840 0.865 4.005 3.045 ;
        RECT 3.645 2.195 4.005 3.045 ;
        RECT 3.840 0.865 4.010 2.730 ;
        RECT 3.645 2.195 4.010 2.730 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.165 0.925 3.990 ;
        RECT 1.655 2.535 1.955 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.090 0.855 0.260 1.965 ;
        RECT 0.170 1.795 0.340 2.280 ;
        RECT 0.090 0.855 0.405 1.025 ;
        RECT 1.835 1.585 2.005 1.965 ;
        RECT 0.090 1.795 2.005 1.965 ;
        RECT 1.835 1.585 2.135 1.755 ;
        RECT 1.145 0.855 1.945 1.025 ;
        RECT 1.775 0.855 1.945 1.405 ;
        RECT 1.775 1.235 2.650 1.405 ;
        RECT 2.480 1.235 2.650 2.315 ;
        RECT 1.145 2.145 2.650 2.315 ;
  END 
END NOR4B2HDMXHT

MACRO NOR4B2HD2XHT
  CLASS  CORE ;
  FOREIGN NOR4B2HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.150 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.205 0.805 1.615 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.900 1.425 3.150 2.360 ;
        RECT 2.900 2.150 3.250 2.360 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.335 1.260 3.655 1.840 ;
    END
  END D
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.030 1.205 1.540 1.615 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.025 ;
        RECT 1.665 -0.300 1.965 0.670 ;
        RECT 2.665 -0.300 2.965 0.485 ;
        RECT 3.765 -0.300 4.065 0.485 ;
        RECT 4.705 -0.300 5.005 1.005 ;
        RECT 5.745 -0.300 6.045 1.055 ;
        RECT 0.000 -0.300 6.150 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.290 0.720 5.460 2.960 ;
        RECT 5.290 1.740 5.710 1.950 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.165 0.925 3.990 ;
        RECT 1.655 2.495 1.955 3.990 ;
        RECT 4.705 2.295 5.005 3.990 ;
        RECT 5.745 2.295 6.045 3.990 ;
        RECT 0.000 3.390 6.150 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.090 0.855 0.260 1.965 ;
        RECT 0.170 1.795 0.340 2.280 ;
        RECT 0.090 0.855 0.405 1.025 ;
        RECT 1.835 1.630 2.005 1.965 ;
        RECT 0.090 1.795 2.005 1.965 ;
        RECT 1.835 1.630 2.175 1.800 ;
        RECT 1.145 0.855 2.035 1.025 ;
        RECT 1.865 0.855 2.035 1.450 ;
        RECT 1.865 1.280 2.630 1.450 ;
        RECT 2.460 1.280 2.630 2.315 ;
        RECT 1.145 2.145 2.630 2.315 ;
        RECT 2.215 0.865 4.005 1.035 ;
        RECT 3.835 0.865 4.005 2.620 ;
        RECT 3.645 2.045 4.005 2.620 ;
        RECT 3.835 1.595 4.665 1.765 ;
        RECT 4.220 1.945 4.390 2.620 ;
        RECT 4.185 1.125 4.485 1.415 ;
        RECT 4.185 1.245 5.110 1.415 ;
        RECT 4.940 1.245 5.110 2.115 ;
        RECT 4.220 1.945 5.110 2.115 ;
  END 
END NOR4B2HD2XHT

MACRO NOR4B2HD1XHT
  CLASS  CORE ;
  FOREIGN NOR4B2HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.740 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.205 0.740 1.615 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.900 1.565 3.150 2.360 ;
        RECT 2.900 2.150 3.250 2.360 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.335 1.260 3.655 1.840 ;
    END
  END D
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.965 1.205 1.540 1.615 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.025 ;
        RECT 1.665 -0.300 1.965 0.670 ;
        RECT 2.665 -0.300 2.965 0.485 ;
        RECT 3.765 -0.300 4.065 0.485 ;
        RECT 4.735 -0.300 5.035 1.055 ;
        RECT 0.000 -0.300 5.740 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.320 0.720 5.490 2.960 ;
        RECT 5.320 1.680 5.640 2.010 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.165 0.925 3.990 ;
        RECT 1.655 2.495 1.955 3.990 ;
        RECT 4.705 2.295 5.005 3.990 ;
        RECT 0.000 3.390 5.740 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.090 0.855 0.260 1.965 ;
        RECT 0.170 1.795 0.340 2.280 ;
        RECT 0.090 0.855 0.405 1.025 ;
        RECT 1.835 1.630 2.005 1.965 ;
        RECT 0.090 1.795 2.005 1.965 ;
        RECT 1.835 1.630 2.175 1.800 ;
        RECT 1.145 0.855 2.035 1.025 ;
        RECT 1.865 0.855 2.035 1.450 ;
        RECT 1.865 1.280 2.630 1.450 ;
        RECT 2.460 1.280 2.630 2.315 ;
        RECT 1.145 2.145 2.630 2.315 ;
        RECT 2.215 0.865 4.005 1.035 ;
        RECT 3.835 0.865 4.005 2.620 ;
        RECT 3.645 2.045 4.005 2.620 ;
        RECT 3.835 1.595 4.665 1.765 ;
        RECT 4.220 1.945 4.390 2.280 ;
        RECT 4.185 1.125 4.485 1.415 ;
        RECT 4.185 1.245 5.140 1.415 ;
        RECT 4.970 1.245 5.140 2.115 ;
        RECT 4.220 1.945 5.140 2.115 ;
  END 
END NOR4B2HD1XHT

MACRO NOR4B1HDMXHT
  CLASS  CORE ;
  FOREIGN NOR4B1HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.485 1.630 1.785 2.360 ;
        RECT 1.260 2.150 1.785 2.360 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.215 0.870 1.620 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.070 1.585 2.410 2.020 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.590 1.585 2.760 3.180 ;
        RECT 2.490 2.970 2.840 3.180 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.035 ;
        RECT 1.665 -0.300 1.965 1.035 ;
        RECT 2.705 -0.300 3.005 1.035 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.940 2.490 3.180 2.730 ;
        RECT 1.210 0.950 1.380 1.405 ;
        RECT 2.250 0.950 2.420 1.405 ;
        RECT 1.210 1.235 3.110 1.405 ;
        RECT 2.970 1.235 3.110 2.840 ;
        RECT 2.940 1.235 3.110 2.730 ;
        RECT 2.970 2.490 3.180 2.840 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.195 0.955 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.090 1.800 0.340 1.975 ;
        RECT 0.090 0.865 0.260 1.975 ;
        RECT 0.170 1.800 0.340 2.280 ;
        RECT 0.090 0.865 0.405 1.035 ;
        RECT 1.070 1.590 1.240 1.970 ;
        RECT 0.090 1.800 1.240 1.970 ;
  END 
END NOR4B1HDMXHT

MACRO NOR4B1HDLXHT
  CLASS  CORE ;
  FOREIGN NOR4B1HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.485 1.650 1.785 2.360 ;
        RECT 1.260 2.150 1.785 2.360 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.215 0.865 1.625 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.070 1.585 2.360 2.235 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.590 1.585 2.760 3.180 ;
        RECT 2.490 2.970 2.840 3.180 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.035 ;
        RECT 1.665 -0.300 1.965 1.035 ;
        RECT 2.705 -0.300 3.005 1.035 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.940 2.490 3.180 2.730 ;
        RECT 1.210 0.800 1.380 1.405 ;
        RECT 2.250 0.800 2.420 1.405 ;
        RECT 1.210 1.235 3.110 1.405 ;
        RECT 2.970 1.235 3.110 2.840 ;
        RECT 2.940 1.235 3.110 2.730 ;
        RECT 2.970 2.490 3.180 2.840 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.155 0.955 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.090 0.865 0.260 1.975 ;
        RECT 0.170 1.805 0.340 2.280 ;
        RECT 0.090 0.865 0.405 1.035 ;
        RECT 1.045 1.590 1.215 1.975 ;
        RECT 0.090 1.805 1.215 1.975 ;
  END 
END NOR4B1HDLXHT

MACRO NOR4B1HD2XHT
  CLASS  CORE ;
  FOREIGN NOR4B1HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.380 1.565 1.680 2.360 ;
        RECT 1.260 2.150 1.680 2.360 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.215 0.850 1.620 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.990 1.565 2.160 2.770 ;
        RECT 1.670 2.560 2.160 2.770 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.470 1.565 2.640 3.180 ;
        RECT 2.470 2.970 2.840 3.180 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.035 ;
        RECT 1.665 -0.300 1.965 1.035 ;
        RECT 2.705 -0.300 3.005 1.035 ;
        RECT 3.885 -0.300 4.185 0.715 ;
        RECT 4.925 -0.300 5.225 1.055 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.470 0.720 4.640 2.960 ;
        RECT 4.470 1.670 4.820 2.020 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.155 0.955 3.990 ;
        RECT 3.885 2.295 4.185 3.990 ;
        RECT 4.925 2.295 5.225 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.090 1.800 0.340 1.975 ;
        RECT 0.090 0.865 0.260 1.975 ;
        RECT 0.170 1.800 0.340 2.280 ;
        RECT 0.090 0.865 0.405 1.035 ;
        RECT 1.030 1.590 1.200 1.970 ;
        RECT 0.090 1.800 1.200 1.970 ;
        RECT 1.210 0.800 1.380 1.385 ;
        RECT 2.250 0.800 2.420 1.385 ;
        RECT 1.210 1.215 2.990 1.385 ;
        RECT 2.820 1.215 2.990 2.620 ;
        RECT 2.820 1.530 3.815 1.700 ;
        RECT 3.400 1.945 3.570 2.620 ;
        RECT 3.335 1.125 4.290 1.295 ;
        RECT 4.120 1.125 4.290 2.115 ;
        RECT 3.400 1.945 4.290 2.115 ;
  END 
END NOR4B1HD2XHT

MACRO NOR3HDMXHT
  CLASS  CORE ;
  FOREIGN NOR3HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.260 0.380 1.735 ;
        RECT 0.100 1.565 0.585 1.735 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.850 1.585 1.040 2.360 ;
        RECT 0.850 2.150 1.200 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.260 1.585 1.610 1.950 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.035 ;
        RECT 1.175 -0.300 1.475 0.485 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.690 0.950 0.860 1.405 ;
        RECT 0.690 1.235 1.960 1.405 ;
        RECT 1.790 0.950 1.880 2.970 ;
        RECT 1.710 0.950 1.880 1.405 ;
        RECT 1.790 1.235 1.960 2.970 ;
        RECT 1.710 2.330 1.960 2.970 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.055 0.405 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
END NOR3HDMXHT

MACRO NOR3HDLXHT
  CLASS  CORE ;
  FOREIGN NOR3HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.255 0.310 1.755 ;
        RECT 0.100 1.585 0.585 1.755 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 2.490 1.130 3.145 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.260 1.565 1.605 1.950 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 0.745 ;
        RECT 1.175 -0.300 1.475 0.745 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.625 1.125 1.955 1.295 ;
        RECT 1.740 2.085 1.955 2.775 ;
        RECT 1.785 1.125 1.955 2.775 ;
        RECT 1.710 2.135 1.955 2.775 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.200 0.405 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
END NOR3HDLXHT

MACRO NOR3HD3XHT
  CLASS  CORE ;
  FOREIGN NOR3HD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.270 0.580 1.815 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 2.560 1.230 3.105 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.260 2.145 1.675 2.365 ;
        RECT 1.505 2.145 1.675 3.085 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.060 ;
        RECT 1.335 -0.300 1.505 1.360 ;
        RECT 2.970 -0.300 3.140 0.950 ;
        RECT 4.010 -0.300 4.180 0.945 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.490 0.595 3.660 1.340 ;
        RECT 3.490 2.010 3.660 3.090 ;
        RECT 3.490 1.140 4.825 1.340 ;
        RECT 3.490 2.010 4.825 2.265 ;
        RECT 4.530 0.595 4.825 3.090 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.295 2.000 0.465 3.990 ;
        RECT 2.970 2.340 3.140 3.990 ;
        RECT 4.010 2.445 4.180 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.815 1.060 0.985 1.750 ;
        RECT 1.855 1.060 2.025 2.640 ;
        RECT 0.815 1.580 2.855 1.750 ;
        RECT 2.450 0.655 2.620 1.305 ;
        RECT 2.450 1.980 2.620 3.005 ;
        RECT 2.450 1.135 3.215 1.305 ;
        RECT 3.045 1.135 3.215 2.150 ;
        RECT 2.450 1.980 3.215 2.150 ;
        RECT 3.045 1.595 4.240 1.765 ;
  END 
END NOR3HD3XHT

MACRO NOR3HD2XHT
  CLASS  CORE ;
  FOREIGN NOR3HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.325 1.495 1.560 2.135 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.910 1.515 1.130 2.430 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.270 0.380 1.800 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.485 ;
        RECT 1.665 -0.300 1.965 0.715 ;
        RECT 2.705 -0.300 3.005 1.055 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 0.840 2.420 1.205 ;
        RECT 2.250 0.840 2.420 2.280 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.665 2.975 1.965 3.990 ;
        RECT 2.705 2.975 3.005 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 2.000 0.340 2.640 ;
        RECT 0.560 0.920 0.730 2.170 ;
        RECT 0.170 2.000 0.730 2.170 ;
        RECT 0.105 0.920 1.970 1.090 ;
        RECT 1.800 0.920 1.970 2.640 ;
        RECT 1.800 2.470 2.870 2.640 ;
        RECT 3.080 1.585 3.090 2.045 ;
        RECT 3.090 1.585 3.100 2.035 ;
        RECT 3.100 1.585 3.110 2.025 ;
        RECT 3.110 1.585 3.120 2.015 ;
        RECT 3.120 1.585 3.130 2.005 ;
        RECT 3.130 1.585 3.140 1.995 ;
        RECT 3.140 1.585 3.150 1.985 ;
        RECT 3.150 1.585 3.160 1.975 ;
        RECT 3.160 1.585 3.170 1.965 ;
        RECT 3.170 1.585 3.180 1.955 ;
        RECT 3.180 1.585 3.190 1.945 ;
        RECT 3.190 1.585 3.200 1.935 ;
        RECT 3.200 1.585 3.210 1.925 ;
        RECT 3.210 1.585 3.220 1.915 ;
        RECT 3.220 1.585 3.230 1.905 ;
        RECT 3.230 1.585 3.240 1.895 ;
        RECT 3.240 1.585 3.250 1.885 ;
        RECT 3.040 1.840 3.050 2.084 ;
        RECT 3.050 1.830 3.060 2.074 ;
        RECT 3.060 1.820 3.070 2.064 ;
        RECT 3.070 1.810 3.080 2.054 ;
        RECT 2.870 2.010 2.880 2.640 ;
        RECT 2.880 2.000 2.890 2.640 ;
        RECT 2.890 1.990 2.900 2.640 ;
        RECT 2.900 1.980 2.910 2.640 ;
        RECT 2.910 1.970 2.920 2.640 ;
        RECT 2.920 1.960 2.930 2.640 ;
        RECT 2.930 1.950 2.940 2.640 ;
        RECT 2.940 1.940 2.950 2.640 ;
        RECT 2.950 1.930 2.960 2.640 ;
        RECT 2.960 1.920 2.970 2.640 ;
        RECT 2.970 1.910 2.980 2.640 ;
        RECT 2.980 1.900 2.990 2.640 ;
        RECT 2.990 1.890 3.000 2.640 ;
        RECT 3.000 1.880 3.010 2.640 ;
        RECT 3.010 1.870 3.020 2.640 ;
        RECT 3.020 1.860 3.030 2.640 ;
        RECT 3.030 1.850 3.040 2.640 ;
        RECT 2.600 1.235 2.770 1.730 ;
        RECT 3.255 1.125 3.600 1.405 ;
        RECT 2.600 1.235 3.600 1.405 ;
        RECT 3.320 2.085 3.490 2.725 ;
        RECT 3.430 1.125 3.600 2.255 ;
        RECT 3.320 2.085 3.600 2.255 ;
  END 
END NOR3HD2XHT

MACRO NOR3HD1XHT
  CLASS  CORE ;
  FOREIGN NOR3HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.260 0.310 1.800 ;
        RECT 0.100 1.500 0.520 1.800 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.870 1.565 1.130 2.430 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.310 1.565 1.540 2.100 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.035 ;
        RECT 1.175 -0.300 1.475 0.485 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.690 1.060 0.860 1.360 ;
        RECT 0.690 1.190 1.890 1.360 ;
        RECT 1.720 1.060 1.880 3.210 ;
        RECT 1.710 1.060 1.880 1.360 ;
        RECT 1.720 1.190 1.890 3.210 ;
        RECT 1.710 2.230 1.950 3.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
END NOR3HD1XHT

MACRO NOR3B1HDMXHT
  CLASS  CORE ;
  FOREIGN NOR3B1HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 1.540 1.550 2.435 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.540 0.520 2.015 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.525 2.020 2.065 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.735 -0.300 1.715 0.595 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.120 0.840 2.370 1.295 ;
        RECT 1.075 1.125 2.370 1.295 ;
        RECT 2.200 0.840 2.290 2.970 ;
        RECT 2.120 2.330 2.290 2.970 ;
        RECT 2.200 0.840 2.370 2.500 ;
        RECT 2.120 2.330 2.370 2.500 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.645 2.735 0.945 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.500 0.340 1.295 ;
        RECT 0.170 1.125 0.890 1.295 ;
        RECT 0.720 1.125 0.890 2.365 ;
        RECT 0.105 2.195 0.890 2.365 ;
        RECT 0.720 1.545 1.070 1.845 ;
  END 
END NOR3B1HDMXHT

MACRO NOR3B1HDLXHT
  CLASS  CORE ;
  FOREIGN NOR3B1HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.260 1.655 1.615 2.360 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.545 0.520 2.015 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.650 2.880 2.175 3.180 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.745 -0.300 1.725 0.745 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.150 1.060 1.320 1.360 ;
        RECT 1.150 1.190 2.360 1.360 ;
        RECT 2.120 0.490 2.280 2.430 ;
        RECT 2.110 0.490 2.280 1.360 ;
        RECT 2.120 1.190 2.290 2.430 ;
        RECT 2.120 1.190 2.360 1.610 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.555 0.955 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 0.960 1.295 ;
        RECT 0.790 1.125 0.960 2.365 ;
        RECT 0.105 2.195 0.960 2.365 ;
        RECT 0.790 1.595 1.070 1.895 ;
  END 
END NOR3B1HDLXHT

MACRO NOR3B1HD2XHT
  CLASS  CORE ;
  FOREIGN NOR3B1HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.270 1.585 1.540 2.050 ;
        RECT 1.270 1.585 1.570 1.885 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.265 0.720 1.845 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.900 1.600 2.070 2.430 ;
        RECT 1.740 2.080 2.070 2.430 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.035 ;
        RECT 1.695 -0.300 1.995 1.035 ;
        RECT 3.275 -0.300 3.575 0.715 ;
        RECT 4.315 -0.300 4.615 1.060 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.860 0.720 4.030 2.840 ;
        RECT 3.790 2.420 4.030 2.840 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.405 0.955 3.990 ;
        RECT 3.275 2.295 3.575 3.990 ;
        RECT 4.315 2.295 4.615 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.090 0.865 0.260 2.215 ;
        RECT 0.090 0.865 0.405 1.035 ;
        RECT 0.920 1.585 1.090 2.215 ;
        RECT 0.090 2.045 1.090 2.215 ;
        RECT 1.240 0.800 1.410 1.405 ;
        RECT 1.240 1.235 2.450 1.405 ;
        RECT 2.280 0.800 2.450 2.620 ;
        RECT 2.280 1.530 3.205 1.700 ;
        RECT 2.790 1.945 2.960 2.620 ;
        RECT 2.725 1.070 3.025 1.305 ;
        RECT 2.725 1.135 3.680 1.305 ;
        RECT 3.510 1.135 3.680 2.115 ;
        RECT 2.790 1.945 3.680 2.115 ;
  END 
END NOR3B1HD2XHT

MACRO NOR3B1HD1XHT
  CLASS  CORE ;
  FOREIGN NOR3B1HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 1.585 1.540 2.430 ;
        RECT 1.330 1.585 1.725 1.885 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.265 0.760 1.845 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.965 1.600 2.360 2.020 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.035 ;
        RECT 1.695 -0.300 1.995 1.035 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.240 1.060 1.410 1.405 ;
        RECT 2.280 1.060 2.450 1.405 ;
        RECT 1.240 1.235 2.770 1.405 ;
        RECT 2.600 1.235 2.770 3.145 ;
        RECT 2.215 2.295 2.770 3.145 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.635 0.955 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.090 0.865 0.260 2.215 ;
        RECT 0.090 0.865 0.405 1.035 ;
        RECT 0.980 1.585 1.150 2.215 ;
        RECT 0.090 2.045 1.150 2.215 ;
  END 
END NOR3B1HD1XHT

MACRO NOR2HDUXHT
  CLASS  CORE ;
  FOREIGN NOR2HDUXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.230 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.090 1.740 0.355 2.490 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.885 1.450 1.130 2.110 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.195 -0.300 0.515 0.510 ;
        RECT 0.775 -0.300 1.075 0.595 ;
        RECT 0.000 -0.300 1.230 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.535 2.350 0.755 2.520 ;
        RECT 0.315 0.860 0.705 1.320 ;
        RECT 0.585 0.860 0.705 3.040 ;
        RECT 0.535 0.860 0.705 2.520 ;
        RECT 0.585 2.350 0.755 3.040 ;
        RECT 0.315 0.860 0.810 1.195 ;
        RECT 0.585 2.740 1.050 3.040 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.740 0.405 3.990 ;
        RECT 0.000 3.390 1.230 3.990 ;
    END
  END VDD
END NOR2HDUXHT

MACRO NOR2HDMXHT
  CLASS  CORE ;
  FOREIGN NOR2HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.260 0.510 1.800 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.735 1.585 1.130 2.020 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.055 ;
        RECT 1.145 -0.300 1.445 1.055 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.690 0.970 0.860 1.405 ;
        RECT 0.690 1.235 1.540 1.405 ;
        RECT 1.370 1.235 1.540 2.840 ;
        RECT 1.210 2.200 1.540 2.840 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.265 0.405 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
END NOR2HDMXHT

MACRO NOR2HDLXHT
  CLASS  CORE ;
  FOREIGN NOR2HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.265 0.310 1.735 ;
        RECT 0.100 1.565 0.585 1.735 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.765 1.585 1.130 2.020 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.055 ;
        RECT 1.145 -0.300 1.445 1.055 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.690 0.820 0.860 1.405 ;
        RECT 0.690 1.235 1.540 1.405 ;
        RECT 1.370 1.235 1.540 2.840 ;
        RECT 1.210 2.250 1.540 2.840 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.315 0.405 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
END NOR2HDLXHT

MACRO NOR2HD3XHT
  CLASS  CORE ;
  FOREIGN NOR2HD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.545 0.370 2.420 ;
        RECT 0.095 1.545 1.585 1.715 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.140 1.545 2.900 1.955 ;
        RECT 2.140 1.545 3.120 1.715 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.750 -0.300 0.920 1.010 ;
        RECT 1.790 -0.300 1.960 1.010 ;
        RECT 2.830 -0.300 3.000 1.010 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.210 0.710 0.380 1.365 ;
        RECT 1.270 0.710 1.440 1.365 ;
        RECT 2.310 0.710 2.480 1.365 ;
        RECT 2.245 2.165 2.545 2.745 ;
        RECT 0.210 1.195 3.600 1.365 ;
        RECT 3.345 1.195 3.600 2.455 ;
        RECT 2.245 2.165 3.600 2.455 ;
        RECT 3.350 0.710 3.600 3.105 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.165 2.635 0.465 3.990 ;
        RECT 1.205 2.295 1.505 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.750 1.915 0.920 2.960 ;
        RECT 0.750 1.915 1.960 2.085 ;
        RECT 1.790 1.915 1.960 3.190 ;
        RECT 2.765 2.635 3.065 3.190 ;
        RECT 1.790 2.965 3.065 3.190 ;
  END 
END NOR2HD3XHT

MACRO NOR2HD1XHT
  CLASS  CORE ;
  FOREIGN NOR2HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.265 0.510 1.800 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.795 1.585 1.190 2.015 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 0.955 ;
        RECT 1.145 -0.300 1.445 0.955 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.690 0.720 0.860 1.405 ;
        RECT 0.690 1.235 1.540 1.405 ;
        RECT 1.370 1.235 1.540 3.210 ;
        RECT 1.215 2.230 1.540 3.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
END NOR2HD1XHT

MACRO NOR2HD2XHT
  CLASS  CORE ;
  FOREIGN NOR2HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.505 1.945 0.690 2.115 ;
        RECT 0.100 1.265 0.445 1.700 ;
        RECT 0.100 1.530 0.675 1.700 ;
        RECT 0.520 1.530 0.675 3.170 ;
        RECT 0.505 1.530 0.675 2.115 ;
        RECT 0.520 1.945 0.690 3.170 ;
        RECT 1.535 2.130 1.705 3.170 ;
        RECT 0.520 3.000 1.705 3.170 ;
        RECT 1.790 1.610 1.960 2.300 ;
        RECT 1.535 2.130 1.960 2.300 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.220 1.540 1.605 1.950 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 0.435 ;
        RECT 2.055 -0.300 2.355 0.435 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.635 0.860 1.040 1.190 ;
        RECT 0.870 0.860 1.040 2.820 ;
        RECT 0.635 0.860 1.210 1.185 ;
        RECT 0.870 2.180 1.230 2.820 ;
        RECT 0.635 1.015 1.880 1.185 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.170 2.230 0.340 3.990 ;
        RECT 1.905 2.635 2.205 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
END NOR2HD2XHT

MACRO NOR2HD1XSPGHT
  CLASS  CORE ;
  FOREIGN NOR2HD1XSPGHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 0.345 0.300 0.885 3.075 ;
      LAYER V7 ;
        RECT 0.435 0.845 0.795 1.205 ;
      LAYER M7 ;
        RECT 0.345 0.835 0.995 1.215 ;
      LAYER V6 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M4 ;
        RECT 0.515 0.835 0.715 1.670 ;
      LAYER V3 ;
        RECT 0.520 1.340 0.710 1.530 ;
      LAYER M3 ;
        RECT 0.425 1.335 1.300 1.535 ;
      LAYER V2 ;
        RECT 0.930 1.340 1.120 1.530 ;
      LAYER M2 ;
        RECT 0.925 1.265 1.125 2.020 ;
      LAYER V1 ;
        RECT 0.930 1.750 1.120 1.940 ;
      LAYER M1 ;
        RECT 0.920 1.265 1.330 2.020 ;
      LAYER M6 ;
        RECT 0.515 0.300 0.715 1.705 ;
      LAYER V5 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M5 ;
        RECT 0.345 0.925 1.345 1.125 ;
      LAYER V4 ;
        RECT 0.520 0.930 0.710 1.120 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 1.575 0.300 2.115 3.075 ;
      LAYER V7 ;
        RECT 1.665 0.845 2.025 1.205 ;
      LAYER M7 ;
        RECT 1.575 0.835 2.355 1.215 ;
      LAYER V6 ;
        RECT 1.750 0.930 1.940 1.120 ;
      LAYER M4 ;
        RECT 2.155 0.835 2.355 1.680 ;
      LAYER V3 ;
        RECT 2.160 1.340 2.350 1.530 ;
      LAYER M3 ;
        RECT 1.555 1.335 2.430 1.535 ;
      LAYER V2 ;
        RECT 1.750 1.340 1.940 1.530 ;
      LAYER M2 ;
        RECT 1.745 1.270 1.945 2.170 ;
      LAYER V1 ;
        RECT 1.750 1.765 1.940 1.955 ;
      LAYER M1 ;
        RECT 1.625 1.585 1.950 2.030 ;
      LAYER M6 ;
        RECT 1.745 0.300 1.945 1.705 ;
      LAYER V5 ;
        RECT 1.750 0.930 1.940 1.120 ;
      LAYER M5 ;
        RECT 1.575 0.835 2.355 1.215 ;
      LAYER V4 ;
        RECT 2.160 0.930 2.350 1.120 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.925 -0.300 1.225 0.955 ;
        RECT 1.965 -0.300 2.265 0.955 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 2.805 0.300 3.345 3.075 ;
      LAYER V7 ;
        RECT 2.895 0.845 3.255 1.205 ;
      LAYER M7 ;
        RECT 2.565 0.835 3.345 1.215 ;
      LAYER V6 ;
        RECT 2.980 0.930 3.170 1.120 ;
      LAYER M4 ;
        RECT 2.565 0.835 2.765 2.245 ;
      LAYER V3 ;
        RECT 2.570 1.750 2.760 1.940 ;
      LAYER M3 ;
        RECT 2.080 1.745 2.900 1.945 ;
      LAYER V2 ;
        RECT 2.160 1.750 2.350 1.940 ;
      LAYER M2 ;
        RECT 2.155 1.670 2.355 2.745 ;
      LAYER V1 ;
        RECT 2.160 2.385 2.350 2.575 ;
      LAYER M1 ;
        RECT 1.510 0.720 1.680 1.405 ;
        RECT 1.510 1.235 2.300 1.405 ;
        RECT 2.130 1.235 2.300 3.190 ;
        RECT 2.035 2.210 2.300 3.190 ;
        RECT 2.035 2.210 2.360 2.745 ;
      LAYER M6 ;
        RECT 2.975 0.300 3.175 1.705 ;
      LAYER V5 ;
        RECT 2.980 0.930 3.170 1.120 ;
      LAYER M5 ;
        RECT 2.565 0.835 3.345 1.215 ;
      LAYER V4 ;
        RECT 2.570 0.930 2.760 1.120 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.925 2.295 1.225 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
END NOR2HD1XSPGHT

MACRO NOR2B1HDUXHT
  CLASS  CORE ;
  FOREIGN NOR2B1HDUXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 1.535 1.555 1.835 ;
        RECT 1.220 1.535 1.555 2.110 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.810 2.910 1.250 3.210 ;
    END
  END AN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.615 -0.300 0.935 0.440 ;
        RECT 1.645 -0.300 1.945 0.660 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.455 1.085 0.625 2.420 ;
        RECT 0.455 2.035 0.810 2.420 ;
        RECT 0.455 1.085 1.375 1.255 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.335 3.180 0.630 3.990 ;
        RECT 1.430 2.795 1.730 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.620 0.275 2.900 ;
        RECT 0.105 2.600 0.610 2.900 ;
        RECT 0.105 0.620 1.465 0.790 ;
  END 
END NOR2B1HDUXHT

MACRO NOR2B1HDMXHT
  CLASS  CORE ;
  FOREIGN NOR2B1HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.300 1.500 1.570 2.085 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.235 0.720 1.735 ;
    END
  END AN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.055 ;
        RECT 1.645 -0.300 1.945 0.505 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.240 0.970 1.410 1.320 ;
        RECT 1.240 1.150 1.935 1.320 ;
        RECT 1.765 1.150 1.935 2.840 ;
        RECT 1.710 2.200 1.950 2.840 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.265 0.955 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.090 0.885 0.260 2.215 ;
        RECT 0.090 0.885 0.405 1.055 ;
        RECT 0.090 1.915 0.405 2.215 ;
        RECT 0.920 1.565 1.090 2.085 ;
        RECT 0.090 1.915 1.090 2.085 ;
  END 
END NOR2B1HDMXHT

MACRO NOR2B1HDLXHT
  CLASS  CORE ;
  FOREIGN NOR2B1HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 1.500 1.585 2.145 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.265 0.720 1.785 ;
    END
  END AN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.055 ;
        RECT 1.645 -0.300 1.945 0.505 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.240 0.820 1.410 1.190 ;
        RECT 1.240 1.020 1.935 1.190 ;
        RECT 1.765 1.020 1.935 2.835 ;
        RECT 1.645 2.315 1.950 2.835 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.315 0.955 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.090 0.885 0.260 2.215 ;
        RECT 0.090 0.885 0.405 1.055 ;
        RECT 0.090 1.965 0.405 2.215 ;
        RECT 0.920 1.565 1.090 2.135 ;
        RECT 0.090 1.965 1.090 2.135 ;
  END 
END NOR2B1HDLXHT

MACRO NOR2B1HD2XHT
  CLASS  CORE ;
  FOREIGN NOR2B1HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.580 1.540 1.950 2.010 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.465 0.720 2.015 ;
    END
  END AN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.945 ;
        RECT 1.695 -0.300 1.995 0.945 ;
        RECT 2.735 -0.300 3.035 0.945 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.240 0.710 1.410 1.350 ;
        RECT 2.150 1.180 2.365 2.755 ;
        RECT 2.280 0.710 2.365 2.755 ;
        RECT 1.695 2.245 2.365 2.755 ;
        RECT 2.280 0.710 2.450 1.350 ;
        RECT 1.240 1.180 2.450 1.350 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.635 0.955 3.990 ;
        RECT 2.895 2.230 3.175 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.090 1.115 0.260 2.365 ;
        RECT 0.090 1.115 0.405 1.285 ;
        RECT 0.900 1.530 1.070 2.365 ;
        RECT 0.090 2.195 1.380 2.365 ;
        RECT 0.900 1.530 1.225 1.700 ;
        RECT 1.210 2.195 1.380 3.170 ;
        RECT 2.545 1.595 2.715 3.170 ;
        RECT 1.210 3.000 2.715 3.170 ;
        RECT 2.545 1.595 2.855 1.765 ;
  END 
END NOR2B1HD2XHT

MACRO NAND4HDMXHT
  CLASS  CORE ;
  FOREIGN NAND4HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 2.495 0.805 2.980 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.850 0.920 1.040 1.820 ;
        RECT 0.850 0.920 1.200 1.130 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.220 1.330 1.610 1.800 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.640 2.490 1.940 3.205 ;
        RECT 1.640 2.490 2.020 2.770 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.235 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.965 1.125 2.360 1.295 ;
        RECT 2.150 1.125 2.360 2.215 ;
        RECT 0.625 2.045 2.360 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.145 0.275 3.990 ;
        RECT 0.105 2.145 0.405 2.315 ;
        RECT 1.055 2.925 1.355 3.990 ;
        RECT 2.120 2.930 2.290 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
END NAND4HDMXHT

MACRO NAND4HDLXHT
  CLASS  CORE ;
  FOREIGN NAND4HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 2.395 0.830 2.840 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.850 0.660 1.200 1.130 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.260 1.330 1.585 1.755 ;
        RECT 1.260 1.330 1.610 1.550 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.630 0.510 2.065 0.880 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.265 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.060 2.200 2.215 ;
        RECT 0.625 2.045 2.200 2.215 ;
        RECT 2.030 1.670 2.360 2.020 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.045 0.275 3.990 ;
        RECT 0.105 2.045 0.405 2.215 ;
        RECT 1.145 2.625 1.445 3.990 ;
        RECT 1.995 2.625 2.295 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
END NAND4HDLXHT

MACRO NAND4HD3XHT
  CLASS  CORE ;
  FOREIGN NAND4HD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.090 1.255 0.635 1.800 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.755 2.460 1.155 2.885 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 0.620 1.695 1.225 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.720 2.460 2.195 2.835 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.060 ;
        RECT 3.430 -0.300 3.600 0.910 ;
        RECT 4.470 -0.300 4.640 0.780 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.950 0.715 4.120 1.355 ;
        RECT 3.950 2.025 4.120 3.005 ;
        RECT 3.950 1.185 5.235 1.355 ;
        RECT 4.885 1.185 5.235 2.360 ;
        RECT 3.950 2.025 5.235 2.360 ;
        RECT 4.990 0.715 5.235 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.295 1.980 0.465 3.990 ;
        RECT 1.335 1.980 1.505 3.990 ;
        RECT 2.375 1.980 2.545 3.990 ;
        RECT 3.430 2.390 3.600 3.990 ;
        RECT 4.470 2.570 4.640 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.815 1.580 0.985 2.280 ;
        RECT 1.855 1.580 2.025 2.280 ;
        RECT 2.375 1.060 2.545 1.750 ;
        RECT 0.815 1.580 3.310 1.750 ;
        RECT 2.910 0.650 3.080 1.290 ;
        RECT 2.910 1.980 3.080 2.960 ;
        RECT 2.910 1.120 3.675 1.290 ;
        RECT 3.505 1.120 3.675 2.150 ;
        RECT 2.910 1.980 3.675 2.150 ;
        RECT 3.505 1.595 4.700 1.765 ;
  END 
END NAND4HD3XHT

MACRO NAND4HD2XHT
  CLASS  CORE ;
  FOREIGN NAND4HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.510 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 2.395 0.875 2.850 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.850 0.660 1.200 1.130 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.260 1.330 1.610 1.820 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.630 0.510 2.065 0.895 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.265 ;
        RECT 3.065 -0.300 3.365 0.935 ;
        RECT 4.105 -0.300 4.405 1.055 ;
        RECT 0.000 -0.300 4.510 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.650 0.720 3.820 2.965 ;
        RECT 3.650 1.740 4.110 1.950 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.045 0.275 3.990 ;
        RECT 0.105 2.045 0.405 2.215 ;
        RECT 1.210 2.560 1.380 3.990 ;
        RECT 2.035 2.625 2.335 3.990 ;
        RECT 3.065 2.335 3.365 3.990 ;
        RECT 4.170 2.230 4.340 3.990 ;
        RECT 0.000 3.390 4.510 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.965 1.125 2.135 2.215 ;
        RECT 0.625 2.045 2.135 2.215 ;
        RECT 1.965 1.125 2.265 1.295 ;
        RECT 1.965 1.585 3.025 1.755 ;
        RECT 2.580 0.720 2.750 1.405 ;
        RECT 2.610 1.935 2.780 2.620 ;
        RECT 2.580 1.235 3.440 1.405 ;
        RECT 3.270 1.235 3.440 2.105 ;
        RECT 2.610 1.935 3.440 2.105 ;
  END 
END NAND4HD2XHT

MACRO NAND4HD1XHT
  CLASS  CORE ;
  FOREIGN NAND4HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.310 2.020 ;
        RECT 0.100 1.585 0.585 1.755 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.850 0.660 1.210 1.130 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.260 1.330 1.610 1.820 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.670 0.510 2.105 0.895 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.295 ;
        RECT 3.095 -0.300 3.395 0.715 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.680 0.720 3.850 2.965 ;
        RECT 3.680 1.670 4.000 2.020 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.595 0.405 3.990 ;
        RECT 1.135 2.595 1.435 3.990 ;
        RECT 2.035 2.595 2.335 3.990 ;
        RECT 3.095 2.295 3.395 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.005 1.125 2.175 2.215 ;
        RECT 0.625 2.045 2.175 2.215 ;
        RECT 2.005 1.125 2.305 1.295 ;
        RECT 2.005 1.585 3.025 1.755 ;
        RECT 2.610 1.935 2.780 2.280 ;
        RECT 2.515 1.125 3.395 1.295 ;
        RECT 3.225 1.125 3.395 2.105 ;
        RECT 2.610 1.935 3.395 2.105 ;
        RECT 3.225 1.520 3.470 1.820 ;
  END 
END NAND4HD1XHT

MACRO NAND4B2HDMXHT
  CLASS  CORE ;
  FOREIGN NAND4B2HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.510 2.905 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.260 2.190 1.730 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.455 1.590 3.295 1.760 ;
        RECT 2.895 1.590 3.295 1.950 ;
    END
  END D
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.240 2.765 3.685 3.180 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.235 ;
        RECT 3.125 -0.300 3.425 1.295 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.365 0.900 1.535 2.215 ;
        RECT 1.365 0.900 2.850 1.080 ;
        RECT 1.175 2.045 2.575 2.215 ;
        RECT 2.560 0.720 2.850 1.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 2.310 0.890 3.990 ;
        RECT 1.790 2.765 1.960 3.990 ;
        RECT 2.890 2.765 3.060 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.135 1.755 ;
        RECT 1.395 2.415 1.565 2.980 ;
        RECT 3.405 2.165 3.575 2.585 ;
        RECT 1.395 2.415 3.575 2.585 ;
        RECT 3.710 1.060 3.880 2.335 ;
        RECT 3.405 2.165 3.880 2.335 ;
  END 
END NAND4B2HDMXHT

MACRO NAND4B2HDLXHT
  CLASS  CORE ;
  FOREIGN NAND4B2HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.510 2.905 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.660 0.660 1.830 1.540 ;
        RECT 1.660 1.330 2.020 1.540 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.075 0.510 2.505 0.895 ;
    END
  END D
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.900 2.745 3.250 3.180 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.715 ;
        RECT 2.735 -0.300 3.035 0.785 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.385 1.125 2.770 1.295 ;
        RECT 2.560 1.125 2.770 2.215 ;
        RECT 1.065 2.045 2.770 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 2.525 0.890 3.990 ;
        RECT 1.615 2.765 1.915 3.990 ;
        RECT 2.420 2.745 2.720 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.065 1.755 ;
        RECT 1.225 2.395 1.545 2.585 ;
        RECT 3.110 2.100 3.280 2.565 ;
        RECT 1.225 2.395 3.280 2.565 ;
        RECT 3.350 0.510 3.520 2.270 ;
        RECT 3.110 2.100 3.520 2.270 ;
  END 
END NAND4B2HDLXHT

MACRO NAND4B2HD2XHT
  CLASS  CORE ;
  FOREIGN NAND4B2HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.150 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.490 2.905 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.965 1.270 3.295 1.820 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.280 0.510 3.755 0.880 ;
    END
  END D
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.850 0.510 1.245 0.925 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.500 -0.300 0.670 0.810 ;
        RECT 1.615 -0.300 1.915 1.265 ;
        RECT 4.690 -0.300 4.990 1.055 ;
        RECT 5.730 -0.300 6.030 1.055 ;
        RECT 0.000 -0.300 6.150 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.275 0.720 5.445 2.965 ;
        RECT 5.275 1.670 5.640 2.050 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.670 2.745 0.970 3.990 ;
        RECT 1.680 1.980 1.850 3.990 ;
        RECT 2.685 2.625 2.985 3.990 ;
        RECT 3.630 2.625 3.930 3.990 ;
        RECT 4.690 2.635 4.990 3.990 ;
        RECT 5.730 2.295 6.030 3.990 ;
        RECT 0.000 3.390 6.150 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 2.110 0.905 2.280 ;
        RECT 0.735 2.110 0.905 2.565 ;
        RECT 0.735 2.395 1.500 2.565 ;
        RECT 1.330 2.395 1.500 2.790 ;
        RECT 1.085 1.125 1.385 2.215 ;
        RECT 1.085 1.525 2.615 1.695 ;
        RECT 3.645 1.060 3.815 2.215 ;
        RECT 2.135 2.045 3.815 2.215 ;
        RECT 3.645 1.585 4.620 1.755 ;
        RECT 4.175 1.060 4.345 1.405 ;
        RECT 4.205 1.935 4.375 2.620 ;
        RECT 4.175 1.235 4.990 1.405 ;
        RECT 4.820 1.235 4.990 2.105 ;
        RECT 4.205 1.935 4.990 2.105 ;
        RECT 4.820 1.520 5.065 1.820 ;
  END 
END NAND4B2HD2XHT

MACRO NAND4B2HD1XHT
  CLASS  CORE ;
  FOREIGN NAND4B2HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.740 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.490 2.905 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.970 1.270 3.230 1.820 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.270 0.510 3.825 0.880 ;
    END
  END D
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.850 0.510 1.245 0.925 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.500 -0.300 0.670 0.810 ;
        RECT 1.610 -0.300 1.910 1.265 ;
        RECT 4.780 -0.300 5.080 1.055 ;
        RECT 0.000 -0.300 5.740 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.365 0.720 5.535 2.965 ;
        RECT 5.365 1.670 5.640 2.050 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.670 2.745 0.970 3.990 ;
        RECT 1.610 2.045 1.910 3.990 ;
        RECT 2.680 2.395 2.980 3.990 ;
        RECT 3.780 2.625 4.080 3.990 ;
        RECT 4.780 2.295 5.080 3.990 ;
        RECT 0.000 3.390 5.740 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 2.110 0.905 2.280 ;
        RECT 0.735 2.110 0.905 2.565 ;
        RECT 0.735 2.395 1.400 2.565 ;
        RECT 1.230 2.395 1.400 3.030 ;
        RECT 1.085 1.125 1.385 1.295 ;
        RECT 1.215 1.125 1.385 2.215 ;
        RECT 1.085 2.045 1.385 2.215 ;
        RECT 1.215 1.590 2.545 1.760 ;
        RECT 2.375 1.525 2.545 1.825 ;
        RECT 3.675 1.060 3.845 2.215 ;
        RECT 2.130 2.045 3.845 2.215 ;
        RECT 3.675 1.585 4.710 1.755 ;
        RECT 4.265 1.060 4.435 1.405 ;
        RECT 4.295 1.935 4.465 2.280 ;
        RECT 4.265 1.235 5.080 1.405 ;
        RECT 4.910 1.235 5.080 2.105 ;
        RECT 4.295 1.935 5.080 2.105 ;
        RECT 4.910 1.520 5.185 1.820 ;
  END 
END NAND4B2HD1XHT

MACRO NAND4B1HDLXHT
  CLASS  CORE ;
  FOREIGN NAND4B1HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.225 0.510 1.610 0.895 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.320 2.840 ;
        RECT 0.100 2.470 0.520 2.705 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.670 1.330 2.025 1.765 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.080 0.510 2.505 0.895 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.715 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.160 2.045 1.330 2.830 ;
        RECT 2.385 1.125 2.770 1.295 ;
        RECT 2.560 1.125 2.770 2.215 ;
        RECT 1.160 2.045 2.770 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.585 2.905 0.885 3.990 ;
        RECT 1.605 2.595 1.905 3.990 ;
        RECT 2.465 2.745 2.765 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.065 1.755 ;
  END 
END NAND4B1HDLXHT

MACRO NAND4B1HD2XHT
  CLASS  CORE ;
  FOREIGN NAND4B1HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.255 0.660 1.610 1.130 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.510 2.905 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.670 1.330 2.020 1.820 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.070 0.510 2.505 0.895 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.715 ;
        RECT 3.465 -0.300 3.765 1.005 ;
        RECT 4.505 -0.300 4.805 1.055 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.050 0.720 4.220 2.965 ;
        RECT 4.050 1.740 4.500 1.950 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.845 0.860 3.990 ;
        RECT 1.650 2.690 1.950 3.990 ;
        RECT 2.435 2.625 2.735 3.990 ;
        RECT 3.465 2.565 3.765 3.990 ;
        RECT 4.505 2.295 4.805 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.065 1.755 ;
        RECT 1.200 2.045 1.370 3.035 ;
        RECT 2.405 1.125 2.705 1.295 ;
        RECT 2.535 1.125 2.705 2.215 ;
        RECT 1.200 2.045 2.705 2.215 ;
        RECT 2.535 1.585 3.425 1.755 ;
        RECT 2.980 1.060 3.150 1.405 ;
        RECT 3.010 1.935 3.180 2.620 ;
        RECT 2.980 1.235 3.870 1.405 ;
        RECT 3.700 1.235 3.870 2.105 ;
        RECT 3.010 1.935 3.870 2.105 ;
  END 
END NAND4B1HD2XHT

MACRO NAND4B1HD1XHT
  CLASS  CORE ;
  FOREIGN NAND4B1HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.510 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.255 0.660 1.610 1.130 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.510 2.905 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.670 1.330 1.960 1.820 ;
        RECT 1.670 1.330 2.020 1.550 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.070 0.510 2.505 0.895 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.715 ;
        RECT 3.495 -0.300 3.795 1.055 ;
        RECT 0.000 -0.300 4.510 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.080 0.720 4.250 2.960 ;
        RECT 4.080 1.670 4.410 2.020 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.845 0.860 3.990 ;
        RECT 1.650 2.690 1.950 3.990 ;
        RECT 2.435 2.625 2.735 3.990 ;
        RECT 3.495 2.295 3.795 3.990 ;
        RECT 0.000 3.390 4.510 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.065 1.755 ;
        RECT 1.200 2.045 1.370 3.035 ;
        RECT 2.405 1.125 2.705 1.295 ;
        RECT 2.535 1.125 2.705 2.215 ;
        RECT 1.200 2.045 2.705 2.215 ;
        RECT 2.535 1.585 3.425 1.755 ;
        RECT 2.980 1.060 3.150 1.405 ;
        RECT 3.010 1.935 3.180 2.280 ;
        RECT 2.980 1.235 3.840 1.405 ;
        RECT 3.670 1.235 3.840 2.105 ;
        RECT 3.010 1.935 3.840 2.105 ;
  END 
END NAND4B1HD1XHT

MACRO NAND3ODHDHT
  CLASS  CORE ;
  FOREIGN NAND3ODHDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.295 1.265 1.540 1.820 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.830 0.510 1.065 0.990 ;
        RECT 0.830 0.510 1.195 0.720 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.395 0.520 2.835 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.415 -0.300 1.715 0.745 ;
        RECT 2.355 -0.300 2.655 0.715 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 2.940 0.720 3.180 1.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 2.530 0.890 3.990 ;
        RECT 1.570 2.595 1.870 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.215 ;
        RECT 1.845 1.520 2.015 2.215 ;
        RECT 0.105 2.045 2.015 2.215 ;
        RECT 1.935 1.125 2.365 1.295 ;
        RECT 2.195 1.125 2.365 2.280 ;
        RECT 2.195 1.585 2.835 1.755 ;
  END 
END NAND3ODHDHT

MACRO NAND3HDMXHT
  CLASS  CORE ;
  FOREIGN NAND3HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.540 0.310 2.015 ;
        RECT 0.100 1.540 0.555 1.840 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.815 1.265 1.135 1.800 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.315 0.505 1.485 1.820 ;
        RECT 1.315 1.520 1.530 1.820 ;
        RECT 1.265 0.505 1.605 0.730 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.300 0.455 1.295 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.665 1.060 1.955 1.360 ;
        RECT 1.735 1.060 1.955 2.215 ;
        RECT 0.625 2.045 1.955 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.375 0.405 3.990 ;
        RECT 1.145 2.925 1.445 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
END NAND3HDMXHT

MACRO NAND3HDLXHT
  CLASS  CORE ;
  FOREIGN NAND3HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 2.395 0.860 2.845 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.880 1.265 1.130 1.820 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.225 0.510 1.485 0.925 ;
        RECT 1.310 0.510 1.485 1.820 ;
        RECT 1.310 1.520 1.530 1.820 ;
        RECT 1.225 0.510 1.605 0.720 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.300 0.455 1.295 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.665 1.060 1.950 1.360 ;
        RECT 1.740 1.060 1.950 2.215 ;
        RECT 0.625 2.045 1.950 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.045 0.275 3.990 ;
        RECT 0.105 2.045 0.405 2.215 ;
        RECT 1.145 2.595 1.445 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
END NAND3HDLXHT

MACRO NAND3HD3XHT
  CLASS  CORE ;
  FOREIGN NAND3HD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.510 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.270 0.495 1.800 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 2.460 0.950 2.770 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.895 0.710 1.130 1.235 ;
        RECT 0.895 0.710 1.635 0.880 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.225 -0.300 0.525 1.060 ;
        RECT 2.610 -0.300 2.780 0.910 ;
        RECT 3.650 -0.300 3.820 0.780 ;
        RECT 0.000 -0.300 4.510 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.130 2.010 3.300 2.990 ;
        RECT 3.125 0.595 3.305 1.340 ;
        RECT 3.125 1.170 4.415 1.340 ;
        RECT 3.130 2.010 4.415 2.265 ;
        RECT 4.170 0.595 4.415 2.990 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.950 0.405 3.990 ;
        RECT 1.150 2.530 1.320 3.990 ;
        RECT 2.610 2.390 2.780 3.990 ;
        RECT 3.650 2.445 3.820 3.990 ;
        RECT 0.000 3.390 4.510 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.580 1.060 1.750 2.215 ;
        RECT 0.535 2.045 1.815 2.215 ;
        RECT 1.580 1.580 2.505 1.750 ;
        RECT 2.090 0.655 2.260 1.300 ;
        RECT 2.090 2.025 2.260 3.005 ;
        RECT 2.090 1.130 2.855 1.300 ;
        RECT 2.685 1.130 2.855 2.195 ;
        RECT 2.090 2.025 2.855 2.195 ;
        RECT 2.685 1.595 3.880 1.765 ;
  END 
END NAND3HD3XHT

MACRO NAND3HD2XHT
  CLASS  CORE ;
  FOREIGN NAND3HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 2.395 0.815 2.880 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.815 1.265 1.130 1.820 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.265 0.510 1.485 0.725 ;
        RECT 1.310 0.510 1.485 1.820 ;
        RECT 1.310 1.520 1.520 1.820 ;
        RECT 1.265 0.510 1.605 0.720 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.295 ;
        RECT 2.590 -0.300 2.890 1.055 ;
        RECT 3.630 -0.300 3.930 1.055 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.175 0.720 3.345 2.965 ;
        RECT 3.175 1.740 3.705 1.950 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.045 0.275 3.990 ;
        RECT 0.105 2.045 0.405 2.215 ;
        RECT 1.145 2.625 1.445 3.990 ;
        RECT 2.590 2.295 2.890 3.990 ;
        RECT 3.630 2.295 3.930 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.665 1.060 1.910 1.360 ;
        RECT 1.735 1.060 1.910 2.215 ;
        RECT 0.625 2.045 1.910 2.215 ;
        RECT 1.735 1.585 2.520 1.755 ;
        RECT 2.010 0.620 2.350 0.790 ;
        RECT 2.180 0.620 2.350 1.405 ;
        RECT 2.240 1.935 2.410 2.735 ;
        RECT 2.040 2.565 2.410 2.735 ;
        RECT 2.180 1.235 2.920 1.405 ;
        RECT 2.750 1.235 2.920 2.105 ;
        RECT 2.240 1.935 2.920 2.105 ;
        RECT 2.750 1.520 2.965 1.820 ;
  END 
END NAND3HD2XHT

MACRO NAND3HD1XHT
  CLASS  CORE ;
  FOREIGN NAND3HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.505 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.870 1.265 1.130 1.820 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.325 1.425 1.555 2.015 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.055 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.000 0.860 2.640 ;
        RECT 0.690 2.195 1.950 2.375 ;
        RECT 1.730 0.715 1.905 1.360 ;
        RECT 1.735 0.715 1.905 2.620 ;
        RECT 1.735 1.980 1.950 2.620 ;
        RECT 1.730 2.195 1.950 2.620 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.285 0.405 3.990 ;
        RECT 1.145 2.625 1.445 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
END NAND3HD1XHT

MACRO NAND3B1HDMXHT
  CLASS  CORE ;
  FOREIGN NAND3B1HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.285 1.265 1.540 1.820 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.510 2.905 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.750 0.510 1.940 1.820 ;
        RECT 1.750 1.520 2.000 1.820 ;
        RECT 1.675 0.510 2.015 0.720 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.095 2.045 2.365 2.215 ;
        RECT 2.120 1.060 2.365 1.360 ;
        RECT 2.180 1.060 2.290 3.160 ;
        RECT 2.120 2.045 2.290 3.160 ;
        RECT 2.180 1.060 2.365 2.425 ;
        RECT 2.120 2.045 2.365 2.425 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 2.860 0.890 3.990 ;
        RECT 1.525 2.925 1.825 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.100 1.755 ;
  END 
END NAND3B1HDMXHT

MACRO NAND3B1HDLXHT
  CLASS  CORE ;
  FOREIGN NAND3B1HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.285 1.265 1.540 1.820 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.510 2.905 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.720 0.510 1.910 1.840 ;
        RECT 1.720 1.540 2.000 1.840 ;
        RECT 1.675 0.510 2.015 0.735 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 0.855 2.370 1.360 ;
        RECT 2.120 1.060 2.370 1.360 ;
        RECT 2.200 0.855 2.290 2.830 ;
        RECT 2.120 2.045 2.290 2.830 ;
        RECT 2.200 0.855 2.370 2.215 ;
        RECT 1.095 2.045 2.370 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 2.530 0.890 3.990 ;
        RECT 1.525 2.595 1.825 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.100 1.755 ;
  END 
END NAND3B1HDLXHT

MACRO NAND3B1HD1XHT
  CLASS  CORE ;
  FOREIGN NAND3B1HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.260 1.200 1.820 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.080 0.510 2.425 0.945 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.425 0.735 2.015 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.730 -0.300 1.900 1.120 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 0.715 0.270 2.750 ;
        RECT 0.100 0.715 0.340 1.360 ;
        RECT 0.100 2.085 0.340 2.750 ;
        RECT 0.100 2.195 1.380 2.365 ;
        RECT 1.210 2.000 1.380 2.640 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.625 0.925 3.990 ;
        RECT 1.665 2.285 1.965 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.500 1.585 2.515 1.755 ;
        RECT 2.215 1.125 2.515 2.215 ;
  END 
END NAND3B1HD1XHT

MACRO NAND2ODHDHT
  CLASS  CORE ;
  FOREIGN NAND2ODHDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.420 0.505 1.000 0.720 ;
        RECT 0.830 0.505 1.000 0.880 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.310 2.015 ;
        RECT 0.100 1.520 0.485 1.820 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.180 -0.300 1.350 1.360 ;
        RECT 1.060 1.060 1.350 1.360 ;
        RECT 1.935 -0.300 2.235 0.715 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 2.520 0.720 2.770 1.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.195 0.405 3.990 ;
        RECT 1.145 2.195 1.445 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 0.835 1.295 ;
        RECT 0.665 1.125 0.835 2.370 ;
        RECT 0.665 2.070 0.860 2.370 ;
        RECT 0.665 1.540 1.525 1.840 ;
        RECT 1.580 1.060 1.900 1.360 ;
        RECT 1.730 1.060 1.900 2.310 ;
        RECT 1.730 1.585 2.415 1.755 ;
  END 
END NAND2ODHDHT

MACRO NAND2HDUXHT
  CLASS  CORE ;
  FOREIGN NAND2HDUXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.230 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.205 0.525 0.690 0.695 ;
        RECT 0.520 0.525 0.690 1.050 ;
        RECT 0.520 0.860 1.140 1.050 ;
        RECT 0.920 0.860 1.140 1.190 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.610 0.390 2.260 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.890 -0.300 1.060 0.500 ;
        RECT 0.000 -0.300 1.230 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.170 1.060 0.340 1.430 ;
        RECT 0.170 1.250 0.750 1.430 ;
        RECT 0.570 1.250 0.750 2.770 ;
        RECT 0.570 2.250 0.865 2.770 ;
        RECT 0.350 2.560 0.865 2.770 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.950 0.405 3.990 ;
        RECT 0.630 2.950 0.930 3.990 ;
        RECT 0.000 3.390 1.230 3.990 ;
    END
  END VDD
END NAND2HDUXHT

MACRO NAND2HDMXHT
  CLASS  CORE ;
  FOREIGN NAND2HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.265 0.585 1.730 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 2.500 0.720 2.980 ;
        RECT 0.510 2.680 1.040 2.980 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.065 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.690 1.915 0.860 2.280 ;
        RECT 1.145 1.125 1.540 1.295 ;
        RECT 1.330 1.125 1.540 2.085 ;
        RECT 0.690 1.915 1.540 2.085 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.160 2.040 0.330 3.990 ;
        RECT 0.160 2.040 0.340 2.340 ;
        RECT 1.145 2.330 1.475 2.500 ;
        RECT 1.305 2.330 1.475 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
END NAND2HDMXHT

MACRO NAND2HDLXHT
  CLASS  CORE ;
  FOREIGN NAND2HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.520 0.510 0.690 0.990 ;
        RECT 0.520 0.510 1.195 0.720 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 2.500 0.720 2.865 ;
        RECT 0.510 2.500 1.125 2.670 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.170 -0.300 0.340 1.360 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.690 1.660 0.860 2.280 ;
        RECT 1.145 1.125 1.540 1.295 ;
        RECT 1.330 1.125 1.540 1.830 ;
        RECT 0.690 1.660 1.540 1.830 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.150 2.040 0.320 3.990 ;
        RECT 0.150 2.040 0.340 2.340 ;
        RECT 1.145 2.105 1.475 2.275 ;
        RECT 1.305 2.105 1.475 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
END NAND2HDLXHT

MACRO NAND2HD2XHT
  CLASS  CORE ;
  FOREIGN NAND2HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.610 0.310 2.625 ;
        RECT 0.100 1.610 0.730 1.780 ;
        RECT 2.150 1.585 2.460 1.755 ;
        RECT 2.290 1.585 2.460 2.625 ;
        RECT 0.100 2.455 2.460 2.625 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.265 1.365 1.820 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.245 -0.300 0.545 1.055 ;
        RECT 2.330 -0.300 2.630 1.055 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.355 0.480 1.525 1.055 ;
        RECT 1.290 0.885 1.770 1.055 ;
        RECT 1.290 0.920 2.020 1.055 ;
        RECT 1.590 0.885 1.770 2.215 ;
        RECT 1.590 0.920 2.020 1.130 ;
        RECT 0.770 2.045 2.110 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.250 2.805 0.550 3.990 ;
        RECT 1.290 2.805 1.590 3.990 ;
        RECT 2.330 2.805 2.630 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
END NAND2HD2XHT

MACRO NAND2HD3XHT
  CLASS  CORE ;
  FOREIGN NAND2HD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.270 0.310 1.795 ;
        RECT 0.100 1.625 1.425 1.795 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.650 1.630 2.015 1.955 ;
        RECT 1.650 1.630 3.135 1.800 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.055 ;
        RECT 1.145 -0.300 1.445 1.055 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.170 1.985 0.340 2.965 ;
        RECT 0.170 1.985 1.380 2.155 ;
        RECT 0.170 2.145 3.595 2.155 ;
        RECT 1.210 1.985 1.380 2.965 ;
        RECT 1.210 2.145 2.480 2.315 ;
        RECT 2.310 1.060 2.480 1.445 ;
        RECT 2.310 1.985 2.480 2.965 ;
        RECT 2.310 1.275 3.595 1.445 ;
        RECT 2.310 1.985 3.595 2.220 ;
        RECT 1.210 2.145 3.595 2.220 ;
        RECT 3.350 0.585 3.595 2.965 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.400 0.860 3.990 ;
        RECT 1.695 2.740 1.995 3.990 ;
        RECT 2.830 2.400 3.000 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 0.720 0.860 1.435 ;
        RECT 1.760 0.500 1.930 1.435 ;
        RECT 0.690 1.265 1.930 1.435 ;
        RECT 1.760 0.500 3.065 0.670 ;
        RECT 2.765 0.500 3.065 1.075 ;
  END 
END NAND2HD3XHT

MACRO NAND2HD1XHT
  CLASS  CORE ;
  FOREIGN NAND2HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.500 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 1.265 1.540 1.820 ;
        RECT 1.030 1.520 1.540 1.820 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.055 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.195 0.405 2.705 ;
        RECT 0.680 0.885 0.850 2.365 ;
        RECT 0.680 2.145 1.445 2.365 ;
        RECT 0.105 2.195 1.445 2.365 ;
        RECT 1.145 2.145 1.445 2.720 ;
        RECT 1.155 0.545 1.455 1.055 ;
        RECT 0.680 0.885 1.455 1.055 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.805 0.925 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
END NAND2HD1XHT

MACRO NAND2HD2XSPGHT
  CLASS  CORE ;
  FOREIGN NAND2HD2XSPGHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 0.345 0.425 0.885 3.075 ;
      LAYER V7 ;
        RECT 0.435 0.845 0.795 1.205 ;
      LAYER M7 ;
        RECT 0.285 0.835 0.950 1.215 ;
      LAYER V6 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M4 ;
        RECT 0.515 0.780 0.715 1.600 ;
      LAYER V3 ;
        RECT 0.520 1.340 0.710 1.530 ;
      LAYER M3 ;
        RECT 0.105 1.270 0.715 1.600 ;
      LAYER V2 ;
        RECT 0.110 1.340 0.300 1.530 ;
      LAYER M2 ;
        RECT 0.105 1.190 0.305 2.070 ;
      LAYER V1 ;
        RECT 0.110 1.750 0.300 1.940 ;
      LAYER M1 ;
        RECT 0.100 1.550 0.310 2.625 ;
        RECT 0.100 1.550 1.150 1.850 ;
        RECT 2.455 1.585 2.875 1.755 ;
        RECT 2.705 1.585 2.875 2.625 ;
        RECT 0.100 2.455 2.875 2.625 ;
      LAYER M6 ;
        RECT 0.515 0.425 0.715 1.670 ;
      LAYER V5 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M5 ;
        RECT 0.285 0.925 1.015 1.125 ;
      LAYER V4 ;
        RECT 0.520 0.930 0.710 1.120 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 1.575 0.425 2.115 3.075 ;
      LAYER V7 ;
        RECT 1.665 0.845 2.025 1.205 ;
      LAYER M7 ;
        RECT 1.235 0.835 2.140 1.215 ;
      LAYER V6 ;
        RECT 1.750 0.930 1.940 1.120 ;
      LAYER M4 ;
        RECT 1.335 0.590 1.535 1.450 ;
      LAYER V3 ;
        RECT 1.340 0.930 1.530 1.120 ;
      LAYER M3 ;
        RECT 0.920 0.860 1.535 1.190 ;
      LAYER V2 ;
        RECT 1.340 0.930 1.530 1.120 ;
      LAYER M2 ;
        RECT 1.335 0.805 1.535 1.670 ;
      LAYER V1 ;
        RECT 1.340 1.340 1.530 1.530 ;
      LAYER M1 ;
        RECT 1.330 1.265 1.540 1.820 ;
        RECT 1.330 1.520 1.700 1.820 ;
      LAYER M6 ;
        RECT 1.745 0.425 1.945 1.670 ;
      LAYER V5 ;
        RECT 1.750 0.930 1.940 1.120 ;
      LAYER M5 ;
        RECT 1.235 0.925 2.240 1.125 ;
      LAYER V4 ;
        RECT 1.340 0.930 1.530 1.120 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.840 -0.300 1.010 1.120 ;
        RECT 2.700 -0.300 2.870 1.120 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 2.805 0.425 3.345 3.075 ;
      LAYER V7 ;
        RECT 2.895 1.665 3.255 2.025 ;
      LAYER M7 ;
        RECT 2.730 1.655 3.345 2.035 ;
      LAYER V6 ;
        RECT 2.980 1.750 3.170 1.940 ;
      LAYER M4 ;
        RECT 2.975 1.445 3.175 2.475 ;
      LAYER V3 ;
        RECT 2.980 2.160 3.170 2.350 ;
      LAYER M3 ;
        RECT 2.005 2.155 3.360 2.355 ;
      LAYER V2 ;
        RECT 2.160 2.160 2.350 2.350 ;
      LAYER M2 ;
        RECT 2.155 0.825 2.355 2.455 ;
      LAYER V1 ;
        RECT 2.160 0.930 2.350 1.120 ;
      LAYER M1 ;
        RECT 1.705 0.480 2.100 1.055 ;
        RECT 1.705 0.850 2.360 1.055 ;
        RECT 1.890 0.480 2.100 2.215 ;
        RECT 1.890 0.850 2.360 1.195 ;
        RECT 1.185 2.045 2.525 2.215 ;
      LAYER M6 ;
        RECT 2.975 1.155 3.175 2.460 ;
      LAYER V5 ;
        RECT 2.980 1.750 3.170 1.940 ;
      LAYER M5 ;
        RECT 2.290 1.745 3.345 1.945 ;
      LAYER V4 ;
        RECT 2.980 1.750 3.170 1.940 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.665 2.805 0.965 3.990 ;
        RECT 1.705 2.805 2.005 3.990 ;
        RECT 2.745 2.805 3.045 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
END NAND2HD2XSPGHT

MACRO NAND2HD1XSPGHT
  CLASS  CORE ;
  FOREIGN NAND2HD1XSPGHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 0.345 0.425 0.885 3.075 ;
      LAYER V7 ;
        RECT 0.435 0.845 0.795 1.205 ;
      LAYER M7 ;
        RECT 0.170 0.835 0.885 1.215 ;
      LAYER V6 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M4 ;
        RECT 0.515 0.810 0.715 1.620 ;
      LAYER V3 ;
        RECT 0.520 1.340 0.710 1.530 ;
      LAYER M3 ;
        RECT 0.105 1.250 0.850 1.620 ;
      LAYER V2 ;
        RECT 0.110 1.340 0.300 1.530 ;
      LAYER M2 ;
        RECT 0.105 1.270 0.305 2.015 ;
      LAYER V1 ;
        RECT 0.110 1.750 0.300 1.940 ;
      LAYER M1 ;
        RECT 0.100 1.520 0.310 2.015 ;
        RECT 0.100 1.520 1.585 1.820 ;
      LAYER M6 ;
        RECT 0.515 0.585 0.715 2.660 ;
      LAYER V5 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M5 ;
        RECT 0.170 0.925 1.230 1.125 ;
      LAYER V4 ;
        RECT 0.520 0.930 0.710 1.120 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 1.575 0.425 2.115 3.075 ;
      LAYER V7 ;
        RECT 1.665 0.845 2.025 1.205 ;
      LAYER M7 ;
        RECT 1.450 0.835 2.320 1.215 ;
      LAYER V6 ;
        RECT 1.750 0.930 1.940 1.120 ;
      LAYER M4 ;
        RECT 1.745 0.730 1.945 1.610 ;
      LAYER V3 ;
        RECT 1.750 0.930 1.940 1.120 ;
      LAYER M3 ;
        RECT 1.465 0.840 2.360 1.210 ;
      LAYER V2 ;
        RECT 2.160 0.930 2.350 1.120 ;
      LAYER M2 ;
        RECT 2.155 0.855 2.355 1.670 ;
      LAYER V1 ;
        RECT 2.160 1.340 2.350 1.530 ;
      LAYER M1 ;
        RECT 2.135 1.265 2.500 1.820 ;
      LAYER M6 ;
        RECT 1.745 0.585 1.945 2.660 ;
      LAYER V5 ;
        RECT 1.750 0.930 1.940 1.120 ;
      LAYER M5 ;
        RECT 1.450 0.925 2.725 1.125 ;
      LAYER V4 ;
        RECT 1.750 0.930 1.940 1.120 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.255 -0.300 1.425 1.120 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 2.805 0.425 3.345 3.075 ;
      LAYER V7 ;
        RECT 2.895 2.075 3.255 2.435 ;
      LAYER M7 ;
        RECT 2.465 2.065 3.345 2.445 ;
      LAYER V6 ;
        RECT 2.980 2.160 3.170 2.350 ;
      LAYER M4 ;
        RECT 2.565 2.070 2.765 2.830 ;
      LAYER V3 ;
        RECT 2.570 2.570 2.760 2.760 ;
      LAYER M3 ;
        RECT 2.035 2.560 2.865 2.770 ;
      LAYER V2 ;
        RECT 2.160 2.570 2.350 2.760 ;
      LAYER M2 ;
        RECT 2.155 1.980 2.355 2.870 ;
      LAYER V1 ;
        RECT 2.160 2.160 2.350 2.350 ;
      LAYER M1 ;
        RECT 1.190 2.195 1.490 2.705 ;
        RECT 1.765 0.885 1.935 2.365 ;
        RECT 1.765 2.145 2.465 2.365 ;
        RECT 1.190 2.195 2.465 2.365 ;
        RECT 2.295 2.145 2.465 2.810 ;
        RECT 2.240 0.480 2.540 1.055 ;
        RECT 1.765 0.885 2.540 1.055 ;
      LAYER M6 ;
        RECT 2.975 0.585 3.175 2.660 ;
      LAYER V5 ;
        RECT 2.980 2.160 3.170 2.350 ;
      LAYER M5 ;
        RECT 2.115 2.155 3.345 2.355 ;
      LAYER V4 ;
        RECT 2.570 2.160 2.760 2.350 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.775 2.740 1.945 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
END NAND2HD1XSPGHT

MACRO NAND2B1HDUXHT
  CLASS  CORE ;
  FOREIGN NAND2B1HDUXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.615 1.690 1.205 1.970 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.615 2.840 ;
    END
  END AN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.425 0.500 ;
        RECT 1.505 -0.300 1.705 1.070 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.455 1.125 0.755 1.430 ;
        RECT 0.455 1.250 1.960 1.430 ;
        RECT 1.515 2.090 1.960 2.420 ;
        RECT 1.775 1.250 1.960 2.420 ;
        RECT 1.145 2.170 1.960 2.420 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.620 3.030 0.920 3.990 ;
        RECT 1.145 3.030 1.445 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.680 0.275 2.320 ;
        RECT 0.105 2.060 0.405 2.320 ;
        RECT 0.105 2.150 0.965 2.320 ;
        RECT 0.795 2.150 0.965 2.770 ;
        RECT 0.705 0.480 1.005 0.875 ;
        RECT 0.105 0.680 1.005 0.875 ;
        RECT 0.795 2.600 1.815 2.770 ;
  END 
END NAND2B1HDUXHT

MACRO NAND2B1HDMXHT
  CLASS  CORE ;
  FOREIGN NAND2B1HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.830 0.920 1.485 1.130 ;
        RECT 1.315 0.920 1.485 1.820 ;
        RECT 1.315 1.520 1.560 1.820 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.495 0.520 2.835 ;
    END
  END AN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.620 -0.300 0.920 0.735 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.675 0.840 1.950 1.360 ;
        RECT 1.765 0.840 1.950 2.215 ;
        RECT 1.170 2.045 1.950 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 2.310 0.890 3.990 ;
        RECT 1.645 2.925 1.945 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.135 1.755 ;
  END 
END NAND2B1HDMXHT

MACRO NAND2B1HDLXHT
  CLASS  CORE ;
  FOREIGN NAND2B1HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.825 0.915 1.485 1.130 ;
        RECT 1.310 0.915 1.485 1.820 ;
        RECT 1.310 1.520 1.560 1.820 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 2.495 0.510 2.835 ;
    END
  END AN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.650 -0.300 0.950 0.735 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.675 0.840 1.950 1.360 ;
        RECT 1.765 0.840 1.950 2.215 ;
        RECT 1.170 2.045 1.950 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.100 0.860 3.990 ;
        RECT 1.645 2.660 1.945 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.580 1.130 1.755 ;
  END 
END NAND2B1HDLXHT

MACRO NAND2B1HD2XHT
  CLASS  CORE ;
  FOREIGN NAND2B1HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 1.240 1.545 1.820 ;
        RECT 1.330 1.520 1.820 1.820 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.495 0.475 2.980 ;
    END
  END AN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.055 ;
        RECT 2.740 -0.300 3.040 1.055 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 0.480 1.950 1.195 ;
        RECT 1.740 0.920 2.180 1.195 ;
        RECT 2.000 0.920 2.180 2.215 ;
        RECT 1.180 2.045 2.520 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.805 0.955 3.990 ;
        RECT 1.700 2.805 2.000 3.990 ;
        RECT 2.740 2.805 3.040 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.815 1.635 0.985 2.575 ;
        RECT 0.170 1.635 1.130 1.820 ;
        RECT 2.560 1.585 2.880 1.755 ;
        RECT 2.700 1.585 2.880 2.575 ;
        RECT 0.815 2.395 2.880 2.575 ;
  END 
END NAND2B1HD2XHT

MACRO MUXI4HDMXHT
  CLASS  CORE ;
  FOREIGN MUXI4HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.200 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.240 2.500 6.520 2.830 ;
        RECT 6.240 2.595 6.750 2.830 ;
    END
  END S1
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.165 1.890 4.420 2.440 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.485 1.730 2.830 2.140 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.060 0.910 2.525 1.385 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 1.200 1.230 1.665 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.665 ;
        RECT 2.375 -0.300 2.675 0.665 ;
        RECT 4.380 -0.300 4.680 0.655 ;
        RECT 5.930 -0.300 6.230 0.665 ;
        RECT 7.275 -0.300 7.445 1.210 ;
        RECT 0.000 -0.300 8.200 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.795 1.060 7.965 2.460 ;
        RECT 7.795 2.025 8.100 2.460 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.675 3.040 0.975 3.990 ;
        RECT 2.385 3.040 2.685 3.990 ;
        RECT 4.280 3.035 4.580 3.990 ;
        RECT 6.080 3.025 6.380 3.990 ;
        RECT 7.180 2.370 7.480 3.990 ;
        RECT 0.000 3.390 8.200 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.500 1.910 0.680 2.420 ;
        RECT 0.500 2.000 0.780 2.420 ;
        RECT 0.500 2.000 1.955 2.170 ;
        RECT 3.300 1.155 3.790 1.325 ;
        RECT 3.620 1.155 3.790 2.125 ;
        RECT 3.620 1.955 3.920 2.125 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.105 1.075 0.275 2.860 ;
        RECT 0.105 1.075 0.405 1.245 ;
        RECT 0.105 2.600 0.405 2.860 ;
        RECT 1.165 2.690 1.335 3.030 ;
        RECT 0.105 2.690 1.335 2.860 ;
        RECT 1.165 2.860 2.045 3.030 ;
        RECT 2.305 2.690 2.765 2.860 ;
        RECT 3.030 2.865 3.035 3.210 ;
        RECT 3.030 3.040 3.325 3.210 ;
        RECT 2.865 2.710 2.875 3.210 ;
        RECT 2.875 2.720 2.885 3.210 ;
        RECT 2.885 2.730 2.895 3.210 ;
        RECT 2.895 2.740 2.905 3.210 ;
        RECT 2.905 2.750 2.915 3.210 ;
        RECT 2.915 2.760 2.925 3.210 ;
        RECT 2.925 2.770 2.935 3.210 ;
        RECT 2.935 2.780 2.945 3.210 ;
        RECT 2.945 2.790 2.955 3.210 ;
        RECT 2.955 2.800 2.965 3.210 ;
        RECT 2.965 2.810 2.975 3.210 ;
        RECT 2.975 2.820 2.985 3.210 ;
        RECT 2.985 2.830 2.995 3.210 ;
        RECT 2.995 2.840 3.005 3.210 ;
        RECT 3.005 2.850 3.015 3.210 ;
        RECT 3.015 2.860 3.025 3.210 ;
        RECT 3.025 2.865 3.031 3.209 ;
        RECT 2.855 2.700 2.865 2.950 ;
        RECT 2.765 2.690 2.775 2.860 ;
        RECT 2.775 2.690 2.785 2.870 ;
        RECT 2.785 2.690 2.795 2.880 ;
        RECT 2.795 2.690 2.805 2.890 ;
        RECT 2.805 2.690 2.815 2.900 ;
        RECT 2.815 2.690 2.825 2.910 ;
        RECT 2.825 2.690 2.835 2.920 ;
        RECT 2.835 2.690 2.845 2.930 ;
        RECT 2.845 2.690 2.855 2.940 ;
        RECT 2.215 2.690 2.225 2.940 ;
        RECT 2.225 2.690 2.235 2.930 ;
        RECT 2.235 2.690 2.245 2.920 ;
        RECT 2.245 2.690 2.255 2.910 ;
        RECT 2.255 2.690 2.265 2.900 ;
        RECT 2.265 2.690 2.275 2.890 ;
        RECT 2.275 2.690 2.285 2.880 ;
        RECT 2.285 2.690 2.295 2.870 ;
        RECT 2.295 2.690 2.305 2.860 ;
        RECT 2.135 2.770 2.145 3.020 ;
        RECT 2.145 2.760 2.155 3.010 ;
        RECT 2.155 2.750 2.165 3.000 ;
        RECT 2.165 2.740 2.175 2.990 ;
        RECT 2.175 2.730 2.185 2.980 ;
        RECT 2.185 2.720 2.195 2.970 ;
        RECT 2.195 2.710 2.205 2.960 ;
        RECT 2.205 2.700 2.215 2.950 ;
        RECT 2.045 2.860 2.055 3.030 ;
        RECT 2.055 2.850 2.065 3.030 ;
        RECT 2.065 2.840 2.075 3.030 ;
        RECT 2.075 2.830 2.085 3.030 ;
        RECT 2.085 2.820 2.095 3.030 ;
        RECT 2.095 2.810 2.105 3.030 ;
        RECT 2.105 2.800 2.115 3.030 ;
        RECT 2.115 2.790 2.125 3.030 ;
        RECT 2.125 2.780 2.135 3.030 ;
        RECT 3.220 1.505 3.270 1.675 ;
        RECT 3.530 2.325 3.740 2.495 ;
        RECT 3.120 0.785 4.140 0.955 ;
        RECT 3.970 0.785 4.140 1.325 ;
        RECT 3.970 1.155 4.785 1.325 ;
        RECT 4.615 1.155 4.785 1.780 ;
        RECT 3.440 2.245 3.450 2.495 ;
        RECT 3.450 2.255 3.460 2.495 ;
        RECT 3.460 2.265 3.470 2.495 ;
        RECT 3.470 2.275 3.480 2.495 ;
        RECT 3.480 2.285 3.490 2.495 ;
        RECT 3.490 2.295 3.500 2.495 ;
        RECT 3.500 2.305 3.510 2.495 ;
        RECT 3.510 2.315 3.520 2.495 ;
        RECT 3.520 2.325 3.530 2.495 ;
        RECT 3.270 1.505 3.280 2.325 ;
        RECT 3.280 1.505 3.290 2.335 ;
        RECT 3.290 1.505 3.300 2.345 ;
        RECT 3.300 1.505 3.310 2.355 ;
        RECT 3.310 1.505 3.320 2.365 ;
        RECT 3.320 1.505 3.330 2.375 ;
        RECT 3.330 1.505 3.340 2.385 ;
        RECT 3.340 1.505 3.350 2.395 ;
        RECT 3.350 1.505 3.360 2.405 ;
        RECT 3.360 1.505 3.370 2.415 ;
        RECT 3.370 1.505 3.380 2.425 ;
        RECT 3.380 1.505 3.390 2.435 ;
        RECT 3.390 1.505 3.400 2.445 ;
        RECT 3.400 1.505 3.410 2.455 ;
        RECT 3.410 1.505 3.420 2.465 ;
        RECT 3.420 1.505 3.430 2.475 ;
        RECT 3.430 1.505 3.440 2.485 ;
        RECT 3.130 1.425 3.140 1.675 ;
        RECT 3.140 1.435 3.150 1.675 ;
        RECT 3.150 1.445 3.160 1.675 ;
        RECT 3.160 1.455 3.170 1.675 ;
        RECT 3.170 1.465 3.180 1.675 ;
        RECT 3.180 1.475 3.190 1.675 ;
        RECT 3.190 1.485 3.200 1.675 ;
        RECT 3.200 1.495 3.210 1.675 ;
        RECT 3.210 1.505 3.220 1.675 ;
        RECT 3.120 1.415 3.130 1.665 ;
        RECT 2.950 0.785 2.960 1.495 ;
        RECT 2.960 0.785 2.970 1.505 ;
        RECT 2.970 0.785 2.980 1.515 ;
        RECT 2.980 0.785 2.990 1.525 ;
        RECT 2.990 0.785 3.000 1.535 ;
        RECT 3.000 0.785 3.010 1.545 ;
        RECT 3.010 0.785 3.020 1.555 ;
        RECT 3.020 0.785 3.030 1.565 ;
        RECT 3.030 0.785 3.040 1.575 ;
        RECT 3.040 0.785 3.050 1.585 ;
        RECT 3.050 0.785 3.060 1.595 ;
        RECT 3.060 0.785 3.070 1.605 ;
        RECT 3.070 0.785 3.080 1.615 ;
        RECT 3.080 0.785 3.090 1.625 ;
        RECT 3.090 0.785 3.100 1.635 ;
        RECT 3.100 0.785 3.110 1.645 ;
        RECT 3.110 0.785 3.120 1.655 ;
        RECT 1.520 0.720 1.690 1.820 ;
        RECT 1.515 2.370 2.015 2.540 ;
        RECT 2.045 2.340 2.105 2.540 ;
        RECT 1.520 1.650 2.305 1.820 ;
        RECT 2.135 1.650 2.305 2.510 ;
        RECT 2.135 2.340 2.935 2.510 ;
        RECT 3.360 2.675 5.700 2.855 ;
        RECT 6.105 1.610 6.165 2.190 ;
        RECT 5.995 1.610 6.005 2.290 ;
        RECT 6.005 1.610 6.015 2.280 ;
        RECT 6.015 1.610 6.025 2.270 ;
        RECT 6.025 1.610 6.035 2.260 ;
        RECT 6.035 1.610 6.045 2.250 ;
        RECT 6.045 1.610 6.055 2.240 ;
        RECT 6.055 1.610 6.065 2.230 ;
        RECT 6.065 1.610 6.075 2.220 ;
        RECT 6.075 1.610 6.085 2.210 ;
        RECT 6.085 1.610 6.095 2.200 ;
        RECT 6.095 1.610 6.105 2.190 ;
        RECT 5.825 2.210 5.835 2.800 ;
        RECT 5.835 2.200 5.845 2.790 ;
        RECT 5.845 2.190 5.855 2.780 ;
        RECT 5.855 2.180 5.865 2.770 ;
        RECT 5.865 2.170 5.875 2.760 ;
        RECT 5.875 2.160 5.885 2.750 ;
        RECT 5.885 2.150 5.895 2.740 ;
        RECT 5.895 2.140 5.905 2.730 ;
        RECT 5.905 2.130 5.915 2.720 ;
        RECT 5.915 2.120 5.925 2.710 ;
        RECT 5.925 2.110 5.935 2.700 ;
        RECT 5.935 2.100 5.945 2.690 ;
        RECT 5.945 2.090 5.955 2.680 ;
        RECT 5.955 2.080 5.965 2.670 ;
        RECT 5.965 2.070 5.975 2.660 ;
        RECT 5.975 2.060 5.985 2.650 ;
        RECT 5.985 2.050 5.995 2.640 ;
        RECT 5.780 2.595 5.790 2.845 ;
        RECT 5.790 2.585 5.800 2.835 ;
        RECT 5.800 2.575 5.810 2.825 ;
        RECT 5.810 2.565 5.820 2.815 ;
        RECT 5.820 2.555 5.826 2.809 ;
        RECT 5.700 2.675 5.710 2.855 ;
        RECT 5.710 2.665 5.720 2.855 ;
        RECT 5.720 2.655 5.730 2.855 ;
        RECT 5.730 2.645 5.740 2.855 ;
        RECT 5.740 2.635 5.750 2.855 ;
        RECT 5.750 2.625 5.760 2.855 ;
        RECT 5.760 2.615 5.770 2.855 ;
        RECT 5.770 2.605 5.780 2.855 ;
        RECT 3.280 2.605 3.290 2.855 ;
        RECT 3.290 2.615 3.300 2.855 ;
        RECT 3.300 2.625 3.310 2.855 ;
        RECT 3.310 2.635 3.320 2.855 ;
        RECT 3.320 2.645 3.330 2.855 ;
        RECT 3.330 2.655 3.340 2.855 ;
        RECT 3.340 2.665 3.350 2.855 ;
        RECT 3.350 2.675 3.360 2.855 ;
        RECT 3.025 2.350 3.035 2.600 ;
        RECT 3.035 2.360 3.045 2.610 ;
        RECT 3.045 2.370 3.055 2.620 ;
        RECT 3.055 2.380 3.065 2.630 ;
        RECT 3.065 2.390 3.075 2.640 ;
        RECT 3.075 2.400 3.085 2.650 ;
        RECT 3.085 2.410 3.095 2.660 ;
        RECT 3.095 2.420 3.105 2.670 ;
        RECT 3.105 2.430 3.115 2.680 ;
        RECT 3.115 2.440 3.125 2.690 ;
        RECT 3.125 2.450 3.135 2.700 ;
        RECT 3.135 2.460 3.145 2.710 ;
        RECT 3.145 2.470 3.155 2.720 ;
        RECT 3.155 2.480 3.165 2.730 ;
        RECT 3.165 2.490 3.175 2.740 ;
        RECT 3.175 2.500 3.185 2.750 ;
        RECT 3.185 2.510 3.195 2.760 ;
        RECT 3.195 2.520 3.205 2.770 ;
        RECT 3.205 2.530 3.215 2.780 ;
        RECT 3.215 2.540 3.225 2.790 ;
        RECT 3.225 2.550 3.235 2.800 ;
        RECT 3.235 2.560 3.245 2.810 ;
        RECT 3.245 2.570 3.255 2.820 ;
        RECT 3.255 2.580 3.265 2.830 ;
        RECT 3.265 2.590 3.275 2.840 ;
        RECT 3.275 2.595 3.281 2.849 ;
        RECT 2.935 2.340 2.945 2.510 ;
        RECT 2.945 2.340 2.955 2.520 ;
        RECT 2.955 2.340 2.965 2.530 ;
        RECT 2.965 2.340 2.975 2.540 ;
        RECT 2.975 2.340 2.985 2.550 ;
        RECT 2.985 2.340 2.995 2.560 ;
        RECT 2.995 2.340 3.005 2.570 ;
        RECT 3.005 2.340 3.015 2.580 ;
        RECT 3.015 2.340 3.025 2.590 ;
        RECT 2.105 2.340 2.115 2.530 ;
        RECT 2.115 2.340 2.125 2.520 ;
        RECT 2.125 2.340 2.135 2.510 ;
        RECT 2.015 2.370 2.025 2.540 ;
        RECT 2.025 2.360 2.035 2.540 ;
        RECT 2.035 2.350 2.045 2.540 ;
        RECT 5.620 1.815 5.700 2.015 ;
        RECT 5.610 1.825 5.806 1.889 ;
        RECT 5.630 1.805 5.700 2.015 ;
        RECT 5.600 1.835 5.806 1.889 ;
        RECT 5.400 1.845 5.700 2.015 ;
        RECT 5.400 1.845 5.710 1.985 ;
        RECT 5.400 1.845 5.720 1.975 ;
        RECT 5.400 1.845 5.730 1.965 ;
        RECT 5.400 1.845 5.740 1.955 ;
        RECT 5.400 1.845 5.750 1.945 ;
        RECT 5.400 1.845 5.760 1.935 ;
        RECT 5.400 1.845 5.770 1.925 ;
        RECT 5.400 1.845 5.780 1.915 ;
        RECT 5.400 1.845 5.790 1.905 ;
        RECT 5.400 1.845 5.800 1.895 ;
        RECT 5.635 1.255 5.806 1.889 ;
        RECT 5.635 1.255 6.865 1.425 ;
        RECT 6.695 1.040 6.865 2.340 ;
        RECT 4.965 1.170 5.135 2.495 ;
        RECT 5.285 0.905 5.455 1.340 ;
        RECT 4.965 1.170 5.455 1.340 ;
        RECT 4.965 2.325 5.520 2.495 ;
        RECT 5.285 0.905 6.310 1.075 ;
        RECT 6.615 0.690 7.095 0.860 ;
        RECT 6.525 0.690 6.535 0.940 ;
        RECT 6.535 0.690 6.545 0.930 ;
        RECT 6.545 0.690 6.555 0.920 ;
        RECT 6.555 0.690 6.565 0.910 ;
        RECT 6.565 0.690 6.575 0.900 ;
        RECT 6.575 0.690 6.585 0.890 ;
        RECT 6.585 0.690 6.595 0.880 ;
        RECT 6.595 0.690 6.605 0.870 ;
        RECT 6.605 0.690 6.615 0.860 ;
        RECT 6.400 0.815 6.410 1.065 ;
        RECT 6.410 0.805 6.420 1.055 ;
        RECT 6.420 0.795 6.430 1.045 ;
        RECT 6.430 0.785 6.440 1.035 ;
        RECT 6.440 0.775 6.450 1.025 ;
        RECT 6.450 0.765 6.460 1.015 ;
        RECT 6.460 0.755 6.470 1.005 ;
        RECT 6.470 0.745 6.480 0.995 ;
        RECT 6.480 0.735 6.490 0.985 ;
        RECT 6.490 0.725 6.500 0.975 ;
        RECT 6.500 0.715 6.510 0.965 ;
        RECT 6.510 0.705 6.520 0.955 ;
        RECT 6.520 0.695 6.526 0.949 ;
        RECT 6.310 0.905 6.320 1.075 ;
        RECT 6.320 0.895 6.330 1.075 ;
        RECT 6.330 0.885 6.340 1.075 ;
        RECT 6.340 0.875 6.350 1.075 ;
        RECT 6.350 0.865 6.360 1.075 ;
        RECT 6.360 0.855 6.370 1.075 ;
        RECT 6.370 0.845 6.380 1.075 ;
        RECT 6.380 0.835 6.390 1.075 ;
        RECT 6.390 0.825 6.400 1.075 ;
  END 
END MUXI4HDMXHT

MACRO MUXI4HDLXHT
  CLASS  CORE ;
  FOREIGN MUXI4HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.200 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.240 2.500 6.525 2.830 ;
        RECT 6.240 2.565 6.750 2.830 ;
    END
  END S1
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.165 1.890 4.420 2.440 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.485 1.730 2.830 2.140 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.060 0.910 2.525 1.385 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 1.200 1.230 1.665 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.665 ;
        RECT 2.375 -0.300 2.675 0.665 ;
        RECT 4.380 -0.300 4.680 0.655 ;
        RECT 5.930 -0.300 6.230 0.665 ;
        RECT 7.275 -0.300 7.445 1.360 ;
        RECT 0.000 -0.300 8.200 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.795 1.060 7.965 2.460 ;
        RECT 7.795 2.055 8.100 2.460 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.675 3.040 0.975 3.990 ;
        RECT 2.385 3.040 2.685 3.990 ;
        RECT 4.280 3.035 4.580 3.990 ;
        RECT 6.080 3.025 6.380 3.990 ;
        RECT 7.180 2.165 7.480 3.990 ;
        RECT 0.000 3.390 8.200 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.500 1.910 0.680 2.420 ;
        RECT 0.500 2.000 0.780 2.420 ;
        RECT 0.500 2.000 1.955 2.170 ;
        RECT 3.300 1.155 3.790 1.325 ;
        RECT 3.620 1.155 3.790 2.125 ;
        RECT 3.620 1.955 3.920 2.125 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.105 1.075 0.275 2.860 ;
        RECT 0.105 1.075 0.405 1.245 ;
        RECT 0.105 2.600 0.405 2.860 ;
        RECT 1.165 2.690 1.335 3.030 ;
        RECT 0.105 2.690 1.335 2.860 ;
        RECT 1.165 2.860 2.045 3.030 ;
        RECT 2.305 2.690 2.765 2.860 ;
        RECT 3.030 2.865 3.035 3.210 ;
        RECT 3.030 3.040 3.325 3.210 ;
        RECT 2.865 2.710 2.875 3.210 ;
        RECT 2.875 2.720 2.885 3.210 ;
        RECT 2.885 2.730 2.895 3.210 ;
        RECT 2.895 2.740 2.905 3.210 ;
        RECT 2.905 2.750 2.915 3.210 ;
        RECT 2.915 2.760 2.925 3.210 ;
        RECT 2.925 2.770 2.935 3.210 ;
        RECT 2.935 2.780 2.945 3.210 ;
        RECT 2.945 2.790 2.955 3.210 ;
        RECT 2.955 2.800 2.965 3.210 ;
        RECT 2.965 2.810 2.975 3.210 ;
        RECT 2.975 2.820 2.985 3.210 ;
        RECT 2.985 2.830 2.995 3.210 ;
        RECT 2.995 2.840 3.005 3.210 ;
        RECT 3.005 2.850 3.015 3.210 ;
        RECT 3.015 2.860 3.025 3.210 ;
        RECT 3.025 2.865 3.031 3.209 ;
        RECT 2.855 2.700 2.865 2.950 ;
        RECT 2.765 2.690 2.775 2.860 ;
        RECT 2.775 2.690 2.785 2.870 ;
        RECT 2.785 2.690 2.795 2.880 ;
        RECT 2.795 2.690 2.805 2.890 ;
        RECT 2.805 2.690 2.815 2.900 ;
        RECT 2.815 2.690 2.825 2.910 ;
        RECT 2.825 2.690 2.835 2.920 ;
        RECT 2.835 2.690 2.845 2.930 ;
        RECT 2.845 2.690 2.855 2.940 ;
        RECT 2.215 2.690 2.225 2.940 ;
        RECT 2.225 2.690 2.235 2.930 ;
        RECT 2.235 2.690 2.245 2.920 ;
        RECT 2.245 2.690 2.255 2.910 ;
        RECT 2.255 2.690 2.265 2.900 ;
        RECT 2.265 2.690 2.275 2.890 ;
        RECT 2.275 2.690 2.285 2.880 ;
        RECT 2.285 2.690 2.295 2.870 ;
        RECT 2.295 2.690 2.305 2.860 ;
        RECT 2.135 2.770 2.145 3.020 ;
        RECT 2.145 2.760 2.155 3.010 ;
        RECT 2.155 2.750 2.165 3.000 ;
        RECT 2.165 2.740 2.175 2.990 ;
        RECT 2.175 2.730 2.185 2.980 ;
        RECT 2.185 2.720 2.195 2.970 ;
        RECT 2.195 2.710 2.205 2.960 ;
        RECT 2.205 2.700 2.215 2.950 ;
        RECT 2.045 2.860 2.055 3.030 ;
        RECT 2.055 2.850 2.065 3.030 ;
        RECT 2.065 2.840 2.075 3.030 ;
        RECT 2.075 2.830 2.085 3.030 ;
        RECT 2.085 2.820 2.095 3.030 ;
        RECT 2.095 2.810 2.105 3.030 ;
        RECT 2.105 2.800 2.115 3.030 ;
        RECT 2.115 2.790 2.125 3.030 ;
        RECT 2.125 2.780 2.135 3.030 ;
        RECT 3.220 1.505 3.270 1.675 ;
        RECT 3.530 2.325 3.740 2.495 ;
        RECT 3.120 0.785 4.140 0.955 ;
        RECT 3.970 0.785 4.140 1.325 ;
        RECT 3.970 1.155 4.785 1.325 ;
        RECT 4.615 1.155 4.785 1.780 ;
        RECT 3.440 2.245 3.450 2.495 ;
        RECT 3.450 2.255 3.460 2.495 ;
        RECT 3.460 2.265 3.470 2.495 ;
        RECT 3.470 2.275 3.480 2.495 ;
        RECT 3.480 2.285 3.490 2.495 ;
        RECT 3.490 2.295 3.500 2.495 ;
        RECT 3.500 2.305 3.510 2.495 ;
        RECT 3.510 2.315 3.520 2.495 ;
        RECT 3.520 2.325 3.530 2.495 ;
        RECT 3.270 1.505 3.280 2.325 ;
        RECT 3.280 1.505 3.290 2.335 ;
        RECT 3.290 1.505 3.300 2.345 ;
        RECT 3.300 1.505 3.310 2.355 ;
        RECT 3.310 1.505 3.320 2.365 ;
        RECT 3.320 1.505 3.330 2.375 ;
        RECT 3.330 1.505 3.340 2.385 ;
        RECT 3.340 1.505 3.350 2.395 ;
        RECT 3.350 1.505 3.360 2.405 ;
        RECT 3.360 1.505 3.370 2.415 ;
        RECT 3.370 1.505 3.380 2.425 ;
        RECT 3.380 1.505 3.390 2.435 ;
        RECT 3.390 1.505 3.400 2.445 ;
        RECT 3.400 1.505 3.410 2.455 ;
        RECT 3.410 1.505 3.420 2.465 ;
        RECT 3.420 1.505 3.430 2.475 ;
        RECT 3.430 1.505 3.440 2.485 ;
        RECT 3.130 1.425 3.140 1.675 ;
        RECT 3.140 1.435 3.150 1.675 ;
        RECT 3.150 1.445 3.160 1.675 ;
        RECT 3.160 1.455 3.170 1.675 ;
        RECT 3.170 1.465 3.180 1.675 ;
        RECT 3.180 1.475 3.190 1.675 ;
        RECT 3.190 1.485 3.200 1.675 ;
        RECT 3.200 1.495 3.210 1.675 ;
        RECT 3.210 1.505 3.220 1.675 ;
        RECT 3.120 1.415 3.130 1.665 ;
        RECT 2.950 0.785 2.960 1.495 ;
        RECT 2.960 0.785 2.970 1.505 ;
        RECT 2.970 0.785 2.980 1.515 ;
        RECT 2.980 0.785 2.990 1.525 ;
        RECT 2.990 0.785 3.000 1.535 ;
        RECT 3.000 0.785 3.010 1.545 ;
        RECT 3.010 0.785 3.020 1.555 ;
        RECT 3.020 0.785 3.030 1.565 ;
        RECT 3.030 0.785 3.040 1.575 ;
        RECT 3.040 0.785 3.050 1.585 ;
        RECT 3.050 0.785 3.060 1.595 ;
        RECT 3.060 0.785 3.070 1.605 ;
        RECT 3.070 0.785 3.080 1.615 ;
        RECT 3.080 0.785 3.090 1.625 ;
        RECT 3.090 0.785 3.100 1.635 ;
        RECT 3.100 0.785 3.110 1.645 ;
        RECT 3.110 0.785 3.120 1.655 ;
        RECT 1.520 0.720 1.690 1.820 ;
        RECT 1.515 2.370 2.015 2.540 ;
        RECT 2.045 2.340 2.105 2.540 ;
        RECT 1.520 1.650 2.305 1.820 ;
        RECT 2.135 1.650 2.305 2.510 ;
        RECT 2.135 2.340 2.935 2.510 ;
        RECT 3.360 2.675 5.715 2.855 ;
        RECT 6.105 1.610 6.165 2.190 ;
        RECT 5.995 1.610 6.005 2.290 ;
        RECT 6.005 1.610 6.015 2.280 ;
        RECT 6.015 1.610 6.025 2.270 ;
        RECT 6.025 1.610 6.035 2.260 ;
        RECT 6.035 1.610 6.045 2.250 ;
        RECT 6.045 1.610 6.055 2.240 ;
        RECT 6.055 1.610 6.065 2.230 ;
        RECT 6.065 1.610 6.075 2.220 ;
        RECT 6.075 1.610 6.085 2.210 ;
        RECT 6.085 1.610 6.095 2.200 ;
        RECT 6.095 1.610 6.105 2.190 ;
        RECT 5.825 2.210 5.835 2.800 ;
        RECT 5.835 2.200 5.845 2.790 ;
        RECT 5.845 2.190 5.855 2.780 ;
        RECT 5.855 2.180 5.865 2.770 ;
        RECT 5.865 2.170 5.875 2.760 ;
        RECT 5.875 2.160 5.885 2.750 ;
        RECT 5.885 2.150 5.895 2.740 ;
        RECT 5.895 2.140 5.905 2.730 ;
        RECT 5.905 2.130 5.915 2.720 ;
        RECT 5.915 2.120 5.925 2.710 ;
        RECT 5.925 2.110 5.935 2.700 ;
        RECT 5.935 2.100 5.945 2.690 ;
        RECT 5.945 2.090 5.955 2.680 ;
        RECT 5.955 2.080 5.965 2.670 ;
        RECT 5.965 2.070 5.975 2.660 ;
        RECT 5.975 2.060 5.985 2.650 ;
        RECT 5.985 2.050 5.995 2.640 ;
        RECT 5.780 2.610 5.790 2.844 ;
        RECT 5.790 2.600 5.800 2.834 ;
        RECT 5.800 2.590 5.810 2.824 ;
        RECT 5.810 2.580 5.820 2.814 ;
        RECT 5.820 2.570 5.826 2.810 ;
        RECT 5.715 2.675 5.725 2.855 ;
        RECT 5.725 2.665 5.735 2.855 ;
        RECT 5.735 2.655 5.745 2.855 ;
        RECT 5.745 2.645 5.755 2.855 ;
        RECT 5.755 2.635 5.765 2.855 ;
        RECT 5.765 2.625 5.775 2.855 ;
        RECT 5.775 2.615 5.781 2.855 ;
        RECT 3.280 2.605 3.290 2.855 ;
        RECT 3.290 2.615 3.300 2.855 ;
        RECT 3.300 2.625 3.310 2.855 ;
        RECT 3.310 2.635 3.320 2.855 ;
        RECT 3.320 2.645 3.330 2.855 ;
        RECT 3.330 2.655 3.340 2.855 ;
        RECT 3.340 2.665 3.350 2.855 ;
        RECT 3.350 2.675 3.360 2.855 ;
        RECT 3.025 2.350 3.035 2.600 ;
        RECT 3.035 2.360 3.045 2.610 ;
        RECT 3.045 2.370 3.055 2.620 ;
        RECT 3.055 2.380 3.065 2.630 ;
        RECT 3.065 2.390 3.075 2.640 ;
        RECT 3.075 2.400 3.085 2.650 ;
        RECT 3.085 2.410 3.095 2.660 ;
        RECT 3.095 2.420 3.105 2.670 ;
        RECT 3.105 2.430 3.115 2.680 ;
        RECT 3.115 2.440 3.125 2.690 ;
        RECT 3.125 2.450 3.135 2.700 ;
        RECT 3.135 2.460 3.145 2.710 ;
        RECT 3.145 2.470 3.155 2.720 ;
        RECT 3.155 2.480 3.165 2.730 ;
        RECT 3.165 2.490 3.175 2.740 ;
        RECT 3.175 2.500 3.185 2.750 ;
        RECT 3.185 2.510 3.195 2.760 ;
        RECT 3.195 2.520 3.205 2.770 ;
        RECT 3.205 2.530 3.215 2.780 ;
        RECT 3.215 2.540 3.225 2.790 ;
        RECT 3.225 2.550 3.235 2.800 ;
        RECT 3.235 2.560 3.245 2.810 ;
        RECT 3.245 2.570 3.255 2.820 ;
        RECT 3.255 2.580 3.265 2.830 ;
        RECT 3.265 2.590 3.275 2.840 ;
        RECT 3.275 2.595 3.281 2.849 ;
        RECT 2.935 2.340 2.945 2.510 ;
        RECT 2.945 2.340 2.955 2.520 ;
        RECT 2.955 2.340 2.965 2.530 ;
        RECT 2.965 2.340 2.975 2.540 ;
        RECT 2.975 2.340 2.985 2.550 ;
        RECT 2.985 2.340 2.995 2.560 ;
        RECT 2.995 2.340 3.005 2.570 ;
        RECT 3.005 2.340 3.015 2.580 ;
        RECT 3.015 2.340 3.025 2.590 ;
        RECT 2.105 2.340 2.115 2.530 ;
        RECT 2.115 2.340 2.125 2.520 ;
        RECT 2.125 2.340 2.135 2.510 ;
        RECT 2.015 2.370 2.025 2.540 ;
        RECT 2.025 2.360 2.035 2.540 ;
        RECT 2.035 2.350 2.045 2.540 ;
        RECT 5.620 1.735 5.700 1.935 ;
        RECT 5.610 1.745 5.806 1.809 ;
        RECT 5.630 1.725 5.700 1.935 ;
        RECT 5.600 1.755 5.806 1.809 ;
        RECT 5.400 1.765 5.700 1.935 ;
        RECT 5.400 1.765 5.710 1.905 ;
        RECT 5.400 1.765 5.720 1.895 ;
        RECT 5.400 1.765 5.730 1.885 ;
        RECT 5.400 1.765 5.740 1.875 ;
        RECT 5.400 1.765 5.750 1.865 ;
        RECT 5.400 1.765 5.760 1.855 ;
        RECT 5.400 1.765 5.770 1.845 ;
        RECT 5.400 1.765 5.780 1.835 ;
        RECT 5.400 1.765 5.790 1.825 ;
        RECT 5.400 1.765 5.800 1.815 ;
        RECT 5.635 1.255 5.806 1.809 ;
        RECT 5.635 1.255 6.865 1.425 ;
        RECT 6.695 1.040 6.865 2.340 ;
        RECT 4.965 1.170 5.135 2.495 ;
        RECT 5.285 0.905 5.455 1.340 ;
        RECT 4.965 1.170 5.455 1.340 ;
        RECT 4.965 2.325 5.520 2.495 ;
        RECT 5.285 0.905 6.310 1.075 ;
        RECT 6.615 0.690 7.095 0.860 ;
        RECT 6.525 0.690 6.535 0.940 ;
        RECT 6.535 0.690 6.545 0.930 ;
        RECT 6.545 0.690 6.555 0.920 ;
        RECT 6.555 0.690 6.565 0.910 ;
        RECT 6.565 0.690 6.575 0.900 ;
        RECT 6.575 0.690 6.585 0.890 ;
        RECT 6.585 0.690 6.595 0.880 ;
        RECT 6.595 0.690 6.605 0.870 ;
        RECT 6.605 0.690 6.615 0.860 ;
        RECT 6.400 0.815 6.410 1.065 ;
        RECT 6.410 0.805 6.420 1.055 ;
        RECT 6.420 0.795 6.430 1.045 ;
        RECT 6.430 0.785 6.440 1.035 ;
        RECT 6.440 0.775 6.450 1.025 ;
        RECT 6.450 0.765 6.460 1.015 ;
        RECT 6.460 0.755 6.470 1.005 ;
        RECT 6.470 0.745 6.480 0.995 ;
        RECT 6.480 0.735 6.490 0.985 ;
        RECT 6.490 0.725 6.500 0.975 ;
        RECT 6.500 0.715 6.510 0.965 ;
        RECT 6.510 0.705 6.520 0.955 ;
        RECT 6.520 0.695 6.526 0.949 ;
        RECT 6.310 0.905 6.320 1.075 ;
        RECT 6.320 0.895 6.330 1.075 ;
        RECT 6.330 0.885 6.340 1.075 ;
        RECT 6.340 0.875 6.350 1.075 ;
        RECT 6.350 0.865 6.360 1.075 ;
        RECT 6.360 0.855 6.370 1.075 ;
        RECT 6.370 0.845 6.380 1.075 ;
        RECT 6.380 0.835 6.390 1.075 ;
        RECT 6.390 0.825 6.400 1.075 ;
  END 
END MUXI4HDLXHT

MACRO MUXI4HD2XHT
  CLASS  CORE ;
  FOREIGN MUXI4HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.430 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.235 1.415 7.070 1.510 ;
        RECT 6.130 1.540 7.165 1.585 ;
        RECT 5.235 1.340 5.405 1.980 ;
        RECT 6.130 1.340 6.365 1.585 ;
        RECT 5.235 1.340 6.365 1.510 ;
        RECT 6.600 1.320 7.070 1.585 ;
        RECT 6.885 1.320 7.070 1.840 ;
        RECT 6.130 1.415 7.070 1.585 ;
        RECT 6.885 1.540 7.165 1.840 ;
    END
  END S1
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.165 1.890 4.420 2.440 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.485 1.730 2.830 2.140 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.060 0.920 2.465 1.130 ;
        RECT 2.165 0.920 2.465 1.385 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 1.200 1.230 1.630 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.665 ;
        RECT 2.375 -0.300 2.675 0.740 ;
        RECT 4.360 -0.300 4.660 1.055 ;
        RECT 6.820 -0.300 7.120 0.635 ;
        RECT 7.895 -0.300 8.065 1.120 ;
        RECT 8.870 -0.300 9.170 1.055 ;
        RECT 0.000 -0.300 9.430 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.200 2.120 8.585 2.415 ;
        RECT 8.415 0.720 8.585 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.675 3.040 0.975 3.990 ;
        RECT 2.335 3.040 2.635 3.990 ;
        RECT 4.280 3.095 4.580 3.990 ;
        RECT 6.790 2.975 7.090 3.990 ;
        RECT 7.830 2.635 8.130 3.990 ;
        RECT 8.870 2.295 9.170 3.990 ;
        RECT 0.000 3.390 9.430 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.455 1.840 0.625 2.420 ;
        RECT 0.455 1.910 0.780 2.420 ;
        RECT 0.455 1.910 1.955 2.080 ;
        RECT 3.300 1.155 3.790 1.325 ;
        RECT 3.620 1.155 3.790 2.125 ;
        RECT 3.620 1.955 3.920 2.125 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.105 1.075 0.275 2.860 ;
        RECT 0.105 1.075 0.405 1.245 ;
        RECT 0.105 2.600 0.405 2.860 ;
        RECT 1.165 2.690 1.335 3.030 ;
        RECT 0.105 2.690 1.335 2.860 ;
        RECT 1.165 2.860 1.995 3.030 ;
        RECT 2.255 2.690 2.765 2.860 ;
        RECT 3.030 2.865 3.035 3.210 ;
        RECT 3.030 3.040 3.325 3.210 ;
        RECT 2.865 2.710 2.875 3.210 ;
        RECT 2.875 2.720 2.885 3.210 ;
        RECT 2.885 2.730 2.895 3.210 ;
        RECT 2.895 2.740 2.905 3.210 ;
        RECT 2.905 2.750 2.915 3.210 ;
        RECT 2.915 2.760 2.925 3.210 ;
        RECT 2.925 2.770 2.935 3.210 ;
        RECT 2.935 2.780 2.945 3.210 ;
        RECT 2.945 2.790 2.955 3.210 ;
        RECT 2.955 2.800 2.965 3.210 ;
        RECT 2.965 2.810 2.975 3.210 ;
        RECT 2.975 2.820 2.985 3.210 ;
        RECT 2.985 2.830 2.995 3.210 ;
        RECT 2.995 2.840 3.005 3.210 ;
        RECT 3.005 2.850 3.015 3.210 ;
        RECT 3.015 2.860 3.025 3.210 ;
        RECT 3.025 2.865 3.031 3.209 ;
        RECT 2.855 2.700 2.865 2.950 ;
        RECT 2.765 2.690 2.775 2.860 ;
        RECT 2.775 2.690 2.785 2.870 ;
        RECT 2.785 2.690 2.795 2.880 ;
        RECT 2.795 2.690 2.805 2.890 ;
        RECT 2.805 2.690 2.815 2.900 ;
        RECT 2.815 2.690 2.825 2.910 ;
        RECT 2.825 2.690 2.835 2.920 ;
        RECT 2.835 2.690 2.845 2.930 ;
        RECT 2.845 2.690 2.855 2.940 ;
        RECT 2.165 2.690 2.175 2.940 ;
        RECT 2.175 2.690 2.185 2.930 ;
        RECT 2.185 2.690 2.195 2.920 ;
        RECT 2.195 2.690 2.205 2.910 ;
        RECT 2.205 2.690 2.215 2.900 ;
        RECT 2.215 2.690 2.225 2.890 ;
        RECT 2.225 2.690 2.235 2.880 ;
        RECT 2.235 2.690 2.245 2.870 ;
        RECT 2.245 2.690 2.255 2.860 ;
        RECT 2.085 2.770 2.095 3.020 ;
        RECT 2.095 2.760 2.105 3.010 ;
        RECT 2.105 2.750 2.115 3.000 ;
        RECT 2.115 2.740 2.125 2.990 ;
        RECT 2.125 2.730 2.135 2.980 ;
        RECT 2.135 2.720 2.145 2.970 ;
        RECT 2.145 2.710 2.155 2.960 ;
        RECT 2.155 2.700 2.165 2.950 ;
        RECT 1.995 2.860 2.005 3.030 ;
        RECT 2.005 2.850 2.015 3.030 ;
        RECT 2.015 2.840 2.025 3.030 ;
        RECT 2.025 2.830 2.035 3.030 ;
        RECT 2.035 2.820 2.045 3.030 ;
        RECT 2.045 2.810 2.055 3.030 ;
        RECT 2.055 2.800 2.065 3.030 ;
        RECT 2.065 2.790 2.075 3.030 ;
        RECT 2.075 2.780 2.085 3.030 ;
        RECT 3.220 1.505 3.270 1.675 ;
        RECT 3.530 2.325 3.740 2.495 ;
        RECT 3.120 0.785 4.140 0.955 ;
        RECT 3.970 0.785 4.140 1.515 ;
        RECT 3.970 1.345 4.705 1.515 ;
        RECT 4.535 1.345 4.705 1.650 ;
        RECT 3.440 2.245 3.450 2.495 ;
        RECT 3.450 2.255 3.460 2.495 ;
        RECT 3.460 2.265 3.470 2.495 ;
        RECT 3.470 2.275 3.480 2.495 ;
        RECT 3.480 2.285 3.490 2.495 ;
        RECT 3.490 2.295 3.500 2.495 ;
        RECT 3.500 2.305 3.510 2.495 ;
        RECT 3.510 2.315 3.520 2.495 ;
        RECT 3.520 2.325 3.530 2.495 ;
        RECT 3.270 1.505 3.280 2.325 ;
        RECT 3.280 1.505 3.290 2.335 ;
        RECT 3.290 1.505 3.300 2.345 ;
        RECT 3.300 1.505 3.310 2.355 ;
        RECT 3.310 1.505 3.320 2.365 ;
        RECT 3.320 1.505 3.330 2.375 ;
        RECT 3.330 1.505 3.340 2.385 ;
        RECT 3.340 1.505 3.350 2.395 ;
        RECT 3.350 1.505 3.360 2.405 ;
        RECT 3.360 1.505 3.370 2.415 ;
        RECT 3.370 1.505 3.380 2.425 ;
        RECT 3.380 1.505 3.390 2.435 ;
        RECT 3.390 1.505 3.400 2.445 ;
        RECT 3.400 1.505 3.410 2.455 ;
        RECT 3.410 1.505 3.420 2.465 ;
        RECT 3.420 1.505 3.430 2.475 ;
        RECT 3.430 1.505 3.440 2.485 ;
        RECT 3.130 1.425 3.140 1.675 ;
        RECT 3.140 1.435 3.150 1.675 ;
        RECT 3.150 1.445 3.160 1.675 ;
        RECT 3.160 1.455 3.170 1.675 ;
        RECT 3.170 1.465 3.180 1.675 ;
        RECT 3.180 1.475 3.190 1.675 ;
        RECT 3.190 1.485 3.200 1.675 ;
        RECT 3.200 1.495 3.210 1.675 ;
        RECT 3.210 1.505 3.220 1.675 ;
        RECT 3.120 1.415 3.130 1.665 ;
        RECT 2.950 0.785 2.960 1.495 ;
        RECT 2.960 0.785 2.970 1.505 ;
        RECT 2.970 0.785 2.980 1.515 ;
        RECT 2.980 0.785 2.990 1.525 ;
        RECT 2.990 0.785 3.000 1.535 ;
        RECT 3.000 0.785 3.010 1.545 ;
        RECT 3.010 0.785 3.020 1.555 ;
        RECT 3.020 0.785 3.030 1.565 ;
        RECT 3.030 0.785 3.040 1.575 ;
        RECT 3.040 0.785 3.050 1.585 ;
        RECT 3.050 0.785 3.060 1.595 ;
        RECT 3.060 0.785 3.070 1.605 ;
        RECT 3.070 0.785 3.080 1.615 ;
        RECT 3.080 0.785 3.090 1.625 ;
        RECT 3.090 0.785 3.100 1.635 ;
        RECT 3.100 0.785 3.110 1.645 ;
        RECT 3.110 0.785 3.120 1.655 ;
        RECT 5.650 1.745 5.950 1.935 ;
        RECT 5.650 1.765 6.690 1.935 ;
        RECT 6.520 1.765 6.690 2.190 ;
        RECT 7.250 1.185 7.550 1.355 ;
        RECT 7.315 2.020 7.485 2.390 ;
        RECT 7.380 1.185 7.550 2.190 ;
        RECT 6.520 2.020 7.550 2.190 ;
        RECT 1.520 0.780 1.690 1.730 ;
        RECT 1.515 2.370 1.965 2.540 ;
        RECT 1.520 1.560 2.030 1.730 ;
        RECT 1.995 2.340 2.055 2.540 ;
        RECT 2.085 2.340 2.135 2.510 ;
        RECT 2.305 2.340 2.935 2.510 ;
        RECT 3.360 2.675 3.595 2.855 ;
        RECT 3.360 2.685 4.930 2.855 ;
        RECT 4.760 2.685 4.930 3.140 ;
        RECT 6.440 2.570 6.610 3.140 ;
        RECT 4.760 2.970 6.610 3.140 ;
        RECT 6.440 2.570 7.625 2.740 ;
        RECT 7.455 2.570 7.625 2.880 ;
        RECT 3.280 2.605 3.290 2.855 ;
        RECT 3.290 2.615 3.300 2.855 ;
        RECT 3.300 2.625 3.310 2.855 ;
        RECT 3.310 2.635 3.320 2.855 ;
        RECT 3.320 2.645 3.330 2.855 ;
        RECT 3.330 2.655 3.340 2.855 ;
        RECT 3.340 2.665 3.350 2.855 ;
        RECT 3.350 2.675 3.360 2.855 ;
        RECT 3.025 2.350 3.035 2.600 ;
        RECT 3.035 2.360 3.045 2.610 ;
        RECT 3.045 2.370 3.055 2.620 ;
        RECT 3.055 2.380 3.065 2.630 ;
        RECT 3.065 2.390 3.075 2.640 ;
        RECT 3.075 2.400 3.085 2.650 ;
        RECT 3.085 2.410 3.095 2.660 ;
        RECT 3.095 2.420 3.105 2.670 ;
        RECT 3.105 2.430 3.115 2.680 ;
        RECT 3.115 2.440 3.125 2.690 ;
        RECT 3.125 2.450 3.135 2.700 ;
        RECT 3.135 2.460 3.145 2.710 ;
        RECT 3.145 2.470 3.155 2.720 ;
        RECT 3.155 2.480 3.165 2.730 ;
        RECT 3.165 2.490 3.175 2.740 ;
        RECT 3.175 2.500 3.185 2.750 ;
        RECT 3.185 2.510 3.195 2.760 ;
        RECT 3.195 2.520 3.205 2.770 ;
        RECT 3.205 2.530 3.215 2.780 ;
        RECT 3.215 2.540 3.225 2.790 ;
        RECT 3.225 2.550 3.235 2.800 ;
        RECT 3.235 2.560 3.245 2.810 ;
        RECT 3.245 2.570 3.255 2.820 ;
        RECT 3.255 2.580 3.265 2.830 ;
        RECT 3.265 2.590 3.275 2.840 ;
        RECT 3.275 2.595 3.281 2.849 ;
        RECT 2.935 2.340 2.945 2.510 ;
        RECT 2.945 2.340 2.955 2.520 ;
        RECT 2.955 2.340 2.965 2.530 ;
        RECT 2.965 2.340 2.975 2.540 ;
        RECT 2.975 2.340 2.985 2.550 ;
        RECT 2.985 2.340 2.995 2.560 ;
        RECT 2.995 2.340 3.005 2.570 ;
        RECT 3.005 2.340 3.015 2.580 ;
        RECT 3.015 2.340 3.025 2.590 ;
        RECT 2.135 1.600 2.145 2.510 ;
        RECT 2.145 1.610 2.155 2.510 ;
        RECT 2.155 1.620 2.165 2.510 ;
        RECT 2.165 1.630 2.175 2.510 ;
        RECT 2.175 1.640 2.185 2.510 ;
        RECT 2.185 1.650 2.195 2.510 ;
        RECT 2.195 1.660 2.205 2.510 ;
        RECT 2.205 1.670 2.215 2.510 ;
        RECT 2.215 1.680 2.225 2.510 ;
        RECT 2.225 1.690 2.235 2.510 ;
        RECT 2.235 1.700 2.245 2.510 ;
        RECT 2.245 1.710 2.255 2.510 ;
        RECT 2.255 1.720 2.265 2.510 ;
        RECT 2.265 1.730 2.275 2.510 ;
        RECT 2.275 1.740 2.285 2.510 ;
        RECT 2.285 1.750 2.295 2.510 ;
        RECT 2.295 1.760 2.305 2.510 ;
        RECT 2.105 1.570 2.115 1.804 ;
        RECT 2.115 1.580 2.125 1.814 ;
        RECT 2.125 1.590 2.135 1.824 ;
        RECT 2.030 1.560 2.040 1.730 ;
        RECT 2.040 1.560 2.050 1.740 ;
        RECT 2.050 1.560 2.060 1.750 ;
        RECT 2.060 1.560 2.070 1.760 ;
        RECT 2.070 1.560 2.080 1.770 ;
        RECT 2.080 1.560 2.090 1.780 ;
        RECT 2.090 1.560 2.100 1.790 ;
        RECT 2.100 1.560 2.106 1.800 ;
        RECT 2.055 2.340 2.065 2.530 ;
        RECT 2.065 2.340 2.075 2.520 ;
        RECT 2.075 2.340 2.085 2.510 ;
        RECT 1.965 2.370 1.975 2.540 ;
        RECT 1.975 2.360 1.985 2.540 ;
        RECT 1.985 2.350 1.995 2.540 ;
        RECT 4.885 0.970 5.055 2.330 ;
        RECT 4.885 2.160 6.095 2.330 ;
        RECT 5.440 0.565 6.085 1.140 ;
        RECT 5.455 2.160 6.095 2.670 ;
        RECT 6.900 0.815 7.070 1.140 ;
        RECT 4.885 0.970 7.070 1.140 ;
        RECT 6.900 0.815 7.695 0.985 ;
  END 
END MUXI4HD2XHT

MACRO MUXI4HD1XHT
  CLASS  CORE ;
  FOREIGN MUXI4HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.200 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.240 2.620 6.750 2.830 ;
        RECT 6.450 2.500 6.520 2.855 ;
        RECT 6.240 2.500 6.520 2.830 ;
        RECT 6.450 2.620 6.750 2.855 ;
    END
  END S1
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.165 1.890 4.420 2.440 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.485 1.730 2.830 2.140 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.060 0.920 2.525 1.450 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 1.200 1.230 1.665 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.665 ;
        RECT 2.375 -0.300 2.675 0.740 ;
        RECT 4.380 -0.300 4.680 0.655 ;
        RECT 5.930 -0.300 6.230 0.665 ;
        RECT 7.275 -0.300 7.445 1.120 ;
        RECT 0.000 -0.300 8.200 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.340 2.120 8.030 2.415 ;
        RECT 7.795 0.720 8.030 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.675 3.040 0.975 3.990 ;
        RECT 2.385 3.040 2.685 3.990 ;
        RECT 4.280 3.035 4.580 3.990 ;
        RECT 6.080 3.025 6.380 3.990 ;
        RECT 7.150 2.635 7.450 3.990 ;
        RECT 0.000 3.390 8.200 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.910 0.680 2.420 ;
        RECT 0.510 2.000 0.720 2.420 ;
        RECT 0.510 2.000 1.955 2.170 ;
        RECT 3.300 1.155 3.790 1.325 ;
        RECT 3.620 1.155 3.790 2.125 ;
        RECT 3.620 1.955 3.920 2.125 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.105 1.075 0.275 2.860 ;
        RECT 0.105 1.075 0.405 1.245 ;
        RECT 0.105 2.600 0.405 2.860 ;
        RECT 1.165 2.690 1.335 3.030 ;
        RECT 0.105 2.690 1.335 2.860 ;
        RECT 1.165 2.860 2.045 3.030 ;
        RECT 2.305 2.690 2.765 2.860 ;
        RECT 3.030 2.865 3.035 3.210 ;
        RECT 3.030 3.040 3.325 3.210 ;
        RECT 2.865 2.710 2.875 3.210 ;
        RECT 2.875 2.720 2.885 3.210 ;
        RECT 2.885 2.730 2.895 3.210 ;
        RECT 2.895 2.740 2.905 3.210 ;
        RECT 2.905 2.750 2.915 3.210 ;
        RECT 2.915 2.760 2.925 3.210 ;
        RECT 2.925 2.770 2.935 3.210 ;
        RECT 2.935 2.780 2.945 3.210 ;
        RECT 2.945 2.790 2.955 3.210 ;
        RECT 2.955 2.800 2.965 3.210 ;
        RECT 2.965 2.810 2.975 3.210 ;
        RECT 2.975 2.820 2.985 3.210 ;
        RECT 2.985 2.830 2.995 3.210 ;
        RECT 2.995 2.840 3.005 3.210 ;
        RECT 3.005 2.850 3.015 3.210 ;
        RECT 3.015 2.860 3.025 3.210 ;
        RECT 3.025 2.865 3.031 3.209 ;
        RECT 2.855 2.700 2.865 2.950 ;
        RECT 2.765 2.690 2.775 2.860 ;
        RECT 2.775 2.690 2.785 2.870 ;
        RECT 2.785 2.690 2.795 2.880 ;
        RECT 2.795 2.690 2.805 2.890 ;
        RECT 2.805 2.690 2.815 2.900 ;
        RECT 2.815 2.690 2.825 2.910 ;
        RECT 2.825 2.690 2.835 2.920 ;
        RECT 2.835 2.690 2.845 2.930 ;
        RECT 2.845 2.690 2.855 2.940 ;
        RECT 2.215 2.690 2.225 2.940 ;
        RECT 2.225 2.690 2.235 2.930 ;
        RECT 2.235 2.690 2.245 2.920 ;
        RECT 2.245 2.690 2.255 2.910 ;
        RECT 2.255 2.690 2.265 2.900 ;
        RECT 2.265 2.690 2.275 2.890 ;
        RECT 2.275 2.690 2.285 2.880 ;
        RECT 2.285 2.690 2.295 2.870 ;
        RECT 2.295 2.690 2.305 2.860 ;
        RECT 2.135 2.770 2.145 3.020 ;
        RECT 2.145 2.760 2.155 3.010 ;
        RECT 2.155 2.750 2.165 3.000 ;
        RECT 2.165 2.740 2.175 2.990 ;
        RECT 2.175 2.730 2.185 2.980 ;
        RECT 2.185 2.720 2.195 2.970 ;
        RECT 2.195 2.710 2.205 2.960 ;
        RECT 2.205 2.700 2.215 2.950 ;
        RECT 2.045 2.860 2.055 3.030 ;
        RECT 2.055 2.850 2.065 3.030 ;
        RECT 2.065 2.840 2.075 3.030 ;
        RECT 2.075 2.830 2.085 3.030 ;
        RECT 2.085 2.820 2.095 3.030 ;
        RECT 2.095 2.810 2.105 3.030 ;
        RECT 2.105 2.800 2.115 3.030 ;
        RECT 2.115 2.790 2.125 3.030 ;
        RECT 2.125 2.780 2.135 3.030 ;
        RECT 3.220 1.505 3.270 1.675 ;
        RECT 3.530 2.325 3.740 2.495 ;
        RECT 3.120 0.785 4.140 0.955 ;
        RECT 3.970 0.785 4.140 1.325 ;
        RECT 3.970 1.155 4.785 1.325 ;
        RECT 4.615 1.155 4.785 1.780 ;
        RECT 3.440 2.245 3.450 2.495 ;
        RECT 3.450 2.255 3.460 2.495 ;
        RECT 3.460 2.265 3.470 2.495 ;
        RECT 3.470 2.275 3.480 2.495 ;
        RECT 3.480 2.285 3.490 2.495 ;
        RECT 3.490 2.295 3.500 2.495 ;
        RECT 3.500 2.305 3.510 2.495 ;
        RECT 3.510 2.315 3.520 2.495 ;
        RECT 3.520 2.325 3.530 2.495 ;
        RECT 3.270 1.505 3.280 2.325 ;
        RECT 3.280 1.505 3.290 2.335 ;
        RECT 3.290 1.505 3.300 2.345 ;
        RECT 3.300 1.505 3.310 2.355 ;
        RECT 3.310 1.505 3.320 2.365 ;
        RECT 3.320 1.505 3.330 2.375 ;
        RECT 3.330 1.505 3.340 2.385 ;
        RECT 3.340 1.505 3.350 2.395 ;
        RECT 3.350 1.505 3.360 2.405 ;
        RECT 3.360 1.505 3.370 2.415 ;
        RECT 3.370 1.505 3.380 2.425 ;
        RECT 3.380 1.505 3.390 2.435 ;
        RECT 3.390 1.505 3.400 2.445 ;
        RECT 3.400 1.505 3.410 2.455 ;
        RECT 3.410 1.505 3.420 2.465 ;
        RECT 3.420 1.505 3.430 2.475 ;
        RECT 3.430 1.505 3.440 2.485 ;
        RECT 3.130 1.425 3.140 1.675 ;
        RECT 3.140 1.435 3.150 1.675 ;
        RECT 3.150 1.445 3.160 1.675 ;
        RECT 3.160 1.455 3.170 1.675 ;
        RECT 3.170 1.465 3.180 1.675 ;
        RECT 3.180 1.475 3.190 1.675 ;
        RECT 3.190 1.485 3.200 1.675 ;
        RECT 3.200 1.495 3.210 1.675 ;
        RECT 3.210 1.505 3.220 1.675 ;
        RECT 3.120 1.415 3.130 1.665 ;
        RECT 2.950 0.785 2.960 1.495 ;
        RECT 2.960 0.785 2.970 1.505 ;
        RECT 2.970 0.785 2.980 1.515 ;
        RECT 2.980 0.785 2.990 1.525 ;
        RECT 2.990 0.785 3.000 1.535 ;
        RECT 3.000 0.785 3.010 1.545 ;
        RECT 3.010 0.785 3.020 1.555 ;
        RECT 3.020 0.785 3.030 1.565 ;
        RECT 3.030 0.785 3.040 1.575 ;
        RECT 3.040 0.785 3.050 1.585 ;
        RECT 3.050 0.785 3.060 1.595 ;
        RECT 3.060 0.785 3.070 1.605 ;
        RECT 3.070 0.785 3.080 1.615 ;
        RECT 3.080 0.785 3.090 1.625 ;
        RECT 3.090 0.785 3.100 1.635 ;
        RECT 3.100 0.785 3.110 1.645 ;
        RECT 3.110 0.785 3.120 1.655 ;
        RECT 1.520 0.720 1.690 1.820 ;
        RECT 1.515 2.370 2.015 2.540 ;
        RECT 2.045 2.340 2.105 2.540 ;
        RECT 1.520 1.650 2.305 1.820 ;
        RECT 2.135 1.650 2.305 2.510 ;
        RECT 2.135 2.340 2.935 2.510 ;
        RECT 3.360 2.675 5.710 2.855 ;
        RECT 6.105 1.610 6.165 2.190 ;
        RECT 5.995 1.610 6.005 2.290 ;
        RECT 6.005 1.610 6.015 2.280 ;
        RECT 6.015 1.610 6.025 2.270 ;
        RECT 6.025 1.610 6.035 2.260 ;
        RECT 6.035 1.610 6.045 2.250 ;
        RECT 6.045 1.610 6.055 2.240 ;
        RECT 6.055 1.610 6.065 2.230 ;
        RECT 6.065 1.610 6.075 2.220 ;
        RECT 6.075 1.610 6.085 2.210 ;
        RECT 6.085 1.610 6.095 2.200 ;
        RECT 6.095 1.610 6.105 2.190 ;
        RECT 5.825 2.210 5.835 2.800 ;
        RECT 5.835 2.200 5.845 2.790 ;
        RECT 5.845 2.190 5.855 2.780 ;
        RECT 5.855 2.180 5.865 2.770 ;
        RECT 5.865 2.170 5.875 2.760 ;
        RECT 5.875 2.160 5.885 2.750 ;
        RECT 5.885 2.150 5.895 2.740 ;
        RECT 5.895 2.140 5.905 2.730 ;
        RECT 5.905 2.130 5.915 2.720 ;
        RECT 5.915 2.120 5.925 2.710 ;
        RECT 5.925 2.110 5.935 2.700 ;
        RECT 5.935 2.100 5.945 2.690 ;
        RECT 5.945 2.090 5.955 2.680 ;
        RECT 5.955 2.080 5.965 2.670 ;
        RECT 5.965 2.070 5.975 2.660 ;
        RECT 5.975 2.060 5.985 2.650 ;
        RECT 5.985 2.050 5.995 2.640 ;
        RECT 5.780 2.605 5.790 2.845 ;
        RECT 5.790 2.595 5.800 2.835 ;
        RECT 5.800 2.585 5.810 2.825 ;
        RECT 5.810 2.575 5.820 2.815 ;
        RECT 5.820 2.565 5.826 2.809 ;
        RECT 5.710 2.675 5.720 2.855 ;
        RECT 5.720 2.665 5.730 2.855 ;
        RECT 5.730 2.655 5.740 2.855 ;
        RECT 5.740 2.645 5.750 2.855 ;
        RECT 5.750 2.635 5.760 2.855 ;
        RECT 5.760 2.625 5.770 2.855 ;
        RECT 5.770 2.615 5.780 2.855 ;
        RECT 3.280 2.605 3.290 2.855 ;
        RECT 3.290 2.615 3.300 2.855 ;
        RECT 3.300 2.625 3.310 2.855 ;
        RECT 3.310 2.635 3.320 2.855 ;
        RECT 3.320 2.645 3.330 2.855 ;
        RECT 3.330 2.655 3.340 2.855 ;
        RECT 3.340 2.665 3.350 2.855 ;
        RECT 3.350 2.675 3.360 2.855 ;
        RECT 3.025 2.350 3.035 2.600 ;
        RECT 3.035 2.360 3.045 2.610 ;
        RECT 3.045 2.370 3.055 2.620 ;
        RECT 3.055 2.380 3.065 2.630 ;
        RECT 3.065 2.390 3.075 2.640 ;
        RECT 3.075 2.400 3.085 2.650 ;
        RECT 3.085 2.410 3.095 2.660 ;
        RECT 3.095 2.420 3.105 2.670 ;
        RECT 3.105 2.430 3.115 2.680 ;
        RECT 3.115 2.440 3.125 2.690 ;
        RECT 3.125 2.450 3.135 2.700 ;
        RECT 3.135 2.460 3.145 2.710 ;
        RECT 3.145 2.470 3.155 2.720 ;
        RECT 3.155 2.480 3.165 2.730 ;
        RECT 3.165 2.490 3.175 2.740 ;
        RECT 3.175 2.500 3.185 2.750 ;
        RECT 3.185 2.510 3.195 2.760 ;
        RECT 3.195 2.520 3.205 2.770 ;
        RECT 3.205 2.530 3.215 2.780 ;
        RECT 3.215 2.540 3.225 2.790 ;
        RECT 3.225 2.550 3.235 2.800 ;
        RECT 3.235 2.560 3.245 2.810 ;
        RECT 3.245 2.570 3.255 2.820 ;
        RECT 3.255 2.580 3.265 2.830 ;
        RECT 3.265 2.590 3.275 2.840 ;
        RECT 3.275 2.595 3.281 2.849 ;
        RECT 2.935 2.340 2.945 2.510 ;
        RECT 2.945 2.340 2.955 2.520 ;
        RECT 2.955 2.340 2.965 2.530 ;
        RECT 2.965 2.340 2.975 2.540 ;
        RECT 2.975 2.340 2.985 2.550 ;
        RECT 2.985 2.340 2.995 2.560 ;
        RECT 2.995 2.340 3.005 2.570 ;
        RECT 3.005 2.340 3.015 2.580 ;
        RECT 3.015 2.340 3.025 2.590 ;
        RECT 2.105 2.340 2.115 2.530 ;
        RECT 2.115 2.340 2.125 2.520 ;
        RECT 2.125 2.340 2.135 2.510 ;
        RECT 2.015 2.370 2.025 2.540 ;
        RECT 2.025 2.360 2.035 2.540 ;
        RECT 2.035 2.350 2.045 2.540 ;
        RECT 5.620 1.795 5.700 1.995 ;
        RECT 5.610 1.805 5.806 1.869 ;
        RECT 5.630 1.785 5.700 1.995 ;
        RECT 5.600 1.815 5.806 1.869 ;
        RECT 5.400 1.825 5.700 1.995 ;
        RECT 5.400 1.825 5.710 1.965 ;
        RECT 5.400 1.825 5.720 1.955 ;
        RECT 5.400 1.825 5.730 1.945 ;
        RECT 5.400 1.825 5.740 1.935 ;
        RECT 5.400 1.825 5.750 1.925 ;
        RECT 5.400 1.825 5.760 1.915 ;
        RECT 5.400 1.825 5.770 1.905 ;
        RECT 5.400 1.825 5.780 1.895 ;
        RECT 5.400 1.825 5.790 1.885 ;
        RECT 5.400 1.825 5.800 1.875 ;
        RECT 5.635 1.255 5.806 1.869 ;
        RECT 5.635 1.255 6.865 1.425 ;
        RECT 6.695 1.040 6.865 2.430 ;
        RECT 4.965 1.170 5.135 2.495 ;
        RECT 5.285 0.905 5.455 1.340 ;
        RECT 4.965 1.170 5.455 1.340 ;
        RECT 4.965 2.325 5.520 2.495 ;
        RECT 5.285 0.905 6.310 1.075 ;
        RECT 6.615 0.690 7.095 0.860 ;
        RECT 6.525 0.690 6.535 0.940 ;
        RECT 6.535 0.690 6.545 0.930 ;
        RECT 6.545 0.690 6.555 0.920 ;
        RECT 6.555 0.690 6.565 0.910 ;
        RECT 6.565 0.690 6.575 0.900 ;
        RECT 6.575 0.690 6.585 0.890 ;
        RECT 6.585 0.690 6.595 0.880 ;
        RECT 6.595 0.690 6.605 0.870 ;
        RECT 6.605 0.690 6.615 0.860 ;
        RECT 6.400 0.815 6.410 1.065 ;
        RECT 6.410 0.805 6.420 1.055 ;
        RECT 6.420 0.795 6.430 1.045 ;
        RECT 6.430 0.785 6.440 1.035 ;
        RECT 6.440 0.775 6.450 1.025 ;
        RECT 6.450 0.765 6.460 1.015 ;
        RECT 6.460 0.755 6.470 1.005 ;
        RECT 6.470 0.745 6.480 0.995 ;
        RECT 6.480 0.735 6.490 0.985 ;
        RECT 6.490 0.725 6.500 0.975 ;
        RECT 6.500 0.715 6.510 0.965 ;
        RECT 6.510 0.705 6.520 0.955 ;
        RECT 6.520 0.695 6.526 0.949 ;
        RECT 6.310 0.905 6.320 1.075 ;
        RECT 6.320 0.895 6.330 1.075 ;
        RECT 6.330 0.885 6.340 1.075 ;
        RECT 6.340 0.875 6.350 1.075 ;
        RECT 6.350 0.865 6.360 1.075 ;
        RECT 6.360 0.855 6.370 1.075 ;
        RECT 6.370 0.845 6.380 1.075 ;
        RECT 6.380 0.835 6.390 1.075 ;
        RECT 6.390 0.825 6.400 1.075 ;
  END 
END MUXI4HD1XHT

MACRO MUXI2HDMXHT
  CLASS  CORE ;
  FOREIGN MUXI2HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.510 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.710 1.570 1.200 1.950 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.240 1.860 2.410 2.360 ;
        RECT 2.240 2.150 2.830 2.360 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 2.405 -0.300 2.705 1.295 ;
        RECT 3.435 -0.300 3.735 1.145 ;
        RECT 0.000 -0.300 4.510 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.955 1.125 4.270 1.295 ;
        RECT 4.100 1.125 4.270 2.215 ;
        RECT 3.955 2.045 4.270 2.215 ;
        RECT 4.100 1.670 4.410 2.010 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.540 0.925 3.990 ;
        RECT 2.405 2.540 2.705 3.990 ;
        RECT 3.435 2.375 3.735 3.990 ;
        RECT 0.000 3.390 4.510 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.200 2.860 1.775 3.180 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.655 ;
        RECT 1.400 1.695 1.570 2.300 ;
        RECT 0.170 2.130 1.570 2.300 ;
        RECT 1.515 1.125 1.920 1.295 ;
        RECT 1.750 1.125 1.920 2.650 ;
        RECT 1.515 2.480 1.920 2.650 ;
        RECT 1.750 1.475 2.890 1.645 ;
        RECT 2.720 1.475 2.890 1.870 ;
        RECT 2.925 1.125 3.240 1.295 ;
        RECT 3.070 1.125 3.240 2.710 ;
        RECT 2.925 2.540 3.240 2.710 ;
        RECT 3.070 1.520 3.850 1.820 ;
  END 
END MUXI2HDMXHT

MACRO MUXI2HDLXHT
  CLASS  CORE ;
  FOREIGN MUXI2HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.510 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.720 1.570 1.200 1.950 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.240 1.860 2.410 2.360 ;
        RECT 2.240 2.150 2.830 2.360 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 2.405 -0.300 2.705 1.295 ;
        RECT 3.435 -0.300 3.735 1.295 ;
        RECT 0.000 -0.300 4.510 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.955 1.125 4.270 1.295 ;
        RECT 4.100 1.125 4.270 2.215 ;
        RECT 3.955 2.045 4.270 2.215 ;
        RECT 4.100 1.670 4.410 2.010 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.540 0.925 3.990 ;
        RECT 2.405 2.540 2.705 3.990 ;
        RECT 3.435 2.165 3.735 3.990 ;
        RECT 0.000 3.390 4.510 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.200 2.860 1.775 3.180 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.655 ;
        RECT 1.400 1.695 1.570 2.300 ;
        RECT 0.170 2.130 1.570 2.300 ;
        RECT 1.515 1.125 1.920 1.295 ;
        RECT 1.750 1.125 1.920 2.650 ;
        RECT 1.515 2.480 1.920 2.650 ;
        RECT 1.750 1.475 2.890 1.645 ;
        RECT 2.720 1.475 2.890 1.870 ;
        RECT 2.925 1.125 3.240 1.295 ;
        RECT 3.070 1.125 3.240 2.710 ;
        RECT 2.925 2.540 3.240 2.710 ;
        RECT 3.070 1.515 3.850 1.815 ;
  END 
END MUXI2HDLXHT

MACRO MUXI2HD3XHT
  CLASS  CORE ;
  FOREIGN MUXI2HD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.740 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.330 1.155 1.540 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.675 2.360 2.430 ;
        RECT 2.150 1.675 2.555 1.845 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.065 ;
        RECT 2.485 -0.300 2.785 1.055 ;
        RECT 3.580 -0.300 3.815 1.120 ;
        RECT 4.555 -0.300 4.855 1.055 ;
        RECT 0.000 -0.300 5.740 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.035 0.720 4.335 1.430 ;
        RECT 4.035 1.980 4.335 2.960 ;
        RECT 4.035 1.235 5.375 1.430 ;
        RECT 4.675 1.235 5.375 2.455 ;
        RECT 4.035 1.980 5.375 2.455 ;
        RECT 5.075 0.720 5.375 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.900 0.955 3.990 ;
        RECT 2.550 2.230 2.720 3.990 ;
        RECT 3.580 2.230 3.815 3.990 ;
        RECT 4.555 2.635 4.855 3.990 ;
        RECT 0.000 3.390 5.740 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 2.550 1.665 2.720 ;
        RECT 1.225 2.550 1.665 2.770 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.090 0.895 0.260 1.890 ;
        RECT 0.170 1.720 0.340 2.290 ;
        RECT 0.090 0.895 0.405 1.065 ;
        RECT 1.430 1.330 1.600 1.890 ;
        RECT 0.090 1.720 1.600 1.890 ;
        RECT 1.545 0.895 1.950 1.065 ;
        RECT 1.780 0.895 1.950 2.315 ;
        RECT 1.545 2.145 1.950 2.315 ;
        RECT 1.780 1.325 2.990 1.495 ;
        RECT 2.755 1.325 2.990 1.730 ;
        RECT 3.005 0.555 3.390 1.065 ;
        RECT 3.190 0.555 3.390 2.960 ;
        RECT 3.005 1.980 3.390 2.960 ;
        RECT 3.190 1.610 4.495 1.780 ;
  END 
END MUXI2HD3XHT

MACRO MUXI2HD2XHT
  CLASS  CORE ;
  FOREIGN MUXI2HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.680 1.570 1.200 1.950 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.240 1.860 2.410 2.360 ;
        RECT 2.240 2.150 2.830 2.360 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 2.405 -0.300 2.705 1.295 ;
        RECT 3.435 -0.300 3.735 1.055 ;
        RECT 4.475 -0.300 4.775 1.055 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.020 0.720 4.270 2.960 ;
        RECT 4.020 1.670 4.410 2.010 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.540 0.925 3.990 ;
        RECT 2.405 2.540 2.705 3.990 ;
        RECT 3.435 2.295 3.735 3.990 ;
        RECT 4.475 2.295 4.775 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.200 2.860 1.775 3.180 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.655 ;
        RECT 1.400 1.695 1.570 2.300 ;
        RECT 0.170 2.130 1.570 2.300 ;
        RECT 1.515 1.125 1.920 1.295 ;
        RECT 1.750 1.125 1.920 2.650 ;
        RECT 1.515 2.480 1.920 2.650 ;
        RECT 1.750 1.475 2.890 1.645 ;
        RECT 2.720 1.475 2.890 1.870 ;
        RECT 2.925 1.125 3.240 1.295 ;
        RECT 3.070 1.125 3.240 2.710 ;
        RECT 2.925 2.540 3.240 2.710 ;
        RECT 3.070 1.610 3.775 1.910 ;
  END 
END MUXI2HD2XHT

MACRO MUXI2HD1XHT
  CLASS  CORE ;
  FOREIGN MUXI2HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.510 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.680 1.570 1.200 1.950 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.175 1.860 2.410 2.360 ;
        RECT 2.175 2.150 2.830 2.360 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 2.405 -0.300 2.705 1.295 ;
        RECT 3.435 -0.300 3.735 1.055 ;
        RECT 0.000 -0.300 4.510 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.020 0.720 4.190 2.960 ;
        RECT 4.020 1.670 4.410 2.010 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.540 0.925 3.990 ;
        RECT 2.405 2.540 2.705 3.990 ;
        RECT 3.435 2.295 3.735 3.990 ;
        RECT 0.000 3.390 4.510 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.200 2.860 1.775 3.180 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.655 ;
        RECT 1.400 1.695 1.570 2.300 ;
        RECT 0.170 2.130 1.570 2.300 ;
        RECT 1.515 1.125 1.920 1.295 ;
        RECT 1.750 1.125 1.920 2.650 ;
        RECT 1.515 2.480 1.920 2.650 ;
        RECT 1.750 1.475 2.890 1.645 ;
        RECT 2.720 1.475 2.890 1.870 ;
        RECT 2.925 1.125 3.240 1.295 ;
        RECT 3.070 1.125 3.240 2.710 ;
        RECT 2.925 2.540 3.240 2.710 ;
        RECT 3.070 1.610 3.775 1.910 ;
  END 
END MUXI2HD1XHT

MACRO MUX4HDMXHT
  CLASS  CORE ;
  FOREIGN MUX4HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.610 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.240 2.500 6.750 2.830 ;
    END
  END S1
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.175 1.890 4.420 2.440 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.485 1.730 2.830 2.140 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.060 0.920 2.525 1.385 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 1.060 1.140 1.665 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.665 ;
        RECT 2.375 -0.300 2.675 0.740 ;
        RECT 4.380 -0.300 4.680 0.680 ;
        RECT 5.930 -0.300 6.230 0.725 ;
        RECT 7.595 -0.300 7.895 0.715 ;
        RECT 0.000 -0.300 8.610 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.760 2.120 8.450 2.415 ;
        RECT 8.215 1.060 8.450 2.450 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.675 3.040 0.975 3.990 ;
        RECT 2.385 3.040 2.685 3.990 ;
        RECT 4.380 3.025 4.680 3.990 ;
        RECT 6.080 3.025 6.380 3.990 ;
        RECT 7.595 2.730 7.895 3.990 ;
        RECT 0.000 3.390 8.610 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.500 1.910 0.680 2.420 ;
        RECT 0.500 2.000 0.780 2.420 ;
        RECT 0.500 2.000 1.955 2.170 ;
        RECT 3.300 1.155 3.790 1.325 ;
        RECT 3.620 1.155 3.790 2.125 ;
        RECT 3.620 1.955 3.920 2.125 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.105 1.075 0.275 2.860 ;
        RECT 0.105 1.075 0.405 1.245 ;
        RECT 0.105 2.600 0.405 2.860 ;
        RECT 1.165 2.690 1.335 3.030 ;
        RECT 0.105 2.690 1.335 2.860 ;
        RECT 1.165 2.860 2.045 3.030 ;
        RECT 2.305 2.690 2.765 2.860 ;
        RECT 3.030 2.865 3.035 3.210 ;
        RECT 3.030 3.040 3.325 3.210 ;
        RECT 2.865 2.710 2.875 3.210 ;
        RECT 2.875 2.720 2.885 3.210 ;
        RECT 2.885 2.730 2.895 3.210 ;
        RECT 2.895 2.740 2.905 3.210 ;
        RECT 2.905 2.750 2.915 3.210 ;
        RECT 2.915 2.760 2.925 3.210 ;
        RECT 2.925 2.770 2.935 3.210 ;
        RECT 2.935 2.780 2.945 3.210 ;
        RECT 2.945 2.790 2.955 3.210 ;
        RECT 2.955 2.800 2.965 3.210 ;
        RECT 2.965 2.810 2.975 3.210 ;
        RECT 2.975 2.820 2.985 3.210 ;
        RECT 2.985 2.830 2.995 3.210 ;
        RECT 2.995 2.840 3.005 3.210 ;
        RECT 3.005 2.850 3.015 3.210 ;
        RECT 3.015 2.860 3.025 3.210 ;
        RECT 3.025 2.865 3.031 3.209 ;
        RECT 2.855 2.700 2.865 2.950 ;
        RECT 2.765 2.690 2.775 2.860 ;
        RECT 2.775 2.690 2.785 2.870 ;
        RECT 2.785 2.690 2.795 2.880 ;
        RECT 2.795 2.690 2.805 2.890 ;
        RECT 2.805 2.690 2.815 2.900 ;
        RECT 2.815 2.690 2.825 2.910 ;
        RECT 2.825 2.690 2.835 2.920 ;
        RECT 2.835 2.690 2.845 2.930 ;
        RECT 2.845 2.690 2.855 2.940 ;
        RECT 2.215 2.690 2.225 2.940 ;
        RECT 2.225 2.690 2.235 2.930 ;
        RECT 2.235 2.690 2.245 2.920 ;
        RECT 2.245 2.690 2.255 2.910 ;
        RECT 2.255 2.690 2.265 2.900 ;
        RECT 2.265 2.690 2.275 2.890 ;
        RECT 2.275 2.690 2.285 2.880 ;
        RECT 2.285 2.690 2.295 2.870 ;
        RECT 2.295 2.690 2.305 2.860 ;
        RECT 2.135 2.770 2.145 3.020 ;
        RECT 2.145 2.760 2.155 3.010 ;
        RECT 2.155 2.750 2.165 3.000 ;
        RECT 2.165 2.740 2.175 2.990 ;
        RECT 2.175 2.730 2.185 2.980 ;
        RECT 2.185 2.720 2.195 2.970 ;
        RECT 2.195 2.710 2.205 2.960 ;
        RECT 2.205 2.700 2.215 2.950 ;
        RECT 2.045 2.860 2.055 3.030 ;
        RECT 2.055 2.850 2.065 3.030 ;
        RECT 2.065 2.840 2.075 3.030 ;
        RECT 2.075 2.830 2.085 3.030 ;
        RECT 2.085 2.820 2.095 3.030 ;
        RECT 2.095 2.810 2.105 3.030 ;
        RECT 2.105 2.800 2.115 3.030 ;
        RECT 2.115 2.790 2.125 3.030 ;
        RECT 2.125 2.780 2.135 3.030 ;
        RECT 3.220 1.505 3.270 1.675 ;
        RECT 3.530 2.325 3.740 2.495 ;
        RECT 3.120 0.785 4.140 0.955 ;
        RECT 3.970 0.785 4.140 1.325 ;
        RECT 3.970 1.155 4.745 1.325 ;
        RECT 4.575 1.155 4.745 1.710 ;
        RECT 3.440 2.245 3.450 2.495 ;
        RECT 3.450 2.255 3.460 2.495 ;
        RECT 3.460 2.265 3.470 2.495 ;
        RECT 3.470 2.275 3.480 2.495 ;
        RECT 3.480 2.285 3.490 2.495 ;
        RECT 3.490 2.295 3.500 2.495 ;
        RECT 3.500 2.305 3.510 2.495 ;
        RECT 3.510 2.315 3.520 2.495 ;
        RECT 3.520 2.325 3.530 2.495 ;
        RECT 3.270 1.505 3.280 2.325 ;
        RECT 3.280 1.505 3.290 2.335 ;
        RECT 3.290 1.505 3.300 2.345 ;
        RECT 3.300 1.505 3.310 2.355 ;
        RECT 3.310 1.505 3.320 2.365 ;
        RECT 3.320 1.505 3.330 2.375 ;
        RECT 3.330 1.505 3.340 2.385 ;
        RECT 3.340 1.505 3.350 2.395 ;
        RECT 3.350 1.505 3.360 2.405 ;
        RECT 3.360 1.505 3.370 2.415 ;
        RECT 3.370 1.505 3.380 2.425 ;
        RECT 3.380 1.505 3.390 2.435 ;
        RECT 3.390 1.505 3.400 2.445 ;
        RECT 3.400 1.505 3.410 2.455 ;
        RECT 3.410 1.505 3.420 2.465 ;
        RECT 3.420 1.505 3.430 2.475 ;
        RECT 3.430 1.505 3.440 2.485 ;
        RECT 3.130 1.425 3.140 1.675 ;
        RECT 3.140 1.435 3.150 1.675 ;
        RECT 3.150 1.445 3.160 1.675 ;
        RECT 3.160 1.455 3.170 1.675 ;
        RECT 3.170 1.465 3.180 1.675 ;
        RECT 3.180 1.475 3.190 1.675 ;
        RECT 3.190 1.485 3.200 1.675 ;
        RECT 3.200 1.495 3.210 1.675 ;
        RECT 3.210 1.505 3.220 1.675 ;
        RECT 3.120 1.415 3.130 1.665 ;
        RECT 2.950 0.785 2.960 1.495 ;
        RECT 2.960 0.785 2.970 1.505 ;
        RECT 2.970 0.785 2.980 1.515 ;
        RECT 2.980 0.785 2.990 1.525 ;
        RECT 2.990 0.785 3.000 1.535 ;
        RECT 3.000 0.785 3.010 1.545 ;
        RECT 3.010 0.785 3.020 1.555 ;
        RECT 3.020 0.785 3.030 1.565 ;
        RECT 3.030 0.785 3.040 1.575 ;
        RECT 3.040 0.785 3.050 1.585 ;
        RECT 3.050 0.785 3.060 1.595 ;
        RECT 3.060 0.785 3.070 1.605 ;
        RECT 3.070 0.785 3.080 1.615 ;
        RECT 3.080 0.785 3.090 1.625 ;
        RECT 3.090 0.785 3.100 1.635 ;
        RECT 3.100 0.785 3.110 1.645 ;
        RECT 3.110 0.785 3.120 1.655 ;
        RECT 1.520 0.720 1.690 1.820 ;
        RECT 1.515 2.370 2.015 2.540 ;
        RECT 2.045 2.340 2.105 2.540 ;
        RECT 1.520 1.650 2.305 1.820 ;
        RECT 2.135 1.650 2.305 2.510 ;
        RECT 2.135 2.340 2.935 2.510 ;
        RECT 3.360 2.675 3.595 2.855 ;
        RECT 3.360 2.675 5.800 2.845 ;
        RECT 6.105 1.610 6.165 2.190 ;
        RECT 5.995 1.610 6.005 2.290 ;
        RECT 6.005 1.610 6.015 2.280 ;
        RECT 6.015 1.610 6.025 2.270 ;
        RECT 6.025 1.610 6.035 2.260 ;
        RECT 6.035 1.610 6.045 2.250 ;
        RECT 6.045 1.610 6.055 2.240 ;
        RECT 6.055 1.610 6.065 2.230 ;
        RECT 6.065 1.610 6.075 2.220 ;
        RECT 6.075 1.610 6.085 2.210 ;
        RECT 6.085 1.610 6.095 2.200 ;
        RECT 6.095 1.610 6.105 2.190 ;
        RECT 5.970 2.065 5.980 2.835 ;
        RECT 5.980 2.055 5.990 2.825 ;
        RECT 5.990 2.045 5.996 2.819 ;
        RECT 5.825 2.210 5.835 2.844 ;
        RECT 5.835 2.200 5.845 2.844 ;
        RECT 5.845 2.190 5.855 2.844 ;
        RECT 5.855 2.180 5.865 2.844 ;
        RECT 5.865 2.170 5.875 2.844 ;
        RECT 5.875 2.160 5.885 2.844 ;
        RECT 5.885 2.150 5.895 2.844 ;
        RECT 5.895 2.140 5.905 2.844 ;
        RECT 5.905 2.130 5.915 2.844 ;
        RECT 5.915 2.120 5.925 2.844 ;
        RECT 5.925 2.110 5.935 2.844 ;
        RECT 5.935 2.100 5.945 2.844 ;
        RECT 5.945 2.090 5.955 2.844 ;
        RECT 5.955 2.080 5.965 2.844 ;
        RECT 5.965 2.070 5.971 2.844 ;
        RECT 5.800 2.675 5.810 2.845 ;
        RECT 5.810 2.665 5.820 2.845 ;
        RECT 5.820 2.655 5.826 2.845 ;
        RECT 3.280 2.605 3.290 2.855 ;
        RECT 3.290 2.615 3.300 2.855 ;
        RECT 3.300 2.625 3.310 2.855 ;
        RECT 3.310 2.635 3.320 2.855 ;
        RECT 3.320 2.645 3.330 2.855 ;
        RECT 3.330 2.655 3.340 2.855 ;
        RECT 3.340 2.665 3.350 2.855 ;
        RECT 3.350 2.675 3.360 2.855 ;
        RECT 3.025 2.350 3.035 2.600 ;
        RECT 3.035 2.360 3.045 2.610 ;
        RECT 3.045 2.370 3.055 2.620 ;
        RECT 3.055 2.380 3.065 2.630 ;
        RECT 3.065 2.390 3.075 2.640 ;
        RECT 3.075 2.400 3.085 2.650 ;
        RECT 3.085 2.410 3.095 2.660 ;
        RECT 3.095 2.420 3.105 2.670 ;
        RECT 3.105 2.430 3.115 2.680 ;
        RECT 3.115 2.440 3.125 2.690 ;
        RECT 3.125 2.450 3.135 2.700 ;
        RECT 3.135 2.460 3.145 2.710 ;
        RECT 3.145 2.470 3.155 2.720 ;
        RECT 3.155 2.480 3.165 2.730 ;
        RECT 3.165 2.490 3.175 2.740 ;
        RECT 3.175 2.500 3.185 2.750 ;
        RECT 3.185 2.510 3.195 2.760 ;
        RECT 3.195 2.520 3.205 2.770 ;
        RECT 3.205 2.530 3.215 2.780 ;
        RECT 3.215 2.540 3.225 2.790 ;
        RECT 3.225 2.550 3.235 2.800 ;
        RECT 3.235 2.560 3.245 2.810 ;
        RECT 3.245 2.570 3.255 2.820 ;
        RECT 3.255 2.580 3.265 2.830 ;
        RECT 3.265 2.590 3.275 2.840 ;
        RECT 3.275 2.595 3.281 2.849 ;
        RECT 2.935 2.340 2.945 2.510 ;
        RECT 2.945 2.340 2.955 2.520 ;
        RECT 2.955 2.340 2.965 2.530 ;
        RECT 2.965 2.340 2.975 2.540 ;
        RECT 2.975 2.340 2.985 2.550 ;
        RECT 2.985 2.340 2.995 2.560 ;
        RECT 2.995 2.340 3.005 2.570 ;
        RECT 3.005 2.340 3.015 2.580 ;
        RECT 3.015 2.340 3.025 2.590 ;
        RECT 2.105 2.340 2.115 2.530 ;
        RECT 2.115 2.340 2.125 2.520 ;
        RECT 2.125 2.340 2.135 2.510 ;
        RECT 2.015 2.370 2.025 2.540 ;
        RECT 2.025 2.360 2.035 2.540 ;
        RECT 2.035 2.350 2.045 2.540 ;
        RECT 5.630 1.805 5.700 1.995 ;
        RECT 5.620 1.815 5.806 1.889 ;
        RECT 5.400 1.825 5.700 1.995 ;
        RECT 5.400 1.825 5.710 1.985 ;
        RECT 5.400 1.825 5.720 1.975 ;
        RECT 5.400 1.825 5.730 1.965 ;
        RECT 5.400 1.825 5.740 1.955 ;
        RECT 5.400 1.825 5.750 1.945 ;
        RECT 5.400 1.825 5.760 1.935 ;
        RECT 5.400 1.825 5.770 1.925 ;
        RECT 5.400 1.825 5.780 1.915 ;
        RECT 5.400 1.825 5.790 1.905 ;
        RECT 5.400 1.825 5.800 1.895 ;
        RECT 5.635 1.255 5.806 1.889 ;
        RECT 6.630 1.105 6.865 1.425 ;
        RECT 5.635 1.255 6.865 1.425 ;
        RECT 6.695 1.105 6.865 2.280 ;
        RECT 6.630 1.105 6.930 1.275 ;
        RECT 4.965 1.170 5.135 2.495 ;
        RECT 5.285 0.905 5.455 1.340 ;
        RECT 4.965 1.170 5.455 1.340 ;
        RECT 4.965 2.325 5.520 2.495 ;
        RECT 5.285 0.905 6.310 1.075 ;
        RECT 6.570 0.735 7.090 0.905 ;
        RECT 6.480 0.735 6.490 0.985 ;
        RECT 6.490 0.735 6.500 0.975 ;
        RECT 6.500 0.735 6.510 0.965 ;
        RECT 6.510 0.735 6.520 0.955 ;
        RECT 6.520 0.735 6.530 0.945 ;
        RECT 6.530 0.735 6.540 0.935 ;
        RECT 6.540 0.735 6.550 0.925 ;
        RECT 6.550 0.735 6.560 0.915 ;
        RECT 6.560 0.735 6.570 0.905 ;
        RECT 6.400 0.815 6.410 1.065 ;
        RECT 6.410 0.805 6.420 1.055 ;
        RECT 6.420 0.795 6.430 1.045 ;
        RECT 6.430 0.785 6.440 1.035 ;
        RECT 6.440 0.775 6.450 1.025 ;
        RECT 6.450 0.765 6.460 1.015 ;
        RECT 6.460 0.755 6.470 1.005 ;
        RECT 6.470 0.745 6.480 0.995 ;
        RECT 6.310 0.905 6.320 1.075 ;
        RECT 6.320 0.895 6.330 1.075 ;
        RECT 6.330 0.885 6.340 1.075 ;
        RECT 6.340 0.875 6.350 1.075 ;
        RECT 6.350 0.865 6.360 1.075 ;
        RECT 6.360 0.855 6.370 1.075 ;
        RECT 6.370 0.845 6.380 1.075 ;
        RECT 6.380 0.835 6.390 1.075 ;
        RECT 6.390 0.825 6.400 1.075 ;
        RECT 7.205 1.060 7.375 2.280 ;
        RECT 7.205 1.590 8.035 1.760 ;
        RECT 7.865 1.525 8.035 1.825 ;
  END 
END MUX4HDMXHT

MACRO MUX4HDLXHT
  CLASS  CORE ;
  FOREIGN MUX4HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.610 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.240 2.500 6.750 2.830 ;
    END
  END S1
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.175 1.890 4.420 2.440 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.485 1.730 2.830 2.140 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.060 0.920 2.525 1.450 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 1.060 1.140 1.665 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.665 ;
        RECT 2.375 -0.300 2.675 0.740 ;
        RECT 4.380 -0.300 4.680 0.680 ;
        RECT 5.930 -0.300 6.230 0.725 ;
        RECT 7.590 -0.300 7.890 0.715 ;
        RECT 0.000 -0.300 8.610 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.215 1.060 8.385 2.360 ;
        RECT 7.810 2.150 8.385 2.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.675 3.040 0.975 3.990 ;
        RECT 2.385 3.040 2.685 3.990 ;
        RECT 4.380 3.025 4.680 3.990 ;
        RECT 6.080 3.025 6.380 3.990 ;
        RECT 7.590 2.715 7.890 3.990 ;
        RECT 0.000 3.390 8.610 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.500 1.910 0.680 2.420 ;
        RECT 0.500 2.000 0.780 2.420 ;
        RECT 0.500 2.000 1.955 2.170 ;
        RECT 3.300 1.155 3.790 1.325 ;
        RECT 3.620 1.155 3.790 2.125 ;
        RECT 3.620 1.955 3.920 2.125 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.105 1.075 0.275 2.860 ;
        RECT 0.105 1.075 0.405 1.245 ;
        RECT 0.105 2.600 0.405 2.860 ;
        RECT 1.165 2.690 1.335 3.030 ;
        RECT 0.105 2.690 1.335 2.860 ;
        RECT 1.165 2.860 2.045 3.030 ;
        RECT 2.305 2.690 2.765 2.860 ;
        RECT 3.030 2.865 3.035 3.210 ;
        RECT 3.030 3.040 3.325 3.210 ;
        RECT 2.865 2.710 2.875 3.210 ;
        RECT 2.875 2.720 2.885 3.210 ;
        RECT 2.885 2.730 2.895 3.210 ;
        RECT 2.895 2.740 2.905 3.210 ;
        RECT 2.905 2.750 2.915 3.210 ;
        RECT 2.915 2.760 2.925 3.210 ;
        RECT 2.925 2.770 2.935 3.210 ;
        RECT 2.935 2.780 2.945 3.210 ;
        RECT 2.945 2.790 2.955 3.210 ;
        RECT 2.955 2.800 2.965 3.210 ;
        RECT 2.965 2.810 2.975 3.210 ;
        RECT 2.975 2.820 2.985 3.210 ;
        RECT 2.985 2.830 2.995 3.210 ;
        RECT 2.995 2.840 3.005 3.210 ;
        RECT 3.005 2.850 3.015 3.210 ;
        RECT 3.015 2.860 3.025 3.210 ;
        RECT 3.025 2.865 3.031 3.209 ;
        RECT 2.855 2.700 2.865 2.950 ;
        RECT 2.765 2.690 2.775 2.860 ;
        RECT 2.775 2.690 2.785 2.870 ;
        RECT 2.785 2.690 2.795 2.880 ;
        RECT 2.795 2.690 2.805 2.890 ;
        RECT 2.805 2.690 2.815 2.900 ;
        RECT 2.815 2.690 2.825 2.910 ;
        RECT 2.825 2.690 2.835 2.920 ;
        RECT 2.835 2.690 2.845 2.930 ;
        RECT 2.845 2.690 2.855 2.940 ;
        RECT 2.215 2.690 2.225 2.940 ;
        RECT 2.225 2.690 2.235 2.930 ;
        RECT 2.235 2.690 2.245 2.920 ;
        RECT 2.245 2.690 2.255 2.910 ;
        RECT 2.255 2.690 2.265 2.900 ;
        RECT 2.265 2.690 2.275 2.890 ;
        RECT 2.275 2.690 2.285 2.880 ;
        RECT 2.285 2.690 2.295 2.870 ;
        RECT 2.295 2.690 2.305 2.860 ;
        RECT 2.135 2.770 2.145 3.020 ;
        RECT 2.145 2.760 2.155 3.010 ;
        RECT 2.155 2.750 2.165 3.000 ;
        RECT 2.165 2.740 2.175 2.990 ;
        RECT 2.175 2.730 2.185 2.980 ;
        RECT 2.185 2.720 2.195 2.970 ;
        RECT 2.195 2.710 2.205 2.960 ;
        RECT 2.205 2.700 2.215 2.950 ;
        RECT 2.045 2.860 2.055 3.030 ;
        RECT 2.055 2.850 2.065 3.030 ;
        RECT 2.065 2.840 2.075 3.030 ;
        RECT 2.075 2.830 2.085 3.030 ;
        RECT 2.085 2.820 2.095 3.030 ;
        RECT 2.095 2.810 2.105 3.030 ;
        RECT 2.105 2.800 2.115 3.030 ;
        RECT 2.115 2.790 2.125 3.030 ;
        RECT 2.125 2.780 2.135 3.030 ;
        RECT 3.220 1.505 3.270 1.675 ;
        RECT 3.530 2.325 3.740 2.495 ;
        RECT 3.120 0.785 4.140 0.955 ;
        RECT 3.970 0.785 4.140 1.325 ;
        RECT 3.970 1.155 4.745 1.325 ;
        RECT 4.575 1.155 4.745 1.710 ;
        RECT 3.440 2.245 3.450 2.495 ;
        RECT 3.450 2.255 3.460 2.495 ;
        RECT 3.460 2.265 3.470 2.495 ;
        RECT 3.470 2.275 3.480 2.495 ;
        RECT 3.480 2.285 3.490 2.495 ;
        RECT 3.490 2.295 3.500 2.495 ;
        RECT 3.500 2.305 3.510 2.495 ;
        RECT 3.510 2.315 3.520 2.495 ;
        RECT 3.520 2.325 3.530 2.495 ;
        RECT 3.270 1.505 3.280 2.325 ;
        RECT 3.280 1.505 3.290 2.335 ;
        RECT 3.290 1.505 3.300 2.345 ;
        RECT 3.300 1.505 3.310 2.355 ;
        RECT 3.310 1.505 3.320 2.365 ;
        RECT 3.320 1.505 3.330 2.375 ;
        RECT 3.330 1.505 3.340 2.385 ;
        RECT 3.340 1.505 3.350 2.395 ;
        RECT 3.350 1.505 3.360 2.405 ;
        RECT 3.360 1.505 3.370 2.415 ;
        RECT 3.370 1.505 3.380 2.425 ;
        RECT 3.380 1.505 3.390 2.435 ;
        RECT 3.390 1.505 3.400 2.445 ;
        RECT 3.400 1.505 3.410 2.455 ;
        RECT 3.410 1.505 3.420 2.465 ;
        RECT 3.420 1.505 3.430 2.475 ;
        RECT 3.430 1.505 3.440 2.485 ;
        RECT 3.130 1.425 3.140 1.675 ;
        RECT 3.140 1.435 3.150 1.675 ;
        RECT 3.150 1.445 3.160 1.675 ;
        RECT 3.160 1.455 3.170 1.675 ;
        RECT 3.170 1.465 3.180 1.675 ;
        RECT 3.180 1.475 3.190 1.675 ;
        RECT 3.190 1.485 3.200 1.675 ;
        RECT 3.200 1.495 3.210 1.675 ;
        RECT 3.210 1.505 3.220 1.675 ;
        RECT 3.120 1.415 3.130 1.665 ;
        RECT 2.950 0.785 2.960 1.495 ;
        RECT 2.960 0.785 2.970 1.505 ;
        RECT 2.970 0.785 2.980 1.515 ;
        RECT 2.980 0.785 2.990 1.525 ;
        RECT 2.990 0.785 3.000 1.535 ;
        RECT 3.000 0.785 3.010 1.545 ;
        RECT 3.010 0.785 3.020 1.555 ;
        RECT 3.020 0.785 3.030 1.565 ;
        RECT 3.030 0.785 3.040 1.575 ;
        RECT 3.040 0.785 3.050 1.585 ;
        RECT 3.050 0.785 3.060 1.595 ;
        RECT 3.060 0.785 3.070 1.605 ;
        RECT 3.070 0.785 3.080 1.615 ;
        RECT 3.080 0.785 3.090 1.625 ;
        RECT 3.090 0.785 3.100 1.635 ;
        RECT 3.100 0.785 3.110 1.645 ;
        RECT 3.110 0.785 3.120 1.655 ;
        RECT 1.520 0.720 1.690 1.820 ;
        RECT 1.515 2.370 2.015 2.540 ;
        RECT 2.045 2.340 2.105 2.540 ;
        RECT 1.520 1.650 2.305 1.820 ;
        RECT 2.135 1.650 2.305 2.510 ;
        RECT 2.135 2.340 2.935 2.510 ;
        RECT 3.360 2.675 3.595 2.855 ;
        RECT 3.360 2.675 5.800 2.845 ;
        RECT 6.105 1.610 6.165 2.190 ;
        RECT 5.995 1.610 6.005 2.290 ;
        RECT 6.005 1.610 6.015 2.280 ;
        RECT 6.015 1.610 6.025 2.270 ;
        RECT 6.025 1.610 6.035 2.260 ;
        RECT 6.035 1.610 6.045 2.250 ;
        RECT 6.045 1.610 6.055 2.240 ;
        RECT 6.055 1.610 6.065 2.230 ;
        RECT 6.065 1.610 6.075 2.220 ;
        RECT 6.075 1.610 6.085 2.210 ;
        RECT 6.085 1.610 6.095 2.200 ;
        RECT 6.095 1.610 6.105 2.190 ;
        RECT 5.970 2.065 5.980 2.835 ;
        RECT 5.980 2.055 5.990 2.825 ;
        RECT 5.990 2.045 5.996 2.819 ;
        RECT 5.825 2.210 5.835 2.844 ;
        RECT 5.835 2.200 5.845 2.844 ;
        RECT 5.845 2.190 5.855 2.844 ;
        RECT 5.855 2.180 5.865 2.844 ;
        RECT 5.865 2.170 5.875 2.844 ;
        RECT 5.875 2.160 5.885 2.844 ;
        RECT 5.885 2.150 5.895 2.844 ;
        RECT 5.895 2.140 5.905 2.844 ;
        RECT 5.905 2.130 5.915 2.844 ;
        RECT 5.915 2.120 5.925 2.844 ;
        RECT 5.925 2.110 5.935 2.844 ;
        RECT 5.935 2.100 5.945 2.844 ;
        RECT 5.945 2.090 5.955 2.844 ;
        RECT 5.955 2.080 5.965 2.844 ;
        RECT 5.965 2.070 5.971 2.844 ;
        RECT 5.800 2.675 5.810 2.845 ;
        RECT 5.810 2.665 5.820 2.845 ;
        RECT 5.820 2.655 5.826 2.845 ;
        RECT 3.280 2.605 3.290 2.855 ;
        RECT 3.290 2.615 3.300 2.855 ;
        RECT 3.300 2.625 3.310 2.855 ;
        RECT 3.310 2.635 3.320 2.855 ;
        RECT 3.320 2.645 3.330 2.855 ;
        RECT 3.330 2.655 3.340 2.855 ;
        RECT 3.340 2.665 3.350 2.855 ;
        RECT 3.350 2.675 3.360 2.855 ;
        RECT 3.025 2.350 3.035 2.600 ;
        RECT 3.035 2.360 3.045 2.610 ;
        RECT 3.045 2.370 3.055 2.620 ;
        RECT 3.055 2.380 3.065 2.630 ;
        RECT 3.065 2.390 3.075 2.640 ;
        RECT 3.075 2.400 3.085 2.650 ;
        RECT 3.085 2.410 3.095 2.660 ;
        RECT 3.095 2.420 3.105 2.670 ;
        RECT 3.105 2.430 3.115 2.680 ;
        RECT 3.115 2.440 3.125 2.690 ;
        RECT 3.125 2.450 3.135 2.700 ;
        RECT 3.135 2.460 3.145 2.710 ;
        RECT 3.145 2.470 3.155 2.720 ;
        RECT 3.155 2.480 3.165 2.730 ;
        RECT 3.165 2.490 3.175 2.740 ;
        RECT 3.175 2.500 3.185 2.750 ;
        RECT 3.185 2.510 3.195 2.760 ;
        RECT 3.195 2.520 3.205 2.770 ;
        RECT 3.205 2.530 3.215 2.780 ;
        RECT 3.215 2.540 3.225 2.790 ;
        RECT 3.225 2.550 3.235 2.800 ;
        RECT 3.235 2.560 3.245 2.810 ;
        RECT 3.245 2.570 3.255 2.820 ;
        RECT 3.255 2.580 3.265 2.830 ;
        RECT 3.265 2.590 3.275 2.840 ;
        RECT 3.275 2.595 3.281 2.849 ;
        RECT 2.935 2.340 2.945 2.510 ;
        RECT 2.945 2.340 2.955 2.520 ;
        RECT 2.955 2.340 2.965 2.530 ;
        RECT 2.965 2.340 2.975 2.540 ;
        RECT 2.975 2.340 2.985 2.550 ;
        RECT 2.985 2.340 2.995 2.560 ;
        RECT 2.995 2.340 3.005 2.570 ;
        RECT 3.005 2.340 3.015 2.580 ;
        RECT 3.015 2.340 3.025 2.590 ;
        RECT 2.105 2.340 2.115 2.530 ;
        RECT 2.115 2.340 2.125 2.520 ;
        RECT 2.125 2.340 2.135 2.510 ;
        RECT 2.015 2.370 2.025 2.540 ;
        RECT 2.025 2.360 2.035 2.540 ;
        RECT 2.035 2.350 2.045 2.540 ;
        RECT 5.630 1.805 5.700 1.995 ;
        RECT 5.620 1.815 5.806 1.889 ;
        RECT 5.400 1.825 5.700 1.995 ;
        RECT 5.400 1.825 5.710 1.985 ;
        RECT 5.400 1.825 5.720 1.975 ;
        RECT 5.400 1.825 5.730 1.965 ;
        RECT 5.400 1.825 5.740 1.955 ;
        RECT 5.400 1.825 5.750 1.945 ;
        RECT 5.400 1.825 5.760 1.935 ;
        RECT 5.400 1.825 5.770 1.925 ;
        RECT 5.400 1.825 5.780 1.915 ;
        RECT 5.400 1.825 5.790 1.905 ;
        RECT 5.400 1.825 5.800 1.895 ;
        RECT 5.635 1.255 5.806 1.889 ;
        RECT 6.630 1.105 6.865 1.425 ;
        RECT 5.635 1.255 6.865 1.425 ;
        RECT 6.695 1.105 6.865 2.280 ;
        RECT 6.630 1.105 6.930 1.275 ;
        RECT 4.965 1.170 5.135 2.495 ;
        RECT 5.285 0.905 5.455 1.340 ;
        RECT 4.965 1.170 5.455 1.340 ;
        RECT 4.965 2.325 5.520 2.495 ;
        RECT 5.285 0.905 6.310 1.075 ;
        RECT 6.595 0.710 7.410 0.880 ;
        RECT 6.505 0.710 6.515 0.960 ;
        RECT 6.515 0.710 6.525 0.950 ;
        RECT 6.525 0.710 6.535 0.940 ;
        RECT 6.535 0.710 6.545 0.930 ;
        RECT 6.545 0.710 6.555 0.920 ;
        RECT 6.555 0.710 6.565 0.910 ;
        RECT 6.565 0.710 6.575 0.900 ;
        RECT 6.575 0.710 6.585 0.890 ;
        RECT 6.585 0.710 6.595 0.880 ;
        RECT 6.400 0.815 6.410 1.065 ;
        RECT 6.410 0.805 6.420 1.055 ;
        RECT 6.420 0.795 6.430 1.045 ;
        RECT 6.430 0.785 6.440 1.035 ;
        RECT 6.440 0.775 6.450 1.025 ;
        RECT 6.450 0.765 6.460 1.015 ;
        RECT 6.460 0.755 6.470 1.005 ;
        RECT 6.470 0.745 6.480 0.995 ;
        RECT 6.480 0.735 6.490 0.985 ;
        RECT 6.490 0.725 6.500 0.975 ;
        RECT 6.500 0.715 6.506 0.969 ;
        RECT 6.310 0.905 6.320 1.075 ;
        RECT 6.320 0.895 6.330 1.075 ;
        RECT 6.330 0.885 6.340 1.075 ;
        RECT 6.340 0.875 6.350 1.075 ;
        RECT 6.350 0.865 6.360 1.075 ;
        RECT 6.360 0.855 6.370 1.075 ;
        RECT 6.370 0.845 6.380 1.075 ;
        RECT 6.380 0.835 6.390 1.075 ;
        RECT 6.390 0.825 6.400 1.075 ;
        RECT 7.205 1.060 7.375 2.280 ;
        RECT 7.205 1.630 8.035 1.800 ;
        RECT 7.865 1.525 8.035 1.825 ;
  END 
END MUX4HDLXHT

MACRO MUX4HD2XHT
  CLASS  CORE ;
  FOREIGN MUX4HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.020 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.190 2.500 6.700 2.830 ;
    END
  END S1
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.175 1.890 4.420 2.440 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.485 1.730 2.830 2.140 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.060 0.920 2.525 1.385 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 1.060 1.140 1.665 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.665 ;
        RECT 2.375 -0.300 2.675 0.740 ;
        RECT 4.360 -0.300 4.660 0.680 ;
        RECT 5.860 -0.300 6.160 0.705 ;
        RECT 7.635 -0.300 7.805 1.220 ;
        RECT 8.610 -0.300 8.910 1.055 ;
        RECT 0.000 -0.300 9.020 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.790 2.150 8.390 2.360 ;
        RECT 8.155 0.720 8.390 3.090 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.675 3.040 0.975 3.990 ;
        RECT 2.385 3.040 2.685 3.990 ;
        RECT 4.360 3.025 4.660 3.990 ;
        RECT 6.030 3.025 6.330 3.990 ;
        RECT 7.540 2.975 7.840 3.990 ;
        RECT 8.610 2.295 8.910 3.990 ;
        RECT 0.000 3.390 9.020 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.910 0.680 2.420 ;
        RECT 0.510 2.000 0.720 2.420 ;
        RECT 0.510 2.000 1.955 2.170 ;
        RECT 3.300 1.155 3.790 1.325 ;
        RECT 3.620 1.155 3.790 2.125 ;
        RECT 3.620 1.955 3.920 2.125 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.105 1.075 0.275 2.860 ;
        RECT 0.105 1.075 0.405 1.245 ;
        RECT 0.105 2.600 0.405 2.860 ;
        RECT 1.165 2.690 1.335 3.030 ;
        RECT 0.105 2.690 1.335 2.860 ;
        RECT 1.165 2.860 2.045 3.030 ;
        RECT 2.305 2.690 2.765 2.860 ;
        RECT 3.030 2.865 3.035 3.210 ;
        RECT 3.030 3.040 3.325 3.210 ;
        RECT 2.865 2.710 2.875 3.210 ;
        RECT 2.875 2.720 2.885 3.210 ;
        RECT 2.885 2.730 2.895 3.210 ;
        RECT 2.895 2.740 2.905 3.210 ;
        RECT 2.905 2.750 2.915 3.210 ;
        RECT 2.915 2.760 2.925 3.210 ;
        RECT 2.925 2.770 2.935 3.210 ;
        RECT 2.935 2.780 2.945 3.210 ;
        RECT 2.945 2.790 2.955 3.210 ;
        RECT 2.955 2.800 2.965 3.210 ;
        RECT 2.965 2.810 2.975 3.210 ;
        RECT 2.975 2.820 2.985 3.210 ;
        RECT 2.985 2.830 2.995 3.210 ;
        RECT 2.995 2.840 3.005 3.210 ;
        RECT 3.005 2.850 3.015 3.210 ;
        RECT 3.015 2.860 3.025 3.210 ;
        RECT 3.025 2.865 3.031 3.209 ;
        RECT 2.855 2.700 2.865 2.950 ;
        RECT 2.765 2.690 2.775 2.860 ;
        RECT 2.775 2.690 2.785 2.870 ;
        RECT 2.785 2.690 2.795 2.880 ;
        RECT 2.795 2.690 2.805 2.890 ;
        RECT 2.805 2.690 2.815 2.900 ;
        RECT 2.815 2.690 2.825 2.910 ;
        RECT 2.825 2.690 2.835 2.920 ;
        RECT 2.835 2.690 2.845 2.930 ;
        RECT 2.845 2.690 2.855 2.940 ;
        RECT 2.215 2.690 2.225 2.940 ;
        RECT 2.225 2.690 2.235 2.930 ;
        RECT 2.235 2.690 2.245 2.920 ;
        RECT 2.245 2.690 2.255 2.910 ;
        RECT 2.255 2.690 2.265 2.900 ;
        RECT 2.265 2.690 2.275 2.890 ;
        RECT 2.275 2.690 2.285 2.880 ;
        RECT 2.285 2.690 2.295 2.870 ;
        RECT 2.295 2.690 2.305 2.860 ;
        RECT 2.135 2.770 2.145 3.020 ;
        RECT 2.145 2.760 2.155 3.010 ;
        RECT 2.155 2.750 2.165 3.000 ;
        RECT 2.165 2.740 2.175 2.990 ;
        RECT 2.175 2.730 2.185 2.980 ;
        RECT 2.185 2.720 2.195 2.970 ;
        RECT 2.195 2.710 2.205 2.960 ;
        RECT 2.205 2.700 2.215 2.950 ;
        RECT 2.045 2.860 2.055 3.030 ;
        RECT 2.055 2.850 2.065 3.030 ;
        RECT 2.065 2.840 2.075 3.030 ;
        RECT 2.075 2.830 2.085 3.030 ;
        RECT 2.085 2.820 2.095 3.030 ;
        RECT 2.095 2.810 2.105 3.030 ;
        RECT 2.105 2.800 2.115 3.030 ;
        RECT 2.115 2.790 2.125 3.030 ;
        RECT 2.125 2.780 2.135 3.030 ;
        RECT 3.220 1.505 3.270 1.675 ;
        RECT 3.530 2.325 3.740 2.495 ;
        RECT 3.120 0.785 4.140 0.955 ;
        RECT 3.970 0.785 4.140 1.325 ;
        RECT 3.970 1.155 4.705 1.325 ;
        RECT 4.535 1.155 4.705 1.710 ;
        RECT 3.440 2.245 3.450 2.495 ;
        RECT 3.450 2.255 3.460 2.495 ;
        RECT 3.460 2.265 3.470 2.495 ;
        RECT 3.470 2.275 3.480 2.495 ;
        RECT 3.480 2.285 3.490 2.495 ;
        RECT 3.490 2.295 3.500 2.495 ;
        RECT 3.500 2.305 3.510 2.495 ;
        RECT 3.510 2.315 3.520 2.495 ;
        RECT 3.520 2.325 3.530 2.495 ;
        RECT 3.270 1.505 3.280 2.325 ;
        RECT 3.280 1.505 3.290 2.335 ;
        RECT 3.290 1.505 3.300 2.345 ;
        RECT 3.300 1.505 3.310 2.355 ;
        RECT 3.310 1.505 3.320 2.365 ;
        RECT 3.320 1.505 3.330 2.375 ;
        RECT 3.330 1.505 3.340 2.385 ;
        RECT 3.340 1.505 3.350 2.395 ;
        RECT 3.350 1.505 3.360 2.405 ;
        RECT 3.360 1.505 3.370 2.415 ;
        RECT 3.370 1.505 3.380 2.425 ;
        RECT 3.380 1.505 3.390 2.435 ;
        RECT 3.390 1.505 3.400 2.445 ;
        RECT 3.400 1.505 3.410 2.455 ;
        RECT 3.410 1.505 3.420 2.465 ;
        RECT 3.420 1.505 3.430 2.475 ;
        RECT 3.430 1.505 3.440 2.485 ;
        RECT 3.130 1.425 3.140 1.675 ;
        RECT 3.140 1.435 3.150 1.675 ;
        RECT 3.150 1.445 3.160 1.675 ;
        RECT 3.160 1.455 3.170 1.675 ;
        RECT 3.170 1.465 3.180 1.675 ;
        RECT 3.180 1.475 3.190 1.675 ;
        RECT 3.190 1.485 3.200 1.675 ;
        RECT 3.200 1.495 3.210 1.675 ;
        RECT 3.210 1.505 3.220 1.675 ;
        RECT 3.120 1.415 3.130 1.665 ;
        RECT 2.950 0.785 2.960 1.495 ;
        RECT 2.960 0.785 2.970 1.505 ;
        RECT 2.970 0.785 2.980 1.515 ;
        RECT 2.980 0.785 2.990 1.525 ;
        RECT 2.990 0.785 3.000 1.535 ;
        RECT 3.000 0.785 3.010 1.545 ;
        RECT 3.010 0.785 3.020 1.555 ;
        RECT 3.020 0.785 3.030 1.565 ;
        RECT 3.030 0.785 3.040 1.575 ;
        RECT 3.040 0.785 3.050 1.585 ;
        RECT 3.050 0.785 3.060 1.595 ;
        RECT 3.060 0.785 3.070 1.605 ;
        RECT 3.070 0.785 3.080 1.615 ;
        RECT 3.080 0.785 3.090 1.625 ;
        RECT 3.090 0.785 3.100 1.635 ;
        RECT 3.100 0.785 3.110 1.645 ;
        RECT 3.110 0.785 3.120 1.655 ;
        RECT 1.520 0.720 1.690 1.820 ;
        RECT 1.515 2.370 2.015 2.540 ;
        RECT 1.520 1.650 2.035 1.820 ;
        RECT 2.045 2.340 2.105 2.540 ;
        RECT 2.275 1.800 2.305 2.510 ;
        RECT 2.275 2.340 2.935 2.510 ;
        RECT 3.360 2.675 5.800 2.845 ;
        RECT 5.945 1.610 5.970 2.845 ;
        RECT 6.105 1.610 6.115 2.190 ;
        RECT 5.995 1.610 6.005 2.290 ;
        RECT 6.005 1.610 6.015 2.280 ;
        RECT 6.015 1.610 6.025 2.270 ;
        RECT 6.025 1.610 6.035 2.260 ;
        RECT 6.035 1.610 6.045 2.250 ;
        RECT 6.045 1.610 6.055 2.240 ;
        RECT 6.055 1.610 6.065 2.230 ;
        RECT 6.065 1.610 6.075 2.220 ;
        RECT 6.075 1.610 6.085 2.210 ;
        RECT 6.085 1.610 6.095 2.200 ;
        RECT 6.095 1.610 6.105 2.190 ;
        RECT 5.970 1.610 5.980 2.834 ;
        RECT 5.980 1.610 5.990 2.824 ;
        RECT 5.990 1.610 5.996 2.820 ;
        RECT 5.825 2.210 5.835 2.844 ;
        RECT 5.835 2.200 5.845 2.844 ;
        RECT 5.845 2.190 5.855 2.844 ;
        RECT 5.855 2.180 5.865 2.844 ;
        RECT 5.865 2.170 5.875 2.844 ;
        RECT 5.875 2.160 5.885 2.844 ;
        RECT 5.885 2.150 5.895 2.844 ;
        RECT 5.895 2.140 5.905 2.844 ;
        RECT 5.905 2.130 5.915 2.844 ;
        RECT 5.915 2.120 5.925 2.844 ;
        RECT 5.925 2.110 5.935 2.844 ;
        RECT 5.935 2.100 5.945 2.844 ;
        RECT 5.800 2.675 5.810 2.845 ;
        RECT 5.810 2.665 5.820 2.845 ;
        RECT 5.820 2.655 5.826 2.845 ;
        RECT 3.270 2.595 3.280 2.845 ;
        RECT 3.280 2.605 3.290 2.845 ;
        RECT 3.290 2.615 3.300 2.845 ;
        RECT 3.300 2.625 3.310 2.845 ;
        RECT 3.310 2.635 3.320 2.845 ;
        RECT 3.320 2.645 3.330 2.845 ;
        RECT 3.330 2.655 3.340 2.845 ;
        RECT 3.340 2.665 3.350 2.845 ;
        RECT 3.350 2.675 3.360 2.845 ;
        RECT 3.025 2.350 3.035 2.600 ;
        RECT 3.035 2.360 3.045 2.610 ;
        RECT 3.045 2.370 3.055 2.620 ;
        RECT 3.055 2.380 3.065 2.630 ;
        RECT 3.065 2.390 3.075 2.640 ;
        RECT 3.075 2.400 3.085 2.650 ;
        RECT 3.085 2.410 3.095 2.660 ;
        RECT 3.095 2.420 3.105 2.670 ;
        RECT 3.105 2.430 3.115 2.680 ;
        RECT 3.115 2.440 3.125 2.690 ;
        RECT 3.125 2.450 3.135 2.700 ;
        RECT 3.135 2.460 3.145 2.710 ;
        RECT 3.145 2.470 3.155 2.720 ;
        RECT 3.155 2.480 3.165 2.730 ;
        RECT 3.165 2.490 3.175 2.740 ;
        RECT 3.175 2.500 3.185 2.750 ;
        RECT 3.185 2.510 3.195 2.760 ;
        RECT 3.195 2.520 3.205 2.770 ;
        RECT 3.205 2.530 3.215 2.780 ;
        RECT 3.215 2.540 3.225 2.790 ;
        RECT 3.225 2.550 3.235 2.800 ;
        RECT 3.235 2.560 3.245 2.810 ;
        RECT 3.245 2.570 3.255 2.820 ;
        RECT 3.255 2.580 3.265 2.830 ;
        RECT 3.265 2.585 3.271 2.839 ;
        RECT 2.935 2.340 2.945 2.510 ;
        RECT 2.945 2.340 2.955 2.520 ;
        RECT 2.955 2.340 2.965 2.530 ;
        RECT 2.965 2.340 2.975 2.540 ;
        RECT 2.975 2.340 2.985 2.550 ;
        RECT 2.985 2.340 2.995 2.560 ;
        RECT 2.995 2.340 3.005 2.570 ;
        RECT 3.005 2.340 3.015 2.580 ;
        RECT 3.015 2.340 3.025 2.590 ;
        RECT 2.135 1.670 2.145 2.510 ;
        RECT 2.145 1.680 2.155 2.510 ;
        RECT 2.155 1.690 2.165 2.510 ;
        RECT 2.165 1.700 2.175 2.510 ;
        RECT 2.175 1.710 2.185 2.510 ;
        RECT 2.185 1.720 2.195 2.510 ;
        RECT 2.195 1.730 2.205 2.510 ;
        RECT 2.205 1.740 2.215 2.510 ;
        RECT 2.215 1.750 2.225 2.510 ;
        RECT 2.225 1.760 2.235 2.510 ;
        RECT 2.235 1.770 2.245 2.510 ;
        RECT 2.245 1.780 2.255 2.510 ;
        RECT 2.255 1.790 2.265 2.510 ;
        RECT 2.265 1.800 2.275 2.510 ;
        RECT 2.125 1.660 2.135 1.910 ;
        RECT 2.105 2.340 2.115 2.530 ;
        RECT 2.115 2.340 2.125 2.520 ;
        RECT 2.125 2.340 2.135 2.510 ;
        RECT 2.035 1.650 2.045 1.820 ;
        RECT 2.045 1.650 2.055 1.830 ;
        RECT 2.055 1.650 2.065 1.840 ;
        RECT 2.065 1.650 2.075 1.850 ;
        RECT 2.075 1.650 2.085 1.860 ;
        RECT 2.085 1.650 2.095 1.870 ;
        RECT 2.095 1.650 2.105 1.880 ;
        RECT 2.105 1.650 2.115 1.890 ;
        RECT 2.115 1.650 2.125 1.900 ;
        RECT 2.015 2.370 2.025 2.540 ;
        RECT 2.025 2.360 2.035 2.540 ;
        RECT 2.035 2.350 2.045 2.540 ;
        RECT 5.580 1.805 5.650 1.995 ;
        RECT 5.570 1.815 5.756 1.889 ;
        RECT 5.350 1.825 5.650 1.995 ;
        RECT 5.350 1.825 5.660 1.985 ;
        RECT 5.350 1.825 5.670 1.975 ;
        RECT 5.350 1.825 5.680 1.965 ;
        RECT 5.350 1.825 5.690 1.955 ;
        RECT 5.350 1.825 5.700 1.945 ;
        RECT 5.350 1.825 5.710 1.935 ;
        RECT 5.350 1.825 5.720 1.925 ;
        RECT 5.350 1.825 5.730 1.915 ;
        RECT 5.350 1.825 5.740 1.905 ;
        RECT 5.350 1.825 5.750 1.895 ;
        RECT 5.585 1.255 5.756 1.889 ;
        RECT 5.585 1.255 6.815 1.425 ;
        RECT 6.605 1.040 6.775 1.425 ;
        RECT 6.645 1.225 6.815 2.280 ;
        RECT 4.915 1.170 5.085 2.495 ;
        RECT 5.235 0.905 5.405 1.340 ;
        RECT 4.915 1.170 5.405 1.340 ;
        RECT 4.915 2.325 5.470 2.495 ;
        RECT 5.235 0.905 6.220 1.075 ;
        RECT 6.525 0.690 6.980 0.860 ;
        RECT 6.435 0.690 6.445 0.940 ;
        RECT 6.445 0.690 6.455 0.930 ;
        RECT 6.455 0.690 6.465 0.920 ;
        RECT 6.465 0.690 6.475 0.910 ;
        RECT 6.475 0.690 6.485 0.900 ;
        RECT 6.485 0.690 6.495 0.890 ;
        RECT 6.495 0.690 6.505 0.880 ;
        RECT 6.505 0.690 6.515 0.870 ;
        RECT 6.515 0.690 6.525 0.860 ;
        RECT 6.310 0.815 6.320 1.065 ;
        RECT 6.320 0.805 6.330 1.055 ;
        RECT 6.330 0.795 6.340 1.045 ;
        RECT 6.340 0.785 6.350 1.035 ;
        RECT 6.350 0.775 6.360 1.025 ;
        RECT 6.360 0.765 6.370 1.015 ;
        RECT 6.370 0.755 6.380 1.005 ;
        RECT 6.380 0.745 6.390 0.995 ;
        RECT 6.390 0.735 6.400 0.985 ;
        RECT 6.400 0.725 6.410 0.975 ;
        RECT 6.410 0.715 6.420 0.965 ;
        RECT 6.420 0.705 6.430 0.955 ;
        RECT 6.430 0.695 6.436 0.949 ;
        RECT 6.220 0.905 6.230 1.075 ;
        RECT 6.230 0.895 6.240 1.075 ;
        RECT 6.240 0.885 6.250 1.075 ;
        RECT 6.250 0.875 6.260 1.075 ;
        RECT 6.260 0.865 6.270 1.075 ;
        RECT 6.270 0.855 6.280 1.075 ;
        RECT 6.280 0.845 6.290 1.075 ;
        RECT 6.290 0.835 6.300 1.075 ;
        RECT 6.300 0.825 6.310 1.075 ;
        RECT 7.115 1.060 7.285 2.740 ;
        RECT 7.085 2.440 7.285 2.740 ;
        RECT 7.115 1.630 7.945 1.800 ;
        RECT 7.775 1.525 7.945 1.825 ;
  END 
END MUX4HD2XHT

MACRO MUX4HD1XHT
  CLASS  CORE ;
  FOREIGN MUX4HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.610 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.240 2.500 6.750 2.830 ;
    END
  END S1
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.175 1.890 4.420 2.440 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.485 1.730 2.830 2.140 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.060 0.910 2.470 1.450 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 1.110 1.140 1.665 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.665 ;
        RECT 2.375 -0.300 2.675 0.665 ;
        RECT 4.380 -0.300 4.680 0.680 ;
        RECT 5.930 -0.300 6.230 0.725 ;
        RECT 7.335 -0.300 7.850 0.780 ;
        RECT 0.000 -0.300 8.610 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.790 2.150 8.385 2.360 ;
        RECT 8.215 0.720 8.385 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.675 3.040 0.975 3.990 ;
        RECT 2.385 3.040 2.685 3.990 ;
        RECT 4.380 3.025 4.680 3.990 ;
        RECT 6.080 3.025 6.380 3.990 ;
        RECT 7.280 2.975 7.920 3.990 ;
        RECT 0.000 3.390 8.610 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.500 1.910 0.680 2.420 ;
        RECT 0.500 2.000 0.780 2.420 ;
        RECT 0.500 2.000 1.955 2.170 ;
        RECT 3.300 1.155 3.790 1.325 ;
        RECT 3.620 1.155 3.790 2.125 ;
        RECT 3.620 1.955 3.920 2.125 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.105 1.075 0.275 2.860 ;
        RECT 0.105 1.075 0.405 1.245 ;
        RECT 0.105 2.600 0.405 2.860 ;
        RECT 1.165 2.690 1.335 3.030 ;
        RECT 0.105 2.690 1.335 2.860 ;
        RECT 1.165 2.860 2.045 3.030 ;
        RECT 2.305 2.690 2.765 2.860 ;
        RECT 3.035 3.040 3.325 3.210 ;
        RECT 2.865 2.710 2.875 3.210 ;
        RECT 2.875 2.720 2.885 3.210 ;
        RECT 2.885 2.730 2.895 3.210 ;
        RECT 2.895 2.740 2.905 3.210 ;
        RECT 2.905 2.750 2.915 3.210 ;
        RECT 2.915 2.760 2.925 3.210 ;
        RECT 2.925 2.770 2.935 3.210 ;
        RECT 2.935 2.780 2.945 3.210 ;
        RECT 2.945 2.790 2.955 3.210 ;
        RECT 2.955 2.800 2.965 3.210 ;
        RECT 2.965 2.810 2.975 3.210 ;
        RECT 2.975 2.820 2.985 3.210 ;
        RECT 2.985 2.830 2.995 3.210 ;
        RECT 2.995 2.840 3.005 3.210 ;
        RECT 3.005 2.850 3.015 3.210 ;
        RECT 3.015 2.860 3.025 3.210 ;
        RECT 3.025 2.870 3.035 3.210 ;
        RECT 2.855 2.700 2.865 2.950 ;
        RECT 2.765 2.690 2.775 2.860 ;
        RECT 2.775 2.690 2.785 2.870 ;
        RECT 2.785 2.690 2.795 2.880 ;
        RECT 2.795 2.690 2.805 2.890 ;
        RECT 2.805 2.690 2.815 2.900 ;
        RECT 2.815 2.690 2.825 2.910 ;
        RECT 2.825 2.690 2.835 2.920 ;
        RECT 2.835 2.690 2.845 2.930 ;
        RECT 2.845 2.690 2.855 2.940 ;
        RECT 2.215 2.690 2.225 2.940 ;
        RECT 2.225 2.690 2.235 2.930 ;
        RECT 2.235 2.690 2.245 2.920 ;
        RECT 2.245 2.690 2.255 2.910 ;
        RECT 2.255 2.690 2.265 2.900 ;
        RECT 2.265 2.690 2.275 2.890 ;
        RECT 2.275 2.690 2.285 2.880 ;
        RECT 2.285 2.690 2.295 2.870 ;
        RECT 2.295 2.690 2.305 2.860 ;
        RECT 2.135 2.770 2.145 3.020 ;
        RECT 2.145 2.760 2.155 3.010 ;
        RECT 2.155 2.750 2.165 3.000 ;
        RECT 2.165 2.740 2.175 2.990 ;
        RECT 2.175 2.730 2.185 2.980 ;
        RECT 2.185 2.720 2.195 2.970 ;
        RECT 2.195 2.710 2.205 2.960 ;
        RECT 2.205 2.700 2.215 2.950 ;
        RECT 2.045 2.860 2.055 3.030 ;
        RECT 2.055 2.850 2.065 3.030 ;
        RECT 2.065 2.840 2.075 3.030 ;
        RECT 2.075 2.830 2.085 3.030 ;
        RECT 2.085 2.820 2.095 3.030 ;
        RECT 2.095 2.810 2.105 3.030 ;
        RECT 2.105 2.800 2.115 3.030 ;
        RECT 2.115 2.790 2.125 3.030 ;
        RECT 2.125 2.780 2.135 3.030 ;
        RECT 3.220 1.505 3.270 1.675 ;
        RECT 3.530 2.325 3.740 2.495 ;
        RECT 3.120 0.785 4.140 0.955 ;
        RECT 3.970 0.785 4.140 1.325 ;
        RECT 3.970 1.155 4.745 1.325 ;
        RECT 4.575 1.155 4.745 1.710 ;
        RECT 3.440 2.245 3.450 2.495 ;
        RECT 3.450 2.255 3.460 2.495 ;
        RECT 3.460 2.265 3.470 2.495 ;
        RECT 3.470 2.275 3.480 2.495 ;
        RECT 3.480 2.285 3.490 2.495 ;
        RECT 3.490 2.295 3.500 2.495 ;
        RECT 3.500 2.305 3.510 2.495 ;
        RECT 3.510 2.315 3.520 2.495 ;
        RECT 3.520 2.325 3.530 2.495 ;
        RECT 3.270 1.505 3.280 2.325 ;
        RECT 3.280 1.505 3.290 2.335 ;
        RECT 3.290 1.505 3.300 2.345 ;
        RECT 3.300 1.505 3.310 2.355 ;
        RECT 3.310 1.505 3.320 2.365 ;
        RECT 3.320 1.505 3.330 2.375 ;
        RECT 3.330 1.505 3.340 2.385 ;
        RECT 3.340 1.505 3.350 2.395 ;
        RECT 3.350 1.505 3.360 2.405 ;
        RECT 3.360 1.505 3.370 2.415 ;
        RECT 3.370 1.505 3.380 2.425 ;
        RECT 3.380 1.505 3.390 2.435 ;
        RECT 3.390 1.505 3.400 2.445 ;
        RECT 3.400 1.505 3.410 2.455 ;
        RECT 3.410 1.505 3.420 2.465 ;
        RECT 3.420 1.505 3.430 2.475 ;
        RECT 3.430 1.505 3.440 2.485 ;
        RECT 3.130 1.425 3.140 1.675 ;
        RECT 3.140 1.435 3.150 1.675 ;
        RECT 3.150 1.445 3.160 1.675 ;
        RECT 3.160 1.455 3.170 1.675 ;
        RECT 3.170 1.465 3.180 1.675 ;
        RECT 3.180 1.475 3.190 1.675 ;
        RECT 3.190 1.485 3.200 1.675 ;
        RECT 3.200 1.495 3.210 1.675 ;
        RECT 3.210 1.505 3.220 1.675 ;
        RECT 3.120 1.415 3.130 1.665 ;
        RECT 2.950 0.785 2.960 1.495 ;
        RECT 2.960 0.785 2.970 1.505 ;
        RECT 2.970 0.785 2.980 1.515 ;
        RECT 2.980 0.785 2.990 1.525 ;
        RECT 2.990 0.785 3.000 1.535 ;
        RECT 3.000 0.785 3.010 1.545 ;
        RECT 3.010 0.785 3.020 1.555 ;
        RECT 3.020 0.785 3.030 1.565 ;
        RECT 3.030 0.785 3.040 1.575 ;
        RECT 3.040 0.785 3.050 1.585 ;
        RECT 3.050 0.785 3.060 1.595 ;
        RECT 3.060 0.785 3.070 1.605 ;
        RECT 3.070 0.785 3.080 1.615 ;
        RECT 3.080 0.785 3.090 1.625 ;
        RECT 3.090 0.785 3.100 1.635 ;
        RECT 3.100 0.785 3.110 1.645 ;
        RECT 3.110 0.785 3.120 1.655 ;
        RECT 1.520 0.720 1.690 1.820 ;
        RECT 1.515 2.370 2.015 2.540 ;
        RECT 2.045 2.340 2.105 2.540 ;
        RECT 1.520 1.650 2.305 1.820 ;
        RECT 2.135 1.650 2.305 2.510 ;
        RECT 2.135 2.340 2.935 2.510 ;
        RECT 3.360 2.675 3.595 2.855 ;
        RECT 3.360 2.675 5.800 2.845 ;
        RECT 6.105 1.610 6.165 2.190 ;
        RECT 5.995 1.610 6.005 2.290 ;
        RECT 6.005 1.610 6.015 2.280 ;
        RECT 6.015 1.610 6.025 2.270 ;
        RECT 6.025 1.610 6.035 2.260 ;
        RECT 6.035 1.610 6.045 2.250 ;
        RECT 6.045 1.610 6.055 2.240 ;
        RECT 6.055 1.610 6.065 2.230 ;
        RECT 6.065 1.610 6.075 2.220 ;
        RECT 6.075 1.610 6.085 2.210 ;
        RECT 6.085 1.610 6.095 2.200 ;
        RECT 6.095 1.610 6.105 2.190 ;
        RECT 5.970 2.065 5.980 2.835 ;
        RECT 5.980 2.055 5.990 2.825 ;
        RECT 5.990 2.045 5.996 2.819 ;
        RECT 5.825 2.210 5.835 2.844 ;
        RECT 5.835 2.200 5.845 2.844 ;
        RECT 5.845 2.190 5.855 2.844 ;
        RECT 5.855 2.180 5.865 2.844 ;
        RECT 5.865 2.170 5.875 2.844 ;
        RECT 5.875 2.160 5.885 2.844 ;
        RECT 5.885 2.150 5.895 2.844 ;
        RECT 5.895 2.140 5.905 2.844 ;
        RECT 5.905 2.130 5.915 2.844 ;
        RECT 5.915 2.120 5.925 2.844 ;
        RECT 5.925 2.110 5.935 2.844 ;
        RECT 5.935 2.100 5.945 2.844 ;
        RECT 5.945 2.090 5.955 2.844 ;
        RECT 5.955 2.080 5.965 2.844 ;
        RECT 5.965 2.070 5.971 2.844 ;
        RECT 5.800 2.675 5.810 2.845 ;
        RECT 5.810 2.665 5.820 2.845 ;
        RECT 5.820 2.655 5.826 2.845 ;
        RECT 3.280 2.605 3.290 2.855 ;
        RECT 3.290 2.615 3.300 2.855 ;
        RECT 3.300 2.625 3.310 2.855 ;
        RECT 3.310 2.635 3.320 2.855 ;
        RECT 3.320 2.645 3.330 2.855 ;
        RECT 3.330 2.655 3.340 2.855 ;
        RECT 3.340 2.665 3.350 2.855 ;
        RECT 3.350 2.675 3.360 2.855 ;
        RECT 3.025 2.350 3.035 2.600 ;
        RECT 3.035 2.360 3.045 2.610 ;
        RECT 3.045 2.370 3.055 2.620 ;
        RECT 3.055 2.380 3.065 2.630 ;
        RECT 3.065 2.390 3.075 2.640 ;
        RECT 3.075 2.400 3.085 2.650 ;
        RECT 3.085 2.410 3.095 2.660 ;
        RECT 3.095 2.420 3.105 2.670 ;
        RECT 3.105 2.430 3.115 2.680 ;
        RECT 3.115 2.440 3.125 2.690 ;
        RECT 3.125 2.450 3.135 2.700 ;
        RECT 3.135 2.460 3.145 2.710 ;
        RECT 3.145 2.470 3.155 2.720 ;
        RECT 3.155 2.480 3.165 2.730 ;
        RECT 3.165 2.490 3.175 2.740 ;
        RECT 3.175 2.500 3.185 2.750 ;
        RECT 3.185 2.510 3.195 2.760 ;
        RECT 3.195 2.520 3.205 2.770 ;
        RECT 3.205 2.530 3.215 2.780 ;
        RECT 3.215 2.540 3.225 2.790 ;
        RECT 3.225 2.550 3.235 2.800 ;
        RECT 3.235 2.560 3.245 2.810 ;
        RECT 3.245 2.570 3.255 2.820 ;
        RECT 3.255 2.580 3.265 2.830 ;
        RECT 3.265 2.590 3.275 2.840 ;
        RECT 3.275 2.595 3.281 2.849 ;
        RECT 2.935 2.340 2.945 2.510 ;
        RECT 2.945 2.340 2.955 2.520 ;
        RECT 2.955 2.340 2.965 2.530 ;
        RECT 2.965 2.340 2.975 2.540 ;
        RECT 2.975 2.340 2.985 2.550 ;
        RECT 2.985 2.340 2.995 2.560 ;
        RECT 2.995 2.340 3.005 2.570 ;
        RECT 3.005 2.340 3.015 2.580 ;
        RECT 3.015 2.340 3.025 2.590 ;
        RECT 2.105 2.340 2.115 2.530 ;
        RECT 2.115 2.340 2.125 2.520 ;
        RECT 2.125 2.340 2.135 2.510 ;
        RECT 2.015 2.370 2.025 2.540 ;
        RECT 2.025 2.360 2.035 2.540 ;
        RECT 2.035 2.350 2.045 2.540 ;
        RECT 5.630 1.805 5.700 1.995 ;
        RECT 5.620 1.815 5.806 1.889 ;
        RECT 5.400 1.825 5.700 1.995 ;
        RECT 5.400 1.825 5.710 1.985 ;
        RECT 5.400 1.825 5.720 1.975 ;
        RECT 5.400 1.825 5.730 1.965 ;
        RECT 5.400 1.825 5.740 1.955 ;
        RECT 5.400 1.825 5.750 1.945 ;
        RECT 5.400 1.825 5.760 1.935 ;
        RECT 5.400 1.825 5.770 1.925 ;
        RECT 5.400 1.825 5.780 1.915 ;
        RECT 5.400 1.825 5.790 1.905 ;
        RECT 5.400 1.825 5.800 1.895 ;
        RECT 5.635 1.255 5.806 1.889 ;
        RECT 6.630 1.105 6.865 1.425 ;
        RECT 5.635 1.255 6.865 1.425 ;
        RECT 6.695 1.105 6.865 2.280 ;
        RECT 6.630 1.105 6.930 1.275 ;
        RECT 4.965 1.170 5.135 2.495 ;
        RECT 5.285 0.905 5.455 1.340 ;
        RECT 4.965 1.170 5.455 1.340 ;
        RECT 4.965 2.325 5.520 2.495 ;
        RECT 5.285 0.905 6.310 1.075 ;
        RECT 6.570 0.735 7.155 0.905 ;
        RECT 6.480 0.735 6.490 0.985 ;
        RECT 6.490 0.735 6.500 0.975 ;
        RECT 6.500 0.735 6.510 0.965 ;
        RECT 6.510 0.735 6.520 0.955 ;
        RECT 6.520 0.735 6.530 0.945 ;
        RECT 6.530 0.735 6.540 0.935 ;
        RECT 6.540 0.735 6.550 0.925 ;
        RECT 6.550 0.735 6.560 0.915 ;
        RECT 6.560 0.735 6.570 0.905 ;
        RECT 6.400 0.815 6.410 1.065 ;
        RECT 6.410 0.805 6.420 1.055 ;
        RECT 6.420 0.795 6.430 1.045 ;
        RECT 6.430 0.785 6.440 1.035 ;
        RECT 6.440 0.775 6.450 1.025 ;
        RECT 6.450 0.765 6.460 1.015 ;
        RECT 6.460 0.755 6.470 1.005 ;
        RECT 6.470 0.745 6.480 0.995 ;
        RECT 6.310 0.905 6.320 1.075 ;
        RECT 6.320 0.895 6.330 1.075 ;
        RECT 6.330 0.885 6.340 1.075 ;
        RECT 6.340 0.875 6.350 1.075 ;
        RECT 6.350 0.865 6.360 1.075 ;
        RECT 6.360 0.855 6.370 1.075 ;
        RECT 6.370 0.845 6.380 1.075 ;
        RECT 6.380 0.835 6.390 1.075 ;
        RECT 6.390 0.825 6.400 1.075 ;
        RECT 7.205 1.125 7.375 2.280 ;
        RECT 7.140 1.125 7.440 1.295 ;
        RECT 7.205 1.590 8.035 1.760 ;
        RECT 7.865 1.525 8.035 1.825 ;
  END 
END MUX4HD1XHT

MACRO MUX2HDUXHT
  CLASS  CORE ;
  FOREIGN MUX2HDUXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.090 2.500 0.385 3.020 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.095 1.160 2.505 1.665 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.660 ;
        RECT 2.345 -0.300 2.645 0.660 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.875 0.655 3.190 0.825 ;
        RECT 2.995 0.655 3.190 3.025 ;
        RECT 2.875 2.390 3.190 3.025 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 2.575 0.865 3.990 ;
        RECT 2.345 2.790 2.645 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.520 1.505 1.555 1.970 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.170 0.840 0.340 2.320 ;
        RECT 0.170 2.150 1.215 2.320 ;
        RECT 1.045 2.150 1.215 2.910 ;
        RECT 1.125 0.500 1.305 1.020 ;
        RECT 0.170 0.840 1.305 1.020 ;
        RECT 1.045 2.740 2.025 2.910 ;
        RECT 1.515 1.125 1.915 1.295 ;
        RECT 1.745 1.125 1.915 2.495 ;
        RECT 1.515 2.325 1.915 2.495 ;
        RECT 1.745 1.890 2.810 2.190 ;
  END 
END MUX2HDUXHT

MACRO MUX2HDMXHT
  CLASS  CORE ;
  FOREIGN MUX2HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.705 1.570 1.200 1.950 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.950 2.485 2.465 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 2.315 -0.300 2.615 0.725 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.930 1.060 3.180 1.360 ;
        RECT 2.970 1.060 3.180 2.540 ;
        RECT 2.865 2.370 3.180 2.540 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.490 0.925 3.990 ;
        RECT 2.315 3.040 2.615 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.200 2.860 1.775 3.180 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.605 ;
        RECT 1.400 1.560 1.570 2.305 ;
        RECT 0.170 2.135 1.570 2.305 ;
        RECT 1.515 1.125 1.920 1.295 ;
        RECT 1.750 1.125 1.920 2.660 ;
        RECT 1.515 2.490 1.920 2.660 ;
        RECT 1.750 1.465 2.780 1.635 ;
        RECT 2.610 1.465 2.780 1.765 ;
  END 
END MUX2HDMXHT

MACRO MUX2HDLXHT
  CLASS  CORE ;
  FOREIGN MUX2HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.800 1.570 1.200 1.950 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.990 2.565 2.425 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 2.445 -0.300 2.745 0.745 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.875 1.125 3.180 1.295 ;
        RECT 2.970 1.125 3.180 2.540 ;
        RECT 2.875 2.370 3.180 2.540 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.490 0.925 3.990 ;
        RECT 2.445 3.095 2.745 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.200 2.860 1.775 3.180 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.605 ;
        RECT 0.170 2.130 0.345 2.605 ;
        RECT 1.400 1.560 1.570 2.300 ;
        RECT 0.170 2.130 1.570 2.300 ;
        RECT 1.515 1.125 1.920 1.295 ;
        RECT 1.750 1.125 1.920 2.660 ;
        RECT 1.515 2.490 1.920 2.660 ;
        RECT 1.750 1.460 2.790 1.630 ;
        RECT 2.620 1.460 2.790 1.760 ;
  END 
END MUX2HDLXHT

MACRO MUX2HD3XHT
  CLASS  CORE ;
  FOREIGN MUX2HD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.900 1.395 1.155 2.105 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.725 1.640 3.180 2.020 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.715 ;
        RECT 3.005 -0.300 3.305 1.055 ;
        RECT 4.140 -0.300 4.315 1.120 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.555 0.505 3.940 1.080 ;
        RECT 3.730 2.220 3.900 3.045 ;
        RECT 3.620 2.405 3.900 3.045 ;
        RECT 3.720 0.505 3.940 1.495 ;
        RECT 3.720 1.325 4.895 1.495 ;
        RECT 4.195 1.325 4.895 2.390 ;
        RECT 3.730 2.220 4.895 2.390 ;
        RECT 4.595 0.720 4.895 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.635 0.955 3.990 ;
        RECT 3.035 2.635 3.335 3.990 ;
        RECT 4.140 2.570 4.375 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.550 1.045 0.720 1.800 ;
        RECT 0.440 1.260 0.720 1.800 ;
        RECT 0.550 1.045 2.005 1.215 ;
        RECT 1.825 1.045 2.005 1.665 ;
        RECT 1.825 1.495 2.125 1.665 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.090 0.710 0.260 2.455 ;
        RECT 0.090 0.710 0.405 0.880 ;
        RECT 0.090 1.990 0.405 2.455 ;
        RECT 1.400 1.430 1.570 2.455 ;
        RECT 0.090 2.285 1.570 2.455 ;
        RECT 2.370 1.610 2.540 2.015 ;
        RECT 1.400 1.845 2.540 2.015 ;
        RECT 2.060 2.230 2.230 3.210 ;
        RECT 1.645 0.655 2.575 0.825 ;
        RECT 2.405 0.655 2.575 1.430 ;
        RECT 2.060 2.230 3.225 2.400 ;
        RECT 2.405 1.260 3.360 1.430 ;
        RECT 3.530 1.675 4.015 1.845 ;
        RECT 3.360 1.260 3.370 2.330 ;
        RECT 3.370 1.260 3.380 2.320 ;
        RECT 3.380 1.260 3.390 2.310 ;
        RECT 3.390 1.260 3.400 2.300 ;
        RECT 3.400 1.260 3.410 2.290 ;
        RECT 3.410 1.260 3.420 2.280 ;
        RECT 3.420 1.260 3.430 2.270 ;
        RECT 3.430 1.260 3.440 2.260 ;
        RECT 3.440 1.260 3.450 2.250 ;
        RECT 3.450 1.260 3.460 2.240 ;
        RECT 3.460 1.260 3.470 2.230 ;
        RECT 3.470 1.260 3.480 2.220 ;
        RECT 3.480 1.260 3.490 2.210 ;
        RECT 3.490 1.260 3.500 2.200 ;
        RECT 3.500 1.260 3.510 2.190 ;
        RECT 3.510 1.260 3.520 2.180 ;
        RECT 3.520 1.260 3.530 2.170 ;
        RECT 3.300 2.155 3.310 2.389 ;
        RECT 3.310 2.145 3.320 2.379 ;
        RECT 3.320 2.135 3.330 2.369 ;
        RECT 3.330 2.125 3.340 2.359 ;
        RECT 3.340 2.115 3.350 2.349 ;
        RECT 3.350 2.105 3.360 2.339 ;
        RECT 3.225 2.230 3.235 2.400 ;
        RECT 3.235 2.220 3.245 2.400 ;
        RECT 3.245 2.210 3.255 2.400 ;
        RECT 3.255 2.200 3.265 2.400 ;
        RECT 3.265 2.190 3.275 2.400 ;
        RECT 3.275 2.180 3.285 2.400 ;
        RECT 3.285 2.170 3.295 2.400 ;
        RECT 3.295 2.160 3.301 2.400 ;
  END 
END MUX2HD3XHT

MACRO MUX2HD1XHT
  CLASS  CORE ;
  FOREIGN MUX2HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.570 1.250 2.010 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.310 1.845 2.480 2.360 ;
        RECT 2.310 2.150 2.885 2.360 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.695 -0.300 0.995 1.295 ;
        RECT 2.595 -0.300 2.895 1.055 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.180 0.720 3.390 1.360 ;
        RECT 3.220 0.720 3.390 2.960 ;
        RECT 3.180 1.980 3.390 2.960 ;
        RECT 3.220 1.670 3.590 2.015 ;
        RECT 3.180 1.980 3.590 2.015 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.695 2.545 0.995 3.990 ;
        RECT 2.595 2.635 2.895 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.475 0.740 2.010 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.160 1.125 0.330 2.595 ;
        RECT 0.160 1.125 0.475 1.295 ;
        RECT 0.160 2.190 0.475 2.595 ;
        RECT 1.470 1.560 1.640 2.360 ;
        RECT 0.160 2.190 1.640 2.360 ;
        RECT 1.585 1.125 1.990 1.295 ;
        RECT 1.820 1.125 1.990 2.715 ;
        RECT 1.585 2.545 1.990 2.715 ;
        RECT 1.820 1.475 3.030 1.645 ;
        RECT 2.860 1.475 3.030 1.870 ;
  END 
END MUX2HD1XHT

MACRO LATNSRHDMXHT
  CLASS  CORE ;
  FOREIGN LATNSRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.430 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.005 1.125 7.305 1.295 ;
        RECT 7.105 1.125 7.305 2.890 ;
        RECT 7.030 2.460 7.305 2.890 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.565 0.965 2.055 ;
        RECT 0.510 1.565 1.000 1.865 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.090 1.060 9.330 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.970 1.255 3.185 1.840 ;
        RECT 2.970 1.540 3.370 1.840 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.980 0.480 5.610 1.215 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 2.265 -0.300 2.565 0.595 ;
        RECT 5.790 -0.300 5.960 1.085 ;
        RECT 7.700 -0.300 8.005 0.745 ;
        RECT 8.505 -0.300 8.805 1.145 ;
        RECT 0.000 -0.300 9.430 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.355 2.745 2.065 3.180 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.905 0.895 3.990 ;
        RECT 2.270 2.745 2.440 3.990 ;
        RECT 5.695 2.545 5.865 3.990 ;
        RECT 7.490 2.220 7.790 3.990 ;
        RECT 8.475 2.560 8.775 3.990 ;
        RECT 0.000 3.390 9.430 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.655 1.125 1.955 1.295 ;
        RECT 1.785 1.125 1.955 2.215 ;
        RECT 1.655 2.045 1.955 2.215 ;
        RECT 1.785 1.675 2.615 1.845 ;
        RECT 3.420 1.125 3.720 1.295 ;
        RECT 3.550 1.125 3.720 2.370 ;
        RECT 3.240 2.200 3.720 2.370 ;
        RECT 1.210 0.625 1.445 1.360 ;
        RECT 1.275 0.625 1.445 2.215 ;
        RECT 1.145 2.045 1.445 2.215 ;
        RECT 1.210 0.625 1.585 0.945 ;
        RECT 2.975 0.605 3.145 0.945 ;
        RECT 1.210 0.775 3.145 0.945 ;
        RECT 2.975 0.605 4.045 0.775 ;
        RECT 0.105 1.125 0.275 2.565 ;
        RECT 0.105 1.125 0.405 1.295 ;
        RECT 0.105 2.345 0.405 2.565 ;
        RECT 2.880 2.395 3.060 2.720 ;
        RECT 0.105 2.395 3.060 2.565 ;
        RECT 2.880 2.550 4.050 2.720 ;
        RECT 3.925 1.030 4.050 2.860 ;
        RECT 4.095 2.690 4.340 2.860 ;
        RECT 4.630 0.705 4.800 1.020 ;
        RECT 4.340 0.820 4.800 1.020 ;
        RECT 4.260 0.820 4.270 1.090 ;
        RECT 4.270 0.820 4.280 1.080 ;
        RECT 4.280 0.820 4.290 1.070 ;
        RECT 4.290 0.820 4.300 1.060 ;
        RECT 4.300 0.820 4.310 1.050 ;
        RECT 4.310 0.820 4.320 1.040 ;
        RECT 4.320 0.820 4.330 1.030 ;
        RECT 4.330 0.820 4.340 1.020 ;
        RECT 4.160 0.920 4.170 1.190 ;
        RECT 4.170 0.910 4.180 1.180 ;
        RECT 4.180 0.900 4.190 1.170 ;
        RECT 4.190 0.890 4.200 1.160 ;
        RECT 4.200 0.880 4.210 1.150 ;
        RECT 4.210 0.870 4.220 1.140 ;
        RECT 4.220 0.860 4.230 1.130 ;
        RECT 4.230 0.850 4.240 1.120 ;
        RECT 4.240 0.840 4.250 1.110 ;
        RECT 4.250 0.830 4.260 1.100 ;
        RECT 4.095 0.985 4.105 1.199 ;
        RECT 4.105 0.975 4.115 1.199 ;
        RECT 4.115 0.965 4.125 1.199 ;
        RECT 4.125 0.955 4.135 1.199 ;
        RECT 4.135 0.945 4.145 1.199 ;
        RECT 4.145 0.935 4.155 1.199 ;
        RECT 4.155 0.925 4.161 1.199 ;
        RECT 4.050 1.030 4.060 2.860 ;
        RECT 4.060 1.020 4.070 2.860 ;
        RECT 4.070 1.010 4.080 2.860 ;
        RECT 4.080 1.000 4.090 2.860 ;
        RECT 4.090 0.990 4.096 2.860 ;
        RECT 2.640 2.890 2.810 3.190 ;
        RECT 2.640 2.900 3.635 3.070 ;
        RECT 4.520 2.900 4.690 3.210 ;
        RECT 3.850 3.040 4.690 3.210 ;
        RECT 4.520 2.900 5.515 3.070 ;
        RECT 5.215 2.900 5.515 3.210 ;
        RECT 3.775 2.975 3.785 3.209 ;
        RECT 3.785 2.985 3.795 3.209 ;
        RECT 3.795 2.995 3.805 3.209 ;
        RECT 3.805 3.005 3.815 3.209 ;
        RECT 3.815 3.015 3.825 3.209 ;
        RECT 3.825 3.025 3.835 3.209 ;
        RECT 3.835 3.035 3.845 3.209 ;
        RECT 3.845 3.040 3.851 3.210 ;
        RECT 3.710 2.910 3.720 3.144 ;
        RECT 3.720 2.920 3.730 3.154 ;
        RECT 3.730 2.930 3.740 3.164 ;
        RECT 3.740 2.940 3.750 3.174 ;
        RECT 3.750 2.950 3.760 3.184 ;
        RECT 3.760 2.960 3.770 3.194 ;
        RECT 3.770 2.965 3.776 3.205 ;
        RECT 3.635 2.900 3.645 3.070 ;
        RECT 3.645 2.900 3.655 3.080 ;
        RECT 3.655 2.900 3.665 3.090 ;
        RECT 3.665 2.900 3.675 3.100 ;
        RECT 3.675 2.900 3.685 3.110 ;
        RECT 3.685 2.900 3.695 3.120 ;
        RECT 3.695 2.900 3.705 3.130 ;
        RECT 3.705 2.900 3.711 3.140 ;
        RECT 4.340 1.275 4.645 1.445 ;
        RECT 4.280 2.200 4.580 2.370 ;
        RECT 4.475 1.275 4.645 2.365 ;
        RECT 6.490 1.060 6.815 1.360 ;
        RECT 6.615 2.005 6.815 2.365 ;
        RECT 4.475 2.175 6.815 2.365 ;
        RECT 6.645 1.060 6.815 2.365 ;
        RECT 6.645 1.565 6.925 1.865 ;
        RECT 6.140 0.710 6.310 1.930 ;
        RECT 4.970 1.760 6.310 1.930 ;
        RECT 6.140 0.710 7.320 0.880 ;
        RECT 7.655 0.960 8.230 1.130 ;
        RECT 8.060 0.960 8.230 2.335 ;
        RECT 8.060 2.035 8.250 2.335 ;
        RECT 8.060 1.480 8.910 1.780 ;
        RECT 7.570 0.885 7.580 1.129 ;
        RECT 7.580 0.895 7.590 1.129 ;
        RECT 7.590 0.905 7.600 1.129 ;
        RECT 7.600 0.915 7.610 1.129 ;
        RECT 7.610 0.925 7.620 1.129 ;
        RECT 7.620 0.935 7.630 1.129 ;
        RECT 7.630 0.945 7.640 1.129 ;
        RECT 7.640 0.955 7.650 1.129 ;
        RECT 7.650 0.960 7.656 1.130 ;
        RECT 7.405 0.720 7.415 0.964 ;
        RECT 7.415 0.730 7.425 0.974 ;
        RECT 7.425 0.740 7.435 0.984 ;
        RECT 7.435 0.750 7.445 0.994 ;
        RECT 7.445 0.760 7.455 1.004 ;
        RECT 7.455 0.770 7.465 1.014 ;
        RECT 7.465 0.780 7.475 1.024 ;
        RECT 7.475 0.790 7.485 1.034 ;
        RECT 7.485 0.800 7.495 1.044 ;
        RECT 7.495 0.810 7.505 1.054 ;
        RECT 7.505 0.820 7.515 1.064 ;
        RECT 7.515 0.830 7.525 1.074 ;
        RECT 7.525 0.840 7.535 1.084 ;
        RECT 7.535 0.850 7.545 1.094 ;
        RECT 7.545 0.860 7.555 1.104 ;
        RECT 7.555 0.870 7.565 1.114 ;
        RECT 7.565 0.875 7.571 1.125 ;
        RECT 7.320 0.710 7.330 0.880 ;
        RECT 7.330 0.710 7.340 0.890 ;
        RECT 7.340 0.710 7.350 0.900 ;
        RECT 7.350 0.710 7.360 0.910 ;
        RECT 7.360 0.710 7.370 0.920 ;
        RECT 7.370 0.710 7.380 0.930 ;
        RECT 7.380 0.710 7.390 0.940 ;
        RECT 7.390 0.710 7.400 0.950 ;
        RECT 7.400 0.710 7.406 0.960 ;
  END 
END LATNSRHDMXHT

MACRO LATNSRHDLXHT
  CLASS  CORE ;
  FOREIGN LATNSRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.020 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 6.660 1.580 7.065 1.750 ;
        RECT 6.895 1.125 6.985 2.280 ;
        RECT 6.660 1.125 6.985 1.750 ;
        RECT 6.895 1.580 7.065 2.280 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.565 0.965 2.030 ;
        RECT 0.510 1.565 1.095 1.865 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.615 1.125 8.920 1.295 ;
        RECT 8.750 1.125 8.920 2.910 ;
        RECT 8.515 2.485 8.920 2.910 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.885 1.235 3.180 1.950 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.770 0.480 5.360 0.720 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.685 -0.300 0.985 1.295 ;
        RECT 2.225 -0.300 2.525 0.595 ;
        RECT 5.540 -0.300 5.710 1.360 ;
        RECT 7.570 -0.300 8.080 0.810 ;
        RECT 0.000 -0.300 9.020 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.355 2.855 2.090 3.180 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.855 0.895 3.990 ;
        RECT 2.270 2.855 2.440 3.990 ;
        RECT 5.400 2.420 5.700 3.990 ;
        RECT 7.415 2.100 7.585 3.990 ;
        RECT 7.995 2.730 8.165 3.990 ;
        RECT 0.000 3.390 9.020 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.775 1.125 2.075 1.295 ;
        RECT 1.905 1.125 2.075 2.325 ;
        RECT 1.655 2.155 2.075 2.325 ;
        RECT 1.905 1.720 2.650 2.020 ;
        RECT 3.360 1.060 3.530 2.390 ;
        RECT 1.275 0.625 1.445 2.215 ;
        RECT 1.145 2.045 1.445 2.215 ;
        RECT 1.275 0.625 1.500 1.360 ;
        RECT 1.275 0.625 1.655 0.945 ;
        RECT 2.975 0.605 3.145 0.945 ;
        RECT 1.275 0.775 3.145 0.945 ;
        RECT 2.975 0.605 3.675 0.775 ;
        RECT 0.105 1.125 0.275 2.675 ;
        RECT 0.105 1.125 0.405 1.295 ;
        RECT 0.105 2.185 0.405 2.675 ;
        RECT 3.005 2.505 3.175 2.740 ;
        RECT 0.105 2.505 3.175 2.675 ;
        RECT 3.005 2.570 3.710 2.740 ;
        RECT 3.635 2.570 3.710 2.840 ;
        RECT 3.880 2.570 3.935 2.840 ;
        RECT 4.265 0.605 4.580 0.955 ;
        RECT 4.020 0.755 4.580 0.955 ;
        RECT 3.955 0.755 3.965 1.009 ;
        RECT 3.965 0.755 3.975 0.999 ;
        RECT 3.975 0.755 3.985 0.989 ;
        RECT 3.985 0.755 3.995 0.979 ;
        RECT 3.995 0.755 4.005 0.969 ;
        RECT 4.005 0.755 4.015 0.959 ;
        RECT 4.015 0.755 4.021 0.955 ;
        RECT 3.880 0.830 3.890 1.084 ;
        RECT 3.890 0.820 3.900 1.074 ;
        RECT 3.900 0.810 3.910 1.064 ;
        RECT 3.910 0.800 3.920 1.054 ;
        RECT 3.920 0.790 3.930 1.044 ;
        RECT 3.930 0.780 3.940 1.034 ;
        RECT 3.940 0.770 3.950 1.024 ;
        RECT 3.950 0.760 3.956 1.020 ;
        RECT 3.710 1.000 3.720 2.840 ;
        RECT 3.720 0.990 3.730 2.840 ;
        RECT 3.730 0.980 3.740 2.840 ;
        RECT 3.740 0.970 3.750 2.840 ;
        RECT 3.750 0.960 3.760 2.840 ;
        RECT 3.760 0.950 3.770 2.840 ;
        RECT 3.770 0.940 3.780 2.840 ;
        RECT 3.780 0.930 3.790 2.840 ;
        RECT 3.790 0.920 3.800 2.840 ;
        RECT 3.800 0.910 3.810 2.840 ;
        RECT 3.810 0.900 3.820 2.840 ;
        RECT 3.820 0.890 3.830 2.840 ;
        RECT 3.830 0.880 3.840 2.840 ;
        RECT 3.840 0.870 3.850 2.840 ;
        RECT 3.850 0.860 3.860 2.840 ;
        RECT 3.860 0.850 3.870 2.840 ;
        RECT 3.870 0.840 3.880 2.840 ;
        RECT 2.640 2.890 2.810 3.190 ;
        RECT 3.285 2.920 3.455 3.190 ;
        RECT 2.640 2.920 3.455 3.090 ;
        RECT 4.115 2.855 4.285 3.190 ;
        RECT 3.285 3.020 4.285 3.190 ;
        RECT 4.115 2.855 5.220 3.025 ;
        RECT 5.050 2.855 5.220 3.155 ;
        RECT 4.115 2.090 4.285 2.390 ;
        RECT 4.135 1.135 4.305 2.240 ;
        RECT 6.240 1.060 6.480 1.360 ;
        RECT 4.135 2.060 6.555 2.240 ;
        RECT 6.285 1.060 6.480 2.240 ;
        RECT 6.385 2.060 6.555 2.815 ;
        RECT 6.385 2.515 7.235 2.815 ;
        RECT 5.890 0.710 6.060 1.845 ;
        RECT 4.710 1.675 6.060 1.845 ;
        RECT 5.890 0.710 7.335 0.880 ;
        RECT 7.165 0.710 7.335 1.295 ;
        RECT 7.165 1.125 8.075 1.295 ;
        RECT 7.905 1.125 8.075 2.280 ;
        RECT 7.905 1.980 8.505 2.280 ;
  END 
END LATNSRHDLXHT

MACRO LATNSRHD2XHT
  CLASS  CORE ;
  FOREIGN LATNSRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.070 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.045 1.125 8.345 1.295 ;
        RECT 8.175 1.125 8.345 2.895 ;
        RECT 8.175 1.740 8.360 2.895 ;
        RECT 7.955 2.045 8.360 2.895 ;
        RECT 8.175 1.740 8.580 1.950 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.565 0.965 2.055 ;
        RECT 0.510 1.565 1.000 1.865 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.210 2.085 10.380 3.065 ;
        RECT 10.145 0.785 10.445 1.295 ;
        RECT 10.145 1.125 10.890 1.295 ;
        RECT 10.720 1.125 10.890 2.360 ;
        RECT 10.210 2.085 10.890 2.360 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.310 1.330 3.655 1.910 ;
        RECT 3.310 1.610 3.795 1.910 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.620 0.500 2.920 0.700 ;
        RECT 2.620 0.530 5.715 0.700 ;
        RECT 5.350 0.500 5.715 0.720 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 2.270 -0.300 2.440 0.660 ;
        RECT 6.255 -0.300 6.555 0.980 ;
        RECT 7.495 -0.300 7.795 0.595 ;
        RECT 8.595 -0.300 8.895 0.595 ;
        RECT 9.625 -0.300 9.925 0.715 ;
        RECT 10.665 -0.300 10.965 0.715 ;
        RECT 0.000 -0.300 11.070 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.355 2.745 2.035 3.180 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.895 0.895 3.990 ;
        RECT 2.270 2.910 2.440 3.990 ;
        RECT 6.090 2.540 6.395 3.990 ;
        RECT 7.435 2.635 7.735 3.990 ;
        RECT 8.540 2.230 8.710 3.990 ;
        RECT 9.625 2.295 9.925 3.990 ;
        RECT 10.665 2.635 10.965 3.990 ;
        RECT 0.000 3.390 11.070 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 0.275 2.565 ;
        RECT 0.105 1.125 0.405 1.295 ;
        RECT 0.105 2.345 0.405 2.565 ;
        RECT 0.105 2.395 2.790 2.565 ;
        RECT 2.620 2.395 2.790 3.075 ;
        RECT 2.620 2.905 3.795 3.075 ;
        RECT 3.495 2.905 3.795 3.190 ;
        RECT 3.845 1.230 4.145 1.400 ;
        RECT 3.975 1.230 4.145 2.320 ;
        RECT 3.320 2.150 4.145 2.320 ;
        RECT 1.210 0.625 1.445 1.360 ;
        RECT 1.275 0.625 1.445 2.215 ;
        RECT 1.145 2.045 1.445 2.215 ;
        RECT 1.210 0.625 1.585 0.945 ;
        RECT 1.210 0.775 2.035 0.945 ;
        RECT 2.230 0.880 4.495 1.050 ;
        RECT 4.325 0.880 4.495 2.720 ;
        RECT 4.325 2.550 5.085 2.720 ;
        RECT 4.785 2.550 5.085 2.840 ;
        RECT 2.140 0.800 2.150 1.050 ;
        RECT 2.150 0.810 2.160 1.050 ;
        RECT 2.160 0.820 2.170 1.050 ;
        RECT 2.170 0.830 2.180 1.050 ;
        RECT 2.180 0.840 2.190 1.050 ;
        RECT 2.190 0.850 2.200 1.050 ;
        RECT 2.200 0.860 2.210 1.050 ;
        RECT 2.210 0.870 2.220 1.050 ;
        RECT 2.220 0.880 2.230 1.050 ;
        RECT 2.125 0.785 2.135 1.035 ;
        RECT 2.135 0.790 2.141 1.044 ;
        RECT 2.035 0.775 2.045 0.945 ;
        RECT 2.045 0.775 2.055 0.955 ;
        RECT 2.055 0.775 2.065 0.965 ;
        RECT 2.065 0.775 2.075 0.975 ;
        RECT 2.075 0.775 2.085 0.985 ;
        RECT 2.085 0.775 2.095 0.995 ;
        RECT 2.095 0.775 2.105 1.005 ;
        RECT 2.105 0.775 2.115 1.015 ;
        RECT 2.115 0.775 2.125 1.025 ;
        RECT 1.655 1.125 1.955 1.295 ;
        RECT 1.785 1.125 1.955 2.215 ;
        RECT 2.450 1.610 2.620 2.215 ;
        RECT 1.655 2.045 3.140 2.215 ;
        RECT 2.970 2.045 3.140 2.725 ;
        RECT 2.970 2.555 4.145 2.725 ;
        RECT 3.975 2.555 4.145 3.085 ;
        RECT 4.535 3.020 5.565 3.095 ;
        RECT 4.545 3.020 5.565 3.105 ;
        RECT 4.555 3.020 5.565 3.115 ;
        RECT 4.565 3.020 5.565 3.125 ;
        RECT 4.575 3.020 5.565 3.135 ;
        RECT 4.585 3.020 5.565 3.145 ;
        RECT 4.595 3.020 5.565 3.155 ;
        RECT 3.975 2.915 4.605 3.085 ;
        RECT 4.605 3.020 5.565 3.165 ;
        RECT 3.975 2.925 4.615 3.085 ;
        RECT 4.615 3.020 5.565 3.175 ;
        RECT 3.975 2.935 4.625 3.085 ;
        RECT 4.625 3.020 5.565 3.184 ;
        RECT 3.975 2.940 4.631 3.085 ;
        RECT 3.975 2.950 4.640 3.085 ;
        RECT 3.975 2.960 4.650 3.085 ;
        RECT 3.975 2.970 4.660 3.085 ;
        RECT 3.975 2.980 4.670 3.085 ;
        RECT 3.975 2.990 4.680 3.085 ;
        RECT 3.975 3.000 4.690 3.085 ;
        RECT 3.975 3.010 4.700 3.085 ;
        RECT 4.630 3.020 5.565 3.190 ;
        RECT 6.850 1.610 7.020 1.970 ;
        RECT 5.845 1.795 7.020 1.970 ;
        RECT 6.825 0.830 7.495 1.065 ;
        RECT 4.675 0.880 4.975 2.370 ;
        RECT 4.675 2.150 5.015 2.370 ;
        RECT 7.355 1.630 7.525 2.360 ;
        RECT 4.675 2.150 7.525 2.360 ;
        RECT 7.460 1.625 7.995 1.800 ;
        RECT 7.355 1.630 7.995 1.800 ;
        RECT 5.365 1.245 5.665 1.760 ;
        RECT 7.695 0.775 7.865 1.430 ;
        RECT 5.365 1.245 7.865 1.430 ;
        RECT 7.695 0.775 9.380 0.945 ;
        RECT 9.210 0.775 9.380 2.555 ;
        RECT 9.025 2.045 9.380 2.555 ;
        RECT 9.210 1.515 10.540 1.815 ;
  END 
END LATNSRHD2XHT

MACRO MUX2HD2XHT
  CLASS  CORE ;
  FOREIGN MUX2HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.510 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.900 1.570 1.180 2.010 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.765 1.650 3.065 2.360 ;
        RECT 2.485 2.150 3.065 2.360 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.715 ;
        RECT 2.975 -0.300 3.275 1.055 ;
        RECT 4.080 -0.300 4.380 1.055 ;
        RECT 0.000 -0.300 4.510 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.510 0.545 3.830 1.055 ;
        RECT 3.660 0.545 3.830 3.030 ;
        RECT 3.595 2.010 3.830 3.030 ;
        RECT 3.660 1.670 4.000 2.120 ;
        RECT 3.595 2.010 4.000 2.120 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.635 0.955 3.990 ;
        RECT 2.635 2.975 3.275 3.990 ;
        RECT 4.050 2.295 4.350 3.990 ;
        RECT 0.000 3.390 4.510 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.400 1.420 2.585 1.520 ;
        RECT 0.520 1.220 0.690 1.885 ;
        RECT 0.440 1.570 0.690 1.885 ;
        RECT 0.520 1.220 1.570 1.390 ;
        RECT 1.330 0.860 1.570 1.390 ;
        RECT 0.520 1.350 2.455 1.390 ;
        RECT 1.400 0.860 1.570 2.010 ;
        RECT 2.285 1.350 2.455 1.590 ;
        RECT 1.400 1.350 2.455 1.520 ;
        RECT 2.285 1.420 2.585 1.590 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.090 1.110 0.260 2.360 ;
        RECT 0.170 0.980 0.340 1.280 ;
        RECT 0.090 1.110 0.340 1.280 ;
        RECT 1.880 1.720 2.050 2.360 ;
        RECT 0.090 2.190 2.050 2.360 ;
        RECT 1.545 2.545 1.845 3.055 ;
        RECT 1.860 0.530 2.030 1.170 ;
        RECT 1.860 1.000 2.590 1.170 ;
        RECT 2.965 1.300 3.480 1.470 ;
        RECT 3.245 1.650 3.415 2.715 ;
        RECT 1.545 2.545 3.415 2.715 ;
        RECT 3.310 1.300 3.480 1.870 ;
        RECT 3.245 1.650 3.480 1.870 ;
        RECT 2.890 1.235 2.900 1.469 ;
        RECT 2.900 1.245 2.910 1.469 ;
        RECT 2.910 1.255 2.920 1.469 ;
        RECT 2.920 1.265 2.930 1.469 ;
        RECT 2.930 1.275 2.940 1.469 ;
        RECT 2.940 1.285 2.950 1.469 ;
        RECT 2.950 1.295 2.960 1.469 ;
        RECT 2.960 1.300 2.966 1.470 ;
        RECT 2.665 1.010 2.675 1.244 ;
        RECT 2.675 1.020 2.685 1.254 ;
        RECT 2.685 1.030 2.695 1.264 ;
        RECT 2.695 1.040 2.705 1.274 ;
        RECT 2.705 1.050 2.715 1.284 ;
        RECT 2.715 1.060 2.725 1.294 ;
        RECT 2.725 1.070 2.735 1.304 ;
        RECT 2.735 1.080 2.745 1.314 ;
        RECT 2.745 1.090 2.755 1.324 ;
        RECT 2.755 1.100 2.765 1.334 ;
        RECT 2.765 1.110 2.775 1.344 ;
        RECT 2.775 1.120 2.785 1.354 ;
        RECT 2.785 1.130 2.795 1.364 ;
        RECT 2.795 1.140 2.805 1.374 ;
        RECT 2.805 1.150 2.815 1.384 ;
        RECT 2.815 1.160 2.825 1.394 ;
        RECT 2.825 1.170 2.835 1.404 ;
        RECT 2.835 1.180 2.845 1.414 ;
        RECT 2.845 1.190 2.855 1.424 ;
        RECT 2.855 1.200 2.865 1.434 ;
        RECT 2.865 1.210 2.875 1.444 ;
        RECT 2.875 1.220 2.885 1.454 ;
        RECT 2.885 1.225 2.891 1.465 ;
        RECT 2.590 1.000 2.600 1.170 ;
        RECT 2.600 1.000 2.610 1.180 ;
        RECT 2.610 1.000 2.620 1.190 ;
        RECT 2.620 1.000 2.630 1.200 ;
        RECT 2.630 1.000 2.640 1.210 ;
        RECT 2.640 1.000 2.650 1.220 ;
        RECT 2.650 1.000 2.660 1.230 ;
        RECT 2.660 1.000 2.666 1.240 ;
  END 
END MUX2HD2XHT

MACRO MUX2HD1XSPGHT
  CLASS  CORE ;
  FOREIGN MUX2HD1XSPGHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 1.575 0.300 2.115 3.055 ;
      LAYER V7 ;
        RECT 1.665 0.845 2.025 1.205 ;
      LAYER M7 ;
        RECT 1.495 0.835 2.355 1.215 ;
      LAYER V6 ;
        RECT 1.750 0.930 1.940 1.120 ;
      LAYER M4 ;
        RECT 2.155 0.840 2.355 2.200 ;
      LAYER V3 ;
        RECT 2.160 1.750 2.350 1.940 ;
      LAYER M3 ;
        RECT 1.680 1.745 2.420 1.945 ;
      LAYER V2 ;
        RECT 1.750 1.750 1.940 1.940 ;
      LAYER M2 ;
        RECT 1.745 1.220 1.945 2.200 ;
      LAYER V1 ;
        RECT 1.750 1.750 1.940 1.940 ;
      LAYER M1 ;
        RECT 1.740 1.475 2.000 2.010 ;
      LAYER M6 ;
        RECT 1.745 0.300 1.945 1.870 ;
      LAYER V5 ;
        RECT 1.750 0.930 1.940 1.120 ;
      LAYER M5 ;
        RECT 1.495 0.925 2.455 1.125 ;
      LAYER V4 ;
        RECT 2.160 0.930 2.350 1.120 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 4.035 0.300 4.575 3.065 ;
      LAYER V7 ;
        RECT 4.125 2.075 4.485 2.435 ;
      LAYER M7 ;
        RECT 3.600 2.065 4.575 2.445 ;
      LAYER V6 ;
        RECT 4.210 2.160 4.400 2.350 ;
      LAYER M4 ;
        RECT 3.795 1.980 3.995 2.850 ;
      LAYER V3 ;
        RECT 3.800 2.570 3.990 2.760 ;
      LAYER M3 ;
        RECT 2.895 2.565 4.100 2.765 ;
      LAYER V2 ;
        RECT 2.980 2.570 3.170 2.760 ;
      LAYER M2 ;
        RECT 2.975 1.870 3.175 2.850 ;
      LAYER V1 ;
        RECT 2.980 2.160 3.170 2.350 ;
      LAYER M1 ;
        RECT 2.970 1.845 3.270 2.420 ;
      LAYER M6 ;
        RECT 4.205 1.535 4.405 2.690 ;
      LAYER V5 ;
        RECT 4.210 2.160 4.400 2.350 ;
      LAYER M5 ;
        RECT 3.600 2.155 4.575 2.355 ;
      LAYER V4 ;
        RECT 3.800 2.160 3.990 2.350 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.445 -0.300 1.745 1.295 ;
        RECT 3.275 -0.300 3.575 1.055 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 2.805 0.300 3.345 3.060 ;
      LAYER V7 ;
        RECT 2.895 0.845 3.255 1.205 ;
      LAYER M7 ;
        RECT 2.725 0.835 3.725 1.215 ;
      LAYER V6 ;
        RECT 2.980 0.930 3.170 1.120 ;
      LAYER M4 ;
        RECT 3.385 0.840 3.585 1.715 ;
      LAYER V3 ;
        RECT 3.390 1.340 3.580 1.530 ;
      LAYER M3 ;
        RECT 3.300 1.335 4.480 1.535 ;
      LAYER V2 ;
        RECT 4.210 1.340 4.400 1.530 ;
      LAYER M2 ;
        RECT 4.205 1.250 4.405 2.015 ;
      LAYER V1 ;
        RECT 4.210 1.750 4.400 1.940 ;
      LAYER M1 ;
        RECT 3.890 0.720 4.030 2.960 ;
        RECT 3.860 1.980 4.030 2.960 ;
        RECT 3.890 0.720 4.060 2.210 ;
        RECT 3.860 1.980 4.060 2.210 ;
        RECT 3.860 0.720 4.070 1.360 ;
        RECT 3.890 1.625 4.410 2.015 ;
        RECT 3.860 1.980 4.410 2.015 ;
      LAYER M6 ;
        RECT 2.975 0.300 3.175 1.870 ;
      LAYER V5 ;
        RECT 2.980 0.930 3.170 1.120 ;
      LAYER M5 ;
        RECT 2.725 0.925 3.725 1.125 ;
      LAYER V4 ;
        RECT 3.390 0.930 3.580 1.120 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.445 2.545 1.745 3.990 ;
        RECT 3.275 2.635 3.575 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 0.345 0.300 0.885 3.070 ;
      LAYER V7 ;
        RECT 0.435 0.845 0.795 1.205 ;
      LAYER M7 ;
        RECT 0.200 0.835 0.885 1.215 ;
      LAYER V6 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M4 ;
        RECT 0.515 0.850 0.715 1.670 ;
      LAYER V3 ;
        RECT 0.520 1.340 0.710 1.530 ;
      LAYER M3 ;
        RECT 0.260 1.335 1.600 1.535 ;
      LAYER V2 ;
        RECT 1.340 1.340 1.530 1.530 ;
      LAYER M2 ;
        RECT 1.335 1.200 1.535 2.010 ;
      LAYER V1 ;
        RECT 1.340 1.750 1.530 1.940 ;
      LAYER M1 ;
        RECT 1.260 1.570 1.540 2.010 ;
      LAYER M6 ;
        RECT 0.515 0.300 0.715 1.870 ;
      LAYER V5 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M5 ;
        RECT 0.200 0.925 1.265 1.125 ;
      LAYER V4 ;
        RECT 0.520 0.930 0.710 1.120 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.910 1.190 1.080 2.595 ;
        RECT 0.990 1.060 1.160 1.360 ;
        RECT 0.910 1.190 1.160 1.360 ;
        RECT 0.910 2.190 1.225 2.595 ;
        RECT 2.220 1.560 2.390 2.360 ;
        RECT 0.910 2.190 2.390 2.360 ;
        RECT 2.335 1.125 2.740 1.295 ;
        RECT 2.570 1.125 2.740 2.715 ;
        RECT 2.335 2.545 2.740 2.715 ;
        RECT 2.570 1.475 3.710 1.645 ;
        RECT 3.540 1.475 3.710 1.870 ;
  END 
END MUX2HD1XSPGHT

MACRO MUX2CLKHD4XHT
  CLASS  CORE ;
  FOREIGN MUX2CLKHD4XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.380 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.900 1.575 1.230 2.020 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.605 1.225 4.875 1.745 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.025 ;
        RECT 2.795 -0.300 3.095 0.975 ;
        RECT 4.875 -0.300 5.175 1.025 ;
        RECT 5.935 -0.300 6.235 1.025 ;
        RECT 6.975 -0.300 7.275 1.045 ;
        RECT 0.000 -0.300 7.380 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.415 1.020 5.715 1.430 ;
        RECT 5.415 2.045 5.745 2.960 ;
        RECT 5.415 1.205 6.755 1.430 ;
        RECT 6.055 1.205 6.755 2.455 ;
        RECT 5.415 2.045 6.755 2.455 ;
        RECT 6.455 1.020 6.755 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.615 0.955 3.990 ;
        RECT 2.795 2.625 3.095 3.990 ;
        RECT 4.895 2.275 5.195 3.990 ;
        RECT 5.935 2.635 6.235 3.990 ;
        RECT 6.975 2.295 7.275 3.990 ;
        RECT 0.000 3.390 7.380 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.670 0.720 2.370 ;
        RECT 1.410 1.675 1.580 2.370 ;
        RECT 0.440 2.200 1.580 2.370 ;
        RECT 1.410 1.675 2.210 1.845 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 1.240 2.550 1.410 3.015 ;
        RECT 2.280 2.560 2.450 3.015 ;
        RECT 1.240 2.845 2.450 3.015 ;
        RECT 1.305 0.505 1.475 1.025 ;
        RECT 1.175 0.855 1.475 1.025 ;
        RECT 1.305 0.505 2.545 0.675 ;
        RECT 2.245 0.505 2.545 0.795 ;
        RECT 0.090 1.225 0.260 2.785 ;
        RECT 0.170 0.790 0.340 1.395 ;
        RECT 0.090 2.615 0.405 2.785 ;
        RECT 0.090 1.225 1.430 1.395 ;
        RECT 1.530 1.225 1.730 1.495 ;
        RECT 1.530 1.325 2.285 1.495 ;
        RECT 2.705 1.675 4.075 1.845 ;
        RECT 2.635 1.615 2.645 1.845 ;
        RECT 2.645 1.625 2.655 1.845 ;
        RECT 2.655 1.635 2.665 1.845 ;
        RECT 2.665 1.645 2.675 1.845 ;
        RECT 2.675 1.655 2.685 1.845 ;
        RECT 2.685 1.665 2.695 1.845 ;
        RECT 2.695 1.675 2.705 1.845 ;
        RECT 2.355 1.335 2.365 1.565 ;
        RECT 2.365 1.345 2.375 1.575 ;
        RECT 2.375 1.355 2.385 1.585 ;
        RECT 2.385 1.365 2.395 1.595 ;
        RECT 2.395 1.375 2.405 1.605 ;
        RECT 2.405 1.385 2.415 1.615 ;
        RECT 2.415 1.395 2.425 1.625 ;
        RECT 2.425 1.405 2.435 1.635 ;
        RECT 2.435 1.415 2.445 1.645 ;
        RECT 2.445 1.425 2.455 1.655 ;
        RECT 2.455 1.435 2.465 1.665 ;
        RECT 2.465 1.445 2.475 1.675 ;
        RECT 2.475 1.455 2.485 1.685 ;
        RECT 2.485 1.465 2.495 1.695 ;
        RECT 2.495 1.475 2.505 1.705 ;
        RECT 2.505 1.485 2.515 1.715 ;
        RECT 2.515 1.495 2.525 1.725 ;
        RECT 2.525 1.505 2.535 1.735 ;
        RECT 2.535 1.515 2.545 1.745 ;
        RECT 2.545 1.525 2.555 1.755 ;
        RECT 2.555 1.535 2.565 1.765 ;
        RECT 2.565 1.545 2.575 1.775 ;
        RECT 2.575 1.555 2.585 1.785 ;
        RECT 2.585 1.565 2.595 1.795 ;
        RECT 2.595 1.575 2.605 1.805 ;
        RECT 2.605 1.585 2.615 1.815 ;
        RECT 2.615 1.595 2.625 1.825 ;
        RECT 2.625 1.605 2.635 1.835 ;
        RECT 2.285 1.325 2.295 1.495 ;
        RECT 2.295 1.325 2.305 1.505 ;
        RECT 2.305 1.325 2.315 1.515 ;
        RECT 2.315 1.325 2.325 1.525 ;
        RECT 2.325 1.325 2.335 1.535 ;
        RECT 2.335 1.325 2.345 1.545 ;
        RECT 2.345 1.325 2.355 1.555 ;
        RECT 1.430 1.225 1.440 1.395 ;
        RECT 1.440 1.225 1.450 1.405 ;
        RECT 1.450 1.225 1.460 1.415 ;
        RECT 1.460 1.225 1.470 1.425 ;
        RECT 1.470 1.225 1.480 1.435 ;
        RECT 1.480 1.225 1.490 1.445 ;
        RECT 1.490 1.225 1.500 1.455 ;
        RECT 1.500 1.225 1.510 1.465 ;
        RECT 1.510 1.225 1.520 1.475 ;
        RECT 1.520 1.225 1.530 1.485 ;
        RECT 3.380 2.560 3.550 3.015 ;
        RECT 4.420 2.550 4.590 3.015 ;
        RECT 3.380 2.845 4.590 3.015 ;
        RECT 3.445 0.505 3.615 0.975 ;
        RECT 3.315 0.805 3.615 0.975 ;
        RECT 3.445 0.505 4.655 0.675 ;
        RECT 4.355 0.505 4.655 1.025 ;
        RECT 1.760 2.025 1.930 2.665 ;
        RECT 1.905 0.855 2.075 1.145 ;
        RECT 1.690 0.855 2.075 1.025 ;
        RECT 1.905 0.975 2.460 1.145 ;
        RECT 3.900 2.025 4.070 2.665 ;
        RECT 3.835 0.855 4.135 1.445 ;
        RECT 2.710 1.155 4.135 1.325 ;
        RECT 3.835 1.275 4.425 1.445 ;
        RECT 4.255 1.275 4.425 2.195 ;
        RECT 1.760 2.025 4.425 2.195 ;
        RECT 4.255 1.925 5.235 2.095 ;
        RECT 5.065 1.610 5.235 2.095 ;
        RECT 5.065 1.610 5.875 1.780 ;
        RECT 2.640 1.095 2.650 1.325 ;
        RECT 2.650 1.105 2.660 1.325 ;
        RECT 2.660 1.115 2.670 1.325 ;
        RECT 2.670 1.125 2.680 1.325 ;
        RECT 2.680 1.135 2.690 1.325 ;
        RECT 2.690 1.145 2.700 1.325 ;
        RECT 2.700 1.155 2.710 1.325 ;
        RECT 2.530 0.985 2.540 1.215 ;
        RECT 2.540 0.995 2.550 1.225 ;
        RECT 2.550 1.005 2.560 1.235 ;
        RECT 2.560 1.015 2.570 1.245 ;
        RECT 2.570 1.025 2.580 1.255 ;
        RECT 2.580 1.035 2.590 1.265 ;
        RECT 2.590 1.045 2.600 1.275 ;
        RECT 2.600 1.055 2.610 1.285 ;
        RECT 2.610 1.065 2.620 1.295 ;
        RECT 2.620 1.075 2.630 1.305 ;
        RECT 2.630 1.085 2.640 1.315 ;
        RECT 2.460 0.975 2.470 1.145 ;
        RECT 2.470 0.975 2.480 1.155 ;
        RECT 2.480 0.975 2.490 1.165 ;
        RECT 2.490 0.975 2.500 1.175 ;
        RECT 2.500 0.975 2.510 1.185 ;
        RECT 2.510 0.975 2.520 1.195 ;
        RECT 2.520 0.975 2.530 1.205 ;
  END 
END MUX2CLKHD4XHT

MACRO MUX2CLKHD3XHT
  CLASS  CORE ;
  FOREIGN MUX2CLKHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.270 1.220 2.085 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.560 1.610 2.925 2.050 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.995 ;
        RECT 2.840 -0.300 3.140 0.995 ;
        RECT 3.915 -0.300 4.215 0.995 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.395 0.910 3.695 1.080 ;
        RECT 3.460 1.980 3.630 2.960 ;
        RECT 3.525 0.910 3.695 1.385 ;
        RECT 3.525 1.215 4.735 1.385 ;
        RECT 4.035 1.215 4.735 2.455 ;
        RECT 3.460 1.980 4.735 2.455 ;
        RECT 4.435 1.060 4.735 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.635 0.955 3.990 ;
        RECT 2.865 2.635 3.165 3.990 ;
        RECT 3.915 2.635 4.215 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.260 0.720 1.985 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.090 0.845 0.260 2.455 ;
        RECT 0.090 0.845 0.405 1.080 ;
        RECT 0.090 2.165 0.405 2.455 ;
        RECT 1.400 1.290 1.570 2.455 ;
        RECT 0.090 2.285 1.570 2.455 ;
        RECT 1.400 1.290 1.580 1.960 ;
        RECT 2.210 1.610 2.380 1.960 ;
        RECT 1.400 1.790 2.380 1.960 ;
        RECT 1.870 2.230 2.040 3.210 ;
        RECT 1.685 0.930 2.495 1.100 ;
        RECT 2.325 0.930 2.495 1.430 ;
        RECT 2.325 1.260 3.280 1.430 ;
        RECT 3.110 1.260 3.280 2.400 ;
        RECT 1.870 2.230 3.280 2.400 ;
        RECT 3.110 1.565 3.855 1.735 ;
  END 
END MUX2CLKHD3XHT

MACRO MUX2CLKHD2XHT
  CLASS  CORE ;
  FOREIGN MUX2CLKHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.270 1.180 2.020 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.675 2.360 2.430 ;
        RECT 2.150 1.675 2.555 1.845 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.065 ;
        RECT 2.500 -0.300 2.670 1.130 ;
        RECT 3.570 -0.300 3.740 1.000 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.900 0.895 3.370 1.130 ;
        RECT 3.170 0.895 3.370 2.960 ;
        RECT 3.050 1.980 3.370 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.555 0.955 3.990 ;
        RECT 2.465 2.635 2.765 3.990 ;
        RECT 3.570 2.230 3.740 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.260 0.720 1.960 ;
    END
  END S0
  OBS 
      LAYER M1 ;
        RECT 0.090 0.895 0.260 2.370 ;
        RECT 0.090 0.895 0.405 1.065 ;
        RECT 0.090 2.175 0.405 2.370 ;
        RECT 1.400 1.330 1.570 2.370 ;
        RECT 0.090 2.200 1.570 2.370 ;
        RECT 1.540 0.895 1.945 1.065 ;
        RECT 1.775 0.895 1.945 2.725 ;
        RECT 1.540 2.555 1.945 2.725 ;
        RECT 1.775 1.325 2.970 1.495 ;
        RECT 2.800 1.325 2.970 1.770 ;
  END 
END MUX2CLKHD2XHT

MACRO LATTSHDMXHT
  CLASS  CORE ;
  FOREIGN LATTSHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.560 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 4.555 0.850 4.725 2.280 ;
        RECT 4.555 0.850 4.820 1.205 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.670 1.520 2.090 1.950 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.770 1.520 6.055 2.020 ;
    END
  END E
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.490 0.520 2.950 ;
    END
  END G
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 1.580 -0.300 1.880 0.815 ;
        RECT 3.605 -0.300 3.775 0.810 ;
        RECT 5.380 -0.300 5.680 1.295 ;
        RECT 0.000 -0.300 6.560 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.700 3.030 1.000 3.990 ;
        RECT 1.625 3.030 1.925 3.990 ;
        RECT 3.490 2.935 3.790 3.990 ;
        RECT 5.475 2.520 5.645 3.990 ;
        RECT 0.000 3.390 6.560 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.590 1.030 1.760 ;
        RECT 0.860 1.520 1.030 2.850 ;
        RECT 0.860 2.680 2.010 2.850 ;
        RECT 2.335 2.930 2.640 3.100 ;
        RECT 2.260 2.865 2.270 3.099 ;
        RECT 2.270 2.875 2.280 3.099 ;
        RECT 2.280 2.885 2.290 3.099 ;
        RECT 2.290 2.895 2.300 3.099 ;
        RECT 2.300 2.905 2.310 3.099 ;
        RECT 2.310 2.915 2.320 3.099 ;
        RECT 2.320 2.925 2.330 3.099 ;
        RECT 2.330 2.930 2.336 3.100 ;
        RECT 2.085 2.690 2.095 2.924 ;
        RECT 2.095 2.700 2.105 2.934 ;
        RECT 2.105 2.710 2.115 2.944 ;
        RECT 2.115 2.720 2.125 2.954 ;
        RECT 2.125 2.730 2.135 2.964 ;
        RECT 2.135 2.740 2.145 2.974 ;
        RECT 2.145 2.750 2.155 2.984 ;
        RECT 2.155 2.760 2.165 2.994 ;
        RECT 2.165 2.770 2.175 3.004 ;
        RECT 2.175 2.780 2.185 3.014 ;
        RECT 2.185 2.790 2.195 3.024 ;
        RECT 2.195 2.800 2.205 3.034 ;
        RECT 2.205 2.810 2.215 3.044 ;
        RECT 2.215 2.820 2.225 3.054 ;
        RECT 2.225 2.830 2.235 3.064 ;
        RECT 2.235 2.840 2.245 3.074 ;
        RECT 2.245 2.850 2.255 3.084 ;
        RECT 2.255 2.855 2.261 3.095 ;
        RECT 2.010 2.680 2.020 2.850 ;
        RECT 2.020 2.680 2.030 2.860 ;
        RECT 2.030 2.680 2.040 2.870 ;
        RECT 2.040 2.680 2.050 2.880 ;
        RECT 2.050 2.680 2.060 2.890 ;
        RECT 2.060 2.680 2.070 2.900 ;
        RECT 2.070 2.680 2.080 2.910 ;
        RECT 2.080 2.680 2.086 2.920 ;
        RECT 1.210 1.060 1.380 2.500 ;
        RECT 1.210 2.330 2.200 2.500 ;
        RECT 2.125 0.605 2.295 1.230 ;
        RECT 1.210 1.060 2.295 1.230 ;
        RECT 2.125 0.605 2.630 0.775 ;
        RECT 2.525 2.580 3.085 2.750 ;
        RECT 2.915 2.580 3.085 3.115 ;
        RECT 2.450 2.515 2.460 2.749 ;
        RECT 2.460 2.525 2.470 2.749 ;
        RECT 2.470 2.535 2.480 2.749 ;
        RECT 2.480 2.545 2.490 2.749 ;
        RECT 2.490 2.555 2.500 2.749 ;
        RECT 2.500 2.565 2.510 2.749 ;
        RECT 2.510 2.575 2.520 2.749 ;
        RECT 2.520 2.580 2.526 2.750 ;
        RECT 2.275 2.340 2.285 2.574 ;
        RECT 2.285 2.350 2.295 2.584 ;
        RECT 2.295 2.360 2.305 2.594 ;
        RECT 2.305 2.370 2.315 2.604 ;
        RECT 2.315 2.380 2.325 2.614 ;
        RECT 2.325 2.390 2.335 2.624 ;
        RECT 2.335 2.400 2.345 2.634 ;
        RECT 2.345 2.410 2.355 2.644 ;
        RECT 2.355 2.420 2.365 2.654 ;
        RECT 2.365 2.430 2.375 2.664 ;
        RECT 2.375 2.440 2.385 2.674 ;
        RECT 2.385 2.450 2.395 2.684 ;
        RECT 2.395 2.460 2.405 2.694 ;
        RECT 2.405 2.470 2.415 2.704 ;
        RECT 2.415 2.480 2.425 2.714 ;
        RECT 2.425 2.490 2.435 2.724 ;
        RECT 2.435 2.500 2.445 2.734 ;
        RECT 2.445 2.505 2.451 2.745 ;
        RECT 2.200 2.330 2.210 2.500 ;
        RECT 2.210 2.330 2.220 2.510 ;
        RECT 2.220 2.330 2.230 2.520 ;
        RECT 2.230 2.330 2.240 2.530 ;
        RECT 2.240 2.330 2.250 2.540 ;
        RECT 2.250 2.330 2.260 2.550 ;
        RECT 2.260 2.330 2.270 2.560 ;
        RECT 2.270 2.330 2.276 2.570 ;
        RECT 3.235 0.480 3.405 1.230 ;
        RECT 3.235 1.060 4.215 1.230 ;
        RECT 4.045 1.060 4.215 2.385 ;
        RECT 2.510 1.125 2.810 1.295 ;
        RECT 2.635 1.125 2.805 2.385 ;
        RECT 2.635 1.125 2.810 1.780 ;
        RECT 2.635 1.610 3.865 1.780 ;
        RECT 3.695 1.610 3.865 2.735 ;
        RECT 5.000 1.585 5.170 2.735 ;
        RECT 3.695 2.565 5.170 2.735 ;
        RECT 5.000 1.585 5.500 1.755 ;
        RECT 5.825 2.200 5.995 3.190 ;
        RECT 5.900 1.125 6.405 1.295 ;
        RECT 6.235 1.125 6.405 2.370 ;
        RECT 5.825 2.200 6.405 2.370 ;
  END 
END LATTSHDMXHT

MACRO LATTSHDLXHT
  CLASS  CORE ;
  FOREIGN LATTSHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.560 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 4.610 1.060 4.845 1.670 ;
        RECT 4.675 1.060 4.845 2.280 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.670 1.520 2.210 1.950 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.765 1.540 6.120 1.950 ;
    END
  END E
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.490 0.520 2.855 ;
    END
  END G
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.825 ;
        RECT 1.655 -0.300 1.955 0.880 ;
        RECT 3.725 -0.300 3.895 0.810 ;
        RECT 5.500 -0.300 5.800 1.295 ;
        RECT 0.000 -0.300 6.560 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.700 3.030 1.000 3.990 ;
        RECT 1.745 3.030 2.045 3.990 ;
        RECT 3.610 2.830 3.910 3.990 ;
        RECT 5.565 2.250 5.735 3.990 ;
        RECT 0.000 3.390 6.560 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.590 1.030 1.760 ;
        RECT 0.860 1.520 1.030 2.850 ;
        RECT 0.860 2.680 2.130 2.850 ;
        RECT 2.475 2.950 2.650 3.120 ;
        RECT 2.350 2.835 2.360 3.119 ;
        RECT 2.360 2.845 2.370 3.119 ;
        RECT 2.370 2.855 2.380 3.119 ;
        RECT 2.380 2.865 2.390 3.119 ;
        RECT 2.390 2.875 2.400 3.119 ;
        RECT 2.400 2.885 2.410 3.119 ;
        RECT 2.410 2.895 2.420 3.119 ;
        RECT 2.420 2.905 2.430 3.119 ;
        RECT 2.430 2.915 2.440 3.119 ;
        RECT 2.440 2.925 2.450 3.119 ;
        RECT 2.450 2.935 2.460 3.119 ;
        RECT 2.460 2.945 2.470 3.119 ;
        RECT 2.470 2.950 2.476 3.120 ;
        RECT 2.205 2.690 2.215 2.924 ;
        RECT 2.215 2.700 2.225 2.934 ;
        RECT 2.225 2.710 2.235 2.944 ;
        RECT 2.235 2.720 2.245 2.954 ;
        RECT 2.245 2.730 2.255 2.964 ;
        RECT 2.255 2.740 2.265 2.974 ;
        RECT 2.265 2.750 2.275 2.984 ;
        RECT 2.275 2.760 2.285 2.994 ;
        RECT 2.285 2.770 2.295 3.004 ;
        RECT 2.295 2.780 2.305 3.014 ;
        RECT 2.305 2.790 2.315 3.024 ;
        RECT 2.315 2.800 2.325 3.034 ;
        RECT 2.325 2.810 2.335 3.044 ;
        RECT 2.335 2.820 2.345 3.054 ;
        RECT 2.345 2.825 2.351 3.065 ;
        RECT 2.130 2.680 2.140 2.850 ;
        RECT 2.140 2.680 2.150 2.860 ;
        RECT 2.150 2.680 2.160 2.870 ;
        RECT 2.160 2.680 2.170 2.880 ;
        RECT 2.170 2.680 2.180 2.890 ;
        RECT 2.180 2.680 2.190 2.900 ;
        RECT 2.190 2.680 2.200 2.910 ;
        RECT 2.200 2.680 2.206 2.920 ;
        RECT 1.210 1.060 1.380 2.500 ;
        RECT 1.210 2.330 2.320 2.500 ;
        RECT 2.190 0.630 2.360 1.230 ;
        RECT 1.210 1.060 2.360 1.230 ;
        RECT 2.190 0.630 2.695 0.800 ;
        RECT 2.665 2.600 3.170 2.770 ;
        RECT 2.590 2.535 2.600 2.769 ;
        RECT 2.600 2.545 2.610 2.769 ;
        RECT 2.610 2.555 2.620 2.769 ;
        RECT 2.620 2.565 2.630 2.769 ;
        RECT 2.630 2.575 2.640 2.769 ;
        RECT 2.640 2.585 2.650 2.769 ;
        RECT 2.650 2.595 2.660 2.769 ;
        RECT 2.660 2.600 2.666 2.770 ;
        RECT 2.395 2.340 2.405 2.574 ;
        RECT 2.405 2.350 2.415 2.584 ;
        RECT 2.415 2.360 2.425 2.594 ;
        RECT 2.425 2.370 2.435 2.604 ;
        RECT 2.435 2.380 2.445 2.614 ;
        RECT 2.445 2.390 2.455 2.624 ;
        RECT 2.455 2.400 2.465 2.634 ;
        RECT 2.465 2.410 2.475 2.644 ;
        RECT 2.475 2.420 2.485 2.654 ;
        RECT 2.485 2.430 2.495 2.664 ;
        RECT 2.495 2.440 2.505 2.674 ;
        RECT 2.505 2.450 2.515 2.684 ;
        RECT 2.515 2.460 2.525 2.694 ;
        RECT 2.525 2.470 2.535 2.704 ;
        RECT 2.535 2.480 2.545 2.714 ;
        RECT 2.545 2.490 2.555 2.724 ;
        RECT 2.555 2.500 2.565 2.734 ;
        RECT 2.565 2.510 2.575 2.744 ;
        RECT 2.575 2.520 2.585 2.754 ;
        RECT 2.585 2.525 2.591 2.765 ;
        RECT 2.320 2.330 2.330 2.500 ;
        RECT 2.330 2.330 2.340 2.510 ;
        RECT 2.340 2.330 2.350 2.520 ;
        RECT 2.350 2.330 2.360 2.530 ;
        RECT 2.360 2.330 2.370 2.540 ;
        RECT 2.370 2.330 2.380 2.550 ;
        RECT 2.380 2.330 2.390 2.560 ;
        RECT 2.390 2.330 2.396 2.570 ;
        RECT 3.355 0.615 3.525 1.230 ;
        RECT 3.355 1.060 4.335 1.230 ;
        RECT 4.165 1.060 4.335 2.300 ;
        RECT 2.605 1.125 2.925 1.295 ;
        RECT 2.755 1.125 2.925 2.420 ;
        RECT 2.755 1.610 3.985 1.780 ;
        RECT 3.815 1.610 3.985 2.650 ;
        RECT 5.105 1.585 5.275 2.650 ;
        RECT 3.815 2.480 5.275 2.650 ;
        RECT 5.105 1.585 5.585 1.755 ;
        RECT 6.060 1.060 6.470 1.360 ;
        RECT 6.060 2.165 6.470 2.335 ;
        RECT 6.300 1.060 6.470 3.005 ;
        RECT 5.915 2.820 6.470 3.005 ;
  END 
END LATTSHDLXHT

MACRO LATTSHD2XHT
  CLASS  CORE ;
  FOREIGN LATTSHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.430 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 8.570 0.720 8.740 2.960 ;
        RECT 8.570 1.330 8.990 1.540 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.625 1.520 2.045 1.950 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.250 1.495 6.695 2.025 ;
    END
  END E
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.490 0.520 2.950 ;
    END
  END G
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 1.535 -0.300 1.835 0.770 ;
        RECT 3.560 -0.300 3.730 0.810 ;
        RECT 4.905 -0.300 5.205 0.715 ;
        RECT 5.975 -0.300 6.275 0.595 ;
        RECT 8.050 -0.300 8.220 1.120 ;
        RECT 9.025 -0.300 9.325 1.055 ;
        RECT 0.000 -0.300 9.430 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.700 3.030 1.000 3.990 ;
        RECT 1.580 3.030 1.880 3.990 ;
        RECT 3.415 2.270 3.715 3.990 ;
        RECT 4.905 2.975 5.205 3.990 ;
        RECT 5.975 3.030 6.275 3.990 ;
        RECT 7.985 2.295 8.285 3.990 ;
        RECT 9.025 2.295 9.325 3.990 ;
        RECT 0.000 3.390 9.430 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.590 1.030 1.760 ;
        RECT 0.860 1.520 1.030 2.850 ;
        RECT 0.860 2.680 1.965 2.850 ;
        RECT 2.290 2.930 2.595 3.100 ;
        RECT 2.215 2.865 2.225 3.099 ;
        RECT 2.225 2.875 2.235 3.099 ;
        RECT 2.235 2.885 2.245 3.099 ;
        RECT 2.245 2.895 2.255 3.099 ;
        RECT 2.255 2.905 2.265 3.099 ;
        RECT 2.265 2.915 2.275 3.099 ;
        RECT 2.275 2.925 2.285 3.099 ;
        RECT 2.285 2.930 2.291 3.100 ;
        RECT 2.040 2.690 2.050 2.924 ;
        RECT 2.050 2.700 2.060 2.934 ;
        RECT 2.060 2.710 2.070 2.944 ;
        RECT 2.070 2.720 2.080 2.954 ;
        RECT 2.080 2.730 2.090 2.964 ;
        RECT 2.090 2.740 2.100 2.974 ;
        RECT 2.100 2.750 2.110 2.984 ;
        RECT 2.110 2.760 2.120 2.994 ;
        RECT 2.120 2.770 2.130 3.004 ;
        RECT 2.130 2.780 2.140 3.014 ;
        RECT 2.140 2.790 2.150 3.024 ;
        RECT 2.150 2.800 2.160 3.034 ;
        RECT 2.160 2.810 2.170 3.044 ;
        RECT 2.170 2.820 2.180 3.054 ;
        RECT 2.180 2.830 2.190 3.064 ;
        RECT 2.190 2.840 2.200 3.074 ;
        RECT 2.200 2.850 2.210 3.084 ;
        RECT 2.210 2.855 2.216 3.095 ;
        RECT 1.965 2.680 1.975 2.850 ;
        RECT 1.975 2.680 1.985 2.860 ;
        RECT 1.985 2.680 1.995 2.870 ;
        RECT 1.995 2.680 2.005 2.880 ;
        RECT 2.005 2.680 2.015 2.890 ;
        RECT 2.015 2.680 2.025 2.900 ;
        RECT 2.025 2.680 2.035 2.910 ;
        RECT 2.035 2.680 2.041 2.920 ;
        RECT 1.210 1.060 1.380 2.500 ;
        RECT 1.210 2.330 2.155 2.500 ;
        RECT 2.065 0.710 2.235 1.230 ;
        RECT 1.210 1.060 2.235 1.230 ;
        RECT 2.065 0.710 2.585 0.880 ;
        RECT 2.480 2.580 3.105 2.750 ;
        RECT 2.805 2.580 3.105 3.050 ;
        RECT 2.405 2.515 2.415 2.749 ;
        RECT 2.415 2.525 2.425 2.749 ;
        RECT 2.425 2.535 2.435 2.749 ;
        RECT 2.435 2.545 2.445 2.749 ;
        RECT 2.445 2.555 2.455 2.749 ;
        RECT 2.455 2.565 2.465 2.749 ;
        RECT 2.465 2.575 2.475 2.749 ;
        RECT 2.475 2.580 2.481 2.750 ;
        RECT 2.230 2.340 2.240 2.574 ;
        RECT 2.240 2.350 2.250 2.584 ;
        RECT 2.250 2.360 2.260 2.594 ;
        RECT 2.260 2.370 2.270 2.604 ;
        RECT 2.270 2.380 2.280 2.614 ;
        RECT 2.280 2.390 2.290 2.624 ;
        RECT 2.290 2.400 2.300 2.634 ;
        RECT 2.300 2.410 2.310 2.644 ;
        RECT 2.310 2.420 2.320 2.654 ;
        RECT 2.320 2.430 2.330 2.664 ;
        RECT 2.330 2.440 2.340 2.674 ;
        RECT 2.340 2.450 2.350 2.684 ;
        RECT 2.350 2.460 2.360 2.694 ;
        RECT 2.360 2.470 2.370 2.704 ;
        RECT 2.370 2.480 2.380 2.714 ;
        RECT 2.380 2.490 2.390 2.724 ;
        RECT 2.390 2.500 2.400 2.734 ;
        RECT 2.400 2.505 2.406 2.745 ;
        RECT 2.155 2.330 2.165 2.500 ;
        RECT 2.165 2.330 2.175 2.510 ;
        RECT 2.175 2.330 2.185 2.520 ;
        RECT 2.185 2.330 2.195 2.530 ;
        RECT 2.195 2.330 2.205 2.540 ;
        RECT 2.205 2.330 2.215 2.550 ;
        RECT 2.215 2.330 2.225 2.560 ;
        RECT 2.225 2.330 2.231 2.570 ;
        RECT 2.465 1.125 2.765 1.295 ;
        RECT 2.590 1.125 2.760 2.385 ;
        RECT 2.590 1.125 2.765 1.845 ;
        RECT 2.590 1.675 3.820 1.845 ;
        RECT 3.650 1.610 3.820 1.910 ;
        RECT 3.190 0.690 3.360 1.230 ;
        RECT 3.190 1.060 4.170 1.230 ;
        RECT 4.000 1.060 4.170 2.385 ;
        RECT 4.510 1.060 4.680 2.280 ;
        RECT 4.510 1.585 5.450 1.755 ;
        RECT 5.850 1.125 6.020 2.375 ;
        RECT 5.850 2.205 6.630 2.375 ;
        RECT 5.850 1.125 6.745 1.295 ;
        RECT 6.965 2.565 7.360 2.735 ;
        RECT 6.885 2.495 6.895 2.735 ;
        RECT 6.895 2.505 6.905 2.735 ;
        RECT 6.905 2.515 6.915 2.735 ;
        RECT 6.915 2.525 6.925 2.735 ;
        RECT 6.925 2.535 6.935 2.735 ;
        RECT 6.935 2.545 6.945 2.735 ;
        RECT 6.945 2.555 6.955 2.735 ;
        RECT 6.955 2.565 6.965 2.735 ;
        RECT 6.800 2.410 6.810 2.650 ;
        RECT 6.810 2.420 6.820 2.660 ;
        RECT 6.820 2.430 6.830 2.670 ;
        RECT 6.830 2.440 6.840 2.680 ;
        RECT 6.840 2.450 6.850 2.690 ;
        RECT 6.850 2.460 6.860 2.700 ;
        RECT 6.860 2.470 6.870 2.710 ;
        RECT 6.870 2.480 6.880 2.720 ;
        RECT 6.880 2.485 6.886 2.729 ;
        RECT 6.630 2.205 6.640 2.479 ;
        RECT 6.640 2.205 6.650 2.489 ;
        RECT 6.650 2.205 6.660 2.499 ;
        RECT 6.660 2.205 6.670 2.509 ;
        RECT 6.670 2.205 6.680 2.519 ;
        RECT 6.680 2.205 6.690 2.529 ;
        RECT 6.690 2.205 6.700 2.539 ;
        RECT 6.700 2.205 6.710 2.549 ;
        RECT 6.710 2.205 6.720 2.559 ;
        RECT 6.720 2.205 6.730 2.569 ;
        RECT 6.730 2.205 6.740 2.579 ;
        RECT 6.740 2.205 6.750 2.589 ;
        RECT 6.750 2.205 6.760 2.599 ;
        RECT 6.760 2.205 6.770 2.609 ;
        RECT 6.770 2.205 6.780 2.619 ;
        RECT 6.780 2.205 6.790 2.629 ;
        RECT 6.790 2.205 6.800 2.639 ;
        RECT 5.490 0.775 5.660 1.220 ;
        RECT 5.490 0.775 7.190 0.945 ;
        RECT 7.020 0.620 7.190 2.280 ;
        RECT 7.020 0.620 7.850 0.790 ;
        RECT 7.680 0.490 7.850 0.790 ;
        RECT 5.490 2.120 5.660 2.780 ;
        RECT 6.025 2.610 6.260 2.785 ;
        RECT 5.490 2.610 6.260 2.780 ;
        RECT 6.025 2.615 6.290 2.785 ;
        RECT 7.540 1.060 7.710 3.085 ;
        RECT 6.665 2.915 7.710 3.085 ;
        RECT 7.540 1.635 8.145 1.805 ;
        RECT 6.590 2.850 6.600 3.084 ;
        RECT 6.600 2.860 6.610 3.084 ;
        RECT 6.610 2.870 6.620 3.084 ;
        RECT 6.620 2.880 6.630 3.084 ;
        RECT 6.630 2.890 6.640 3.084 ;
        RECT 6.640 2.900 6.650 3.084 ;
        RECT 6.650 2.910 6.660 3.084 ;
        RECT 6.660 2.915 6.666 3.085 ;
        RECT 6.365 2.625 6.375 2.859 ;
        RECT 6.375 2.635 6.385 2.869 ;
        RECT 6.385 2.645 6.395 2.879 ;
        RECT 6.395 2.655 6.405 2.889 ;
        RECT 6.405 2.665 6.415 2.899 ;
        RECT 6.415 2.675 6.425 2.909 ;
        RECT 6.425 2.685 6.435 2.919 ;
        RECT 6.435 2.695 6.445 2.929 ;
        RECT 6.445 2.705 6.455 2.939 ;
        RECT 6.455 2.715 6.465 2.949 ;
        RECT 6.465 2.725 6.475 2.959 ;
        RECT 6.475 2.735 6.485 2.969 ;
        RECT 6.485 2.745 6.495 2.979 ;
        RECT 6.495 2.755 6.505 2.989 ;
        RECT 6.505 2.765 6.515 2.999 ;
        RECT 6.515 2.775 6.525 3.009 ;
        RECT 6.525 2.785 6.535 3.019 ;
        RECT 6.535 2.795 6.545 3.029 ;
        RECT 6.545 2.805 6.555 3.039 ;
        RECT 6.555 2.815 6.565 3.049 ;
        RECT 6.565 2.825 6.575 3.059 ;
        RECT 6.575 2.835 6.585 3.069 ;
        RECT 6.585 2.840 6.591 3.080 ;
        RECT 6.290 2.615 6.300 2.785 ;
        RECT 6.300 2.615 6.310 2.795 ;
        RECT 6.310 2.615 6.320 2.805 ;
        RECT 6.320 2.615 6.330 2.815 ;
        RECT 6.330 2.615 6.340 2.825 ;
        RECT 6.340 2.615 6.350 2.835 ;
        RECT 6.350 2.615 6.360 2.845 ;
        RECT 6.360 2.615 6.366 2.855 ;
  END 
END LATTSHD2XHT

MACRO LATTSHD1XHT
  CLASS  CORE ;
  FOREIGN LATTSHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.790 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 4.555 2.045 4.725 2.620 ;
        RECT 4.490 1.125 6.630 1.295 ;
        RECT 6.250 1.125 6.630 1.610 ;
        RECT 6.460 1.125 6.630 2.215 ;
        RECT 4.490 2.045 6.630 2.215 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.670 1.520 2.090 1.950 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.120 0.480 4.800 0.650 ;
        RECT 4.630 0.480 4.800 0.945 ;
        RECT 6.455 0.510 6.655 0.945 ;
        RECT 4.630 0.775 6.655 0.945 ;
        RECT 6.455 0.510 6.965 0.875 ;
        RECT 6.455 0.705 7.180 0.875 ;
        RECT 4.630 0.775 7.180 0.875 ;
    END
  END E
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.490 0.520 2.950 ;
    END
  END G
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 1.580 -0.300 1.880 0.815 ;
        RECT 3.605 -0.300 3.775 0.810 ;
        RECT 5.410 -0.300 5.710 0.595 ;
        RECT 7.360 -0.300 7.660 1.295 ;
        RECT 0.000 -0.300 7.790 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.700 3.030 1.000 3.990 ;
        RECT 1.625 3.030 1.925 3.990 ;
        RECT 3.460 2.270 3.760 3.990 ;
        RECT 5.410 2.925 5.710 3.990 ;
        RECT 7.360 2.165 7.660 3.990 ;
        RECT 0.000 3.390 7.790 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.590 1.030 1.760 ;
        RECT 0.860 1.520 1.030 2.850 ;
        RECT 0.860 2.680 2.010 2.850 ;
        RECT 2.335 2.930 2.640 3.100 ;
        RECT 2.260 2.865 2.270 3.099 ;
        RECT 2.270 2.875 2.280 3.099 ;
        RECT 2.280 2.885 2.290 3.099 ;
        RECT 2.290 2.895 2.300 3.099 ;
        RECT 2.300 2.905 2.310 3.099 ;
        RECT 2.310 2.915 2.320 3.099 ;
        RECT 2.320 2.925 2.330 3.099 ;
        RECT 2.330 2.930 2.336 3.100 ;
        RECT 2.085 2.690 2.095 2.924 ;
        RECT 2.095 2.700 2.105 2.934 ;
        RECT 2.105 2.710 2.115 2.944 ;
        RECT 2.115 2.720 2.125 2.954 ;
        RECT 2.125 2.730 2.135 2.964 ;
        RECT 2.135 2.740 2.145 2.974 ;
        RECT 2.145 2.750 2.155 2.984 ;
        RECT 2.155 2.760 2.165 2.994 ;
        RECT 2.165 2.770 2.175 3.004 ;
        RECT 2.175 2.780 2.185 3.014 ;
        RECT 2.185 2.790 2.195 3.024 ;
        RECT 2.195 2.800 2.205 3.034 ;
        RECT 2.205 2.810 2.215 3.044 ;
        RECT 2.215 2.820 2.225 3.054 ;
        RECT 2.225 2.830 2.235 3.064 ;
        RECT 2.235 2.840 2.245 3.074 ;
        RECT 2.245 2.850 2.255 3.084 ;
        RECT 2.255 2.855 2.261 3.095 ;
        RECT 2.010 2.680 2.020 2.850 ;
        RECT 2.020 2.680 2.030 2.860 ;
        RECT 2.030 2.680 2.040 2.870 ;
        RECT 2.040 2.680 2.050 2.880 ;
        RECT 2.050 2.680 2.060 2.890 ;
        RECT 2.060 2.680 2.070 2.900 ;
        RECT 2.070 2.680 2.080 2.910 ;
        RECT 2.080 2.680 2.086 2.920 ;
        RECT 1.210 1.060 1.380 2.500 ;
        RECT 1.210 2.330 2.200 2.500 ;
        RECT 2.095 0.605 2.265 1.230 ;
        RECT 1.210 1.060 2.265 1.230 ;
        RECT 2.095 0.605 2.620 0.775 ;
        RECT 2.525 2.580 3.150 2.750 ;
        RECT 2.850 2.580 3.150 3.050 ;
        RECT 2.450 2.515 2.460 2.749 ;
        RECT 2.460 2.525 2.470 2.749 ;
        RECT 2.470 2.535 2.480 2.749 ;
        RECT 2.480 2.545 2.490 2.749 ;
        RECT 2.490 2.555 2.500 2.749 ;
        RECT 2.500 2.565 2.510 2.749 ;
        RECT 2.510 2.575 2.520 2.749 ;
        RECT 2.520 2.580 2.526 2.750 ;
        RECT 2.275 2.340 2.285 2.574 ;
        RECT 2.285 2.350 2.295 2.584 ;
        RECT 2.295 2.360 2.305 2.594 ;
        RECT 2.305 2.370 2.315 2.604 ;
        RECT 2.315 2.380 2.325 2.614 ;
        RECT 2.325 2.390 2.335 2.624 ;
        RECT 2.335 2.400 2.345 2.634 ;
        RECT 2.345 2.410 2.355 2.644 ;
        RECT 2.355 2.420 2.365 2.654 ;
        RECT 2.365 2.430 2.375 2.664 ;
        RECT 2.375 2.440 2.385 2.674 ;
        RECT 2.385 2.450 2.395 2.684 ;
        RECT 2.395 2.460 2.405 2.694 ;
        RECT 2.405 2.470 2.415 2.704 ;
        RECT 2.415 2.480 2.425 2.714 ;
        RECT 2.425 2.490 2.435 2.724 ;
        RECT 2.435 2.500 2.445 2.734 ;
        RECT 2.445 2.505 2.451 2.745 ;
        RECT 2.200 2.330 2.210 2.500 ;
        RECT 2.210 2.330 2.220 2.510 ;
        RECT 2.220 2.330 2.230 2.520 ;
        RECT 2.230 2.330 2.240 2.530 ;
        RECT 2.240 2.330 2.250 2.540 ;
        RECT 2.250 2.330 2.260 2.550 ;
        RECT 2.260 2.330 2.270 2.560 ;
        RECT 2.270 2.330 2.276 2.570 ;
        RECT 2.510 1.125 2.810 1.295 ;
        RECT 2.635 1.125 2.805 2.385 ;
        RECT 2.635 1.125 2.810 1.845 ;
        RECT 2.635 1.675 3.865 1.845 ;
        RECT 3.695 1.610 3.865 1.910 ;
        RECT 3.235 0.655 3.405 1.230 ;
        RECT 3.235 1.060 4.215 1.230 ;
        RECT 4.045 1.060 4.215 2.385 ;
        RECT 4.415 1.520 4.585 1.820 ;
        RECT 4.415 1.585 5.880 1.755 ;
        RECT 5.000 2.510 5.170 3.170 ;
        RECT 4.120 3.000 5.170 3.170 ;
        RECT 6.765 2.510 6.935 3.170 ;
        RECT 6.905 1.060 7.075 2.680 ;
        RECT 5.000 2.510 7.075 2.680 ;
  END 
END LATTSHD1XHT

MACRO LATSRHDMXHT
  CLASS  CORE ;
  FOREIGN LATSRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.430 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.005 1.125 7.305 1.295 ;
        RECT 7.135 1.125 7.305 2.875 ;
        RECT 7.030 2.485 7.305 2.875 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.090 1.060 9.330 2.400 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.970 1.240 3.180 1.840 ;
        RECT 2.970 1.540 3.370 1.840 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.565 0.965 2.055 ;
    END
  END G
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.980 0.480 5.610 1.215 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 2.265 -0.300 2.565 0.595 ;
        RECT 5.790 -0.300 5.960 1.085 ;
        RECT 7.700 -0.300 8.005 0.745 ;
        RECT 8.505 -0.300 8.805 1.145 ;
        RECT 0.000 -0.300 9.430 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.490 2.745 2.035 3.180 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.905 0.895 3.990 ;
        RECT 2.270 2.745 2.440 3.990 ;
        RECT 5.695 2.610 5.865 3.990 ;
        RECT 5.630 2.610 5.930 2.780 ;
        RECT 7.490 2.220 7.790 3.990 ;
        RECT 8.505 2.495 8.805 3.990 ;
        RECT 0.000 3.390 9.430 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.655 1.125 2.550 1.295 ;
        RECT 2.380 1.125 2.550 2.215 ;
        RECT 1.655 2.045 2.550 2.215 ;
        RECT 3.420 1.125 3.720 1.295 ;
        RECT 3.550 1.125 3.720 2.370 ;
        RECT 3.240 2.200 3.720 2.370 ;
        RECT 1.210 0.775 1.380 2.215 ;
        RECT 1.145 2.045 1.445 2.215 ;
        RECT 2.975 0.605 3.145 0.945 ;
        RECT 1.210 0.775 3.145 0.945 ;
        RECT 2.975 0.605 4.080 0.775 ;
        RECT 0.105 1.125 0.275 2.565 ;
        RECT 0.105 1.125 0.405 1.295 ;
        RECT 0.105 2.345 0.405 2.565 ;
        RECT 1.075 2.395 1.245 2.950 ;
        RECT 2.880 2.395 3.060 2.720 ;
        RECT 0.105 2.395 3.060 2.565 ;
        RECT 3.925 0.975 4.095 2.860 ;
        RECT 2.880 2.550 4.095 2.720 ;
        RECT 3.925 0.975 4.140 1.145 ;
        RECT 3.925 2.690 4.340 2.860 ;
        RECT 4.630 0.705 4.800 1.020 ;
        RECT 4.340 0.850 4.800 1.020 ;
        RECT 4.265 0.850 4.275 1.084 ;
        RECT 4.275 0.850 4.285 1.074 ;
        RECT 4.285 0.850 4.295 1.064 ;
        RECT 4.295 0.850 4.305 1.054 ;
        RECT 4.305 0.850 4.315 1.044 ;
        RECT 4.315 0.850 4.325 1.034 ;
        RECT 4.325 0.850 4.335 1.024 ;
        RECT 4.335 0.850 4.341 1.020 ;
        RECT 4.215 0.900 4.225 1.134 ;
        RECT 4.225 0.890 4.235 1.124 ;
        RECT 4.235 0.880 4.245 1.114 ;
        RECT 4.245 0.870 4.255 1.104 ;
        RECT 4.255 0.860 4.265 1.094 ;
        RECT 4.140 0.975 4.150 1.145 ;
        RECT 4.150 0.965 4.160 1.145 ;
        RECT 4.160 0.955 4.170 1.145 ;
        RECT 4.170 0.945 4.180 1.145 ;
        RECT 4.180 0.935 4.190 1.145 ;
        RECT 4.190 0.925 4.200 1.145 ;
        RECT 4.200 0.915 4.210 1.145 ;
        RECT 4.210 0.905 4.216 1.145 ;
        RECT 2.640 2.890 2.810 3.190 ;
        RECT 3.670 3.040 5.515 3.120 ;
        RECT 3.680 3.040 5.515 3.130 ;
        RECT 3.690 3.040 5.515 3.140 ;
        RECT 3.700 3.040 4.690 3.150 ;
        RECT 3.710 3.040 4.690 3.160 ;
        RECT 3.720 3.040 4.690 3.170 ;
        RECT 3.730 3.040 4.690 3.180 ;
        RECT 3.740 3.040 4.690 3.190 ;
        RECT 2.640 2.940 3.750 3.110 ;
        RECT 3.750 3.040 4.690 3.200 ;
        RECT 2.640 2.950 3.760 3.110 ;
        RECT 2.640 2.960 3.770 3.110 ;
        RECT 2.640 2.970 3.780 3.110 ;
        RECT 2.640 2.980 3.790 3.110 ;
        RECT 2.640 2.990 3.800 3.110 ;
        RECT 2.640 3.000 3.810 3.110 ;
        RECT 2.640 3.010 3.820 3.110 ;
        RECT 2.640 3.020 3.830 3.110 ;
        RECT 2.640 3.030 3.840 3.110 ;
        RECT 4.520 2.975 4.690 3.210 ;
        RECT 3.760 3.040 4.690 3.210 ;
        RECT 4.520 2.975 5.515 3.145 ;
        RECT 5.215 2.975 5.515 3.210 ;
        RECT 4.340 1.275 4.510 2.370 ;
        RECT 4.340 1.275 4.640 1.445 ;
        RECT 6.490 1.060 6.785 1.360 ;
        RECT 6.615 1.060 6.785 2.370 ;
        RECT 4.280 2.200 6.785 2.370 ;
        RECT 6.615 1.565 6.925 1.865 ;
        RECT 6.140 0.710 6.310 1.930 ;
        RECT 4.970 1.735 6.310 1.930 ;
        RECT 6.140 0.710 7.320 0.880 ;
        RECT 7.655 1.125 8.295 1.295 ;
        RECT 8.080 1.125 8.250 2.335 ;
        RECT 8.080 1.125 8.295 1.780 ;
        RECT 8.080 1.480 8.910 1.780 ;
        RECT 7.485 0.800 7.495 1.294 ;
        RECT 7.495 0.810 7.505 1.294 ;
        RECT 7.505 0.820 7.515 1.294 ;
        RECT 7.515 0.830 7.525 1.294 ;
        RECT 7.525 0.840 7.535 1.294 ;
        RECT 7.535 0.850 7.545 1.294 ;
        RECT 7.545 0.860 7.555 1.294 ;
        RECT 7.555 0.870 7.565 1.294 ;
        RECT 7.565 0.880 7.575 1.294 ;
        RECT 7.575 0.890 7.585 1.294 ;
        RECT 7.585 0.900 7.595 1.294 ;
        RECT 7.595 0.910 7.605 1.294 ;
        RECT 7.605 0.920 7.615 1.294 ;
        RECT 7.615 0.930 7.625 1.294 ;
        RECT 7.625 0.940 7.635 1.294 ;
        RECT 7.635 0.950 7.645 1.294 ;
        RECT 7.645 0.960 7.655 1.294 ;
        RECT 7.405 0.720 7.415 0.964 ;
        RECT 7.415 0.730 7.425 0.974 ;
        RECT 7.425 0.740 7.435 0.984 ;
        RECT 7.435 0.750 7.445 0.994 ;
        RECT 7.445 0.760 7.455 1.004 ;
        RECT 7.455 0.770 7.465 1.014 ;
        RECT 7.465 0.780 7.475 1.024 ;
        RECT 7.475 0.790 7.485 1.034 ;
        RECT 7.320 0.710 7.330 0.880 ;
        RECT 7.330 0.710 7.340 0.890 ;
        RECT 7.340 0.710 7.350 0.900 ;
        RECT 7.350 0.710 7.360 0.910 ;
        RECT 7.360 0.710 7.370 0.920 ;
        RECT 7.370 0.710 7.380 0.930 ;
        RECT 7.380 0.710 7.390 0.940 ;
        RECT 7.390 0.710 7.400 0.950 ;
        RECT 7.400 0.710 7.406 0.960 ;
  END 
END LATSRHDMXHT

MACRO LATSRHDLXHT
  CLASS  CORE ;
  FOREIGN LATSRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.020 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 6.660 1.505 7.065 1.675 ;
        RECT 6.895 1.125 6.985 2.280 ;
        RECT 6.660 1.125 6.985 1.675 ;
        RECT 6.895 1.505 7.065 2.280 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.615 1.125 8.920 1.295 ;
        RECT 8.710 1.125 8.920 2.910 ;
        RECT 8.515 2.610 8.920 2.910 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.960 1.235 3.180 1.950 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.565 0.965 2.030 ;
    END
  END G
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.770 0.480 5.360 0.720 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.685 -0.300 0.985 1.295 ;
        RECT 2.225 -0.300 2.525 0.595 ;
        RECT 5.540 -0.300 5.710 1.360 ;
        RECT 7.555 -0.300 8.065 0.810 ;
        RECT 0.000 -0.300 9.020 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.560 2.855 2.035 3.180 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.855 0.895 3.990 ;
        RECT 2.240 2.855 2.440 3.990 ;
        RECT 5.400 2.420 5.700 3.990 ;
        RECT 7.415 2.100 7.585 3.990 ;
        RECT 7.995 2.730 8.165 3.990 ;
        RECT 0.000 3.390 9.020 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.775 1.125 2.230 1.295 ;
        RECT 2.060 1.125 2.230 2.325 ;
        RECT 1.655 2.155 2.230 2.325 ;
        RECT 2.060 1.785 2.715 1.955 ;
        RECT 3.360 1.060 3.530 2.390 ;
        RECT 1.275 0.775 1.445 2.215 ;
        RECT 1.145 2.045 1.445 2.215 ;
        RECT 1.275 0.775 1.500 1.360 ;
        RECT 2.975 0.605 3.145 0.945 ;
        RECT 1.275 0.775 3.145 0.945 ;
        RECT 2.975 0.605 3.715 0.775 ;
        RECT 0.105 1.125 0.275 2.675 ;
        RECT 0.105 1.125 0.405 1.295 ;
        RECT 0.105 2.185 0.405 2.675 ;
        RECT 0.105 2.490 1.245 2.675 ;
        RECT 1.075 2.490 1.245 2.790 ;
        RECT 0.105 2.505 3.170 2.675 ;
        RECT 3.005 2.570 3.710 2.740 ;
        RECT 3.635 2.570 3.710 2.795 ;
        RECT 3.880 2.570 3.935 2.795 ;
        RECT 4.265 0.605 4.580 0.955 ;
        RECT 4.060 0.785 4.580 0.955 ;
        RECT 3.965 0.785 3.975 1.039 ;
        RECT 3.975 0.785 3.985 1.029 ;
        RECT 3.985 0.785 3.995 1.019 ;
        RECT 3.995 0.785 4.005 1.009 ;
        RECT 4.005 0.785 4.015 0.999 ;
        RECT 4.015 0.785 4.025 0.989 ;
        RECT 4.025 0.785 4.035 0.979 ;
        RECT 4.035 0.785 4.045 0.969 ;
        RECT 4.045 0.785 4.055 0.959 ;
        RECT 4.055 0.785 4.061 0.955 ;
        RECT 3.880 0.870 3.890 1.124 ;
        RECT 3.890 0.860 3.900 1.114 ;
        RECT 3.900 0.850 3.910 1.104 ;
        RECT 3.910 0.840 3.920 1.094 ;
        RECT 3.920 0.830 3.930 1.084 ;
        RECT 3.930 0.820 3.940 1.074 ;
        RECT 3.940 0.810 3.950 1.064 ;
        RECT 3.950 0.800 3.960 1.054 ;
        RECT 3.960 0.790 3.966 1.050 ;
        RECT 3.710 1.040 3.720 2.794 ;
        RECT 3.720 1.030 3.730 2.794 ;
        RECT 3.730 1.020 3.740 2.794 ;
        RECT 3.740 1.010 3.750 2.794 ;
        RECT 3.750 1.000 3.760 2.794 ;
        RECT 3.760 0.990 3.770 2.794 ;
        RECT 3.770 0.980 3.780 2.794 ;
        RECT 3.780 0.970 3.790 2.794 ;
        RECT 3.790 0.960 3.800 2.794 ;
        RECT 3.800 0.950 3.810 2.794 ;
        RECT 3.810 0.940 3.820 2.794 ;
        RECT 3.820 0.930 3.830 2.794 ;
        RECT 3.830 0.920 3.840 2.794 ;
        RECT 3.840 0.910 3.850 2.794 ;
        RECT 3.850 0.900 3.860 2.794 ;
        RECT 3.860 0.890 3.870 2.794 ;
        RECT 3.870 0.880 3.880 2.794 ;
        RECT 2.640 2.890 2.810 3.190 ;
        RECT 3.425 3.020 4.285 3.100 ;
        RECT 3.435 3.020 4.285 3.110 ;
        RECT 3.445 3.020 4.285 3.120 ;
        RECT 3.455 3.020 4.285 3.130 ;
        RECT 3.465 3.020 4.285 3.140 ;
        RECT 3.475 3.020 4.285 3.150 ;
        RECT 3.485 3.020 4.285 3.160 ;
        RECT 3.495 3.020 4.285 3.170 ;
        RECT 2.640 2.920 3.505 3.090 ;
        RECT 3.505 3.020 4.285 3.180 ;
        RECT 2.640 2.930 3.515 3.090 ;
        RECT 2.640 2.940 3.525 3.090 ;
        RECT 2.640 2.950 3.535 3.090 ;
        RECT 2.640 2.960 3.545 3.090 ;
        RECT 2.640 2.970 3.555 3.090 ;
        RECT 2.640 2.980 3.565 3.090 ;
        RECT 2.640 2.990 3.575 3.090 ;
        RECT 2.640 3.000 3.585 3.090 ;
        RECT 2.640 3.010 3.595 3.090 ;
        RECT 4.115 2.855 4.285 3.190 ;
        RECT 3.515 3.020 4.285 3.190 ;
        RECT 4.115 2.855 5.220 3.025 ;
        RECT 5.050 2.855 5.220 3.155 ;
        RECT 4.135 1.135 4.350 1.435 ;
        RECT 4.115 2.060 4.285 2.390 ;
        RECT 4.180 1.135 4.350 2.225 ;
        RECT 6.240 1.060 6.480 1.360 ;
        RECT 4.180 2.055 6.555 2.225 ;
        RECT 6.285 1.060 6.480 2.225 ;
        RECT 6.385 2.055 6.555 2.640 ;
        RECT 6.385 2.470 7.235 2.640 ;
        RECT 7.065 2.470 7.235 2.770 ;
        RECT 5.890 0.710 6.060 1.845 ;
        RECT 4.710 1.675 6.060 1.845 ;
        RECT 5.890 0.710 7.335 0.880 ;
        RECT 7.165 0.710 7.335 1.295 ;
        RECT 7.165 1.125 8.135 1.295 ;
        RECT 7.965 1.125 8.135 2.280 ;
        RECT 7.965 1.640 8.505 2.280 ;
  END 
END LATSRHDLXHT

MACRO LATSRHD2XHT
  CLASS  CORE ;
  FOREIGN LATSRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.070 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.045 1.125 8.345 1.295 ;
        RECT 8.175 1.125 8.190 2.960 ;
        RECT 8.020 1.980 8.190 2.960 ;
        RECT 8.175 1.125 8.345 2.170 ;
        RECT 8.020 1.980 8.345 2.170 ;
        RECT 8.175 1.740 8.580 1.950 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.145 0.785 10.445 1.335 ;
        RECT 10.145 2.150 10.445 3.000 ;
        RECT 10.145 1.105 10.955 1.335 ;
        RECT 10.785 1.105 10.955 2.360 ;
        RECT 10.145 2.150 10.955 2.360 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.380 1.265 3.590 1.925 ;
        RECT 3.380 1.755 3.795 1.925 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.565 0.965 2.055 ;
    END
  END G
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.620 0.500 2.920 0.700 ;
        RECT 2.620 0.530 5.745 0.700 ;
        RECT 5.325 0.500 5.745 0.720 ;
        RECT 5.315 0.530 5.745 0.720 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 2.270 -0.300 2.440 0.660 ;
        RECT 6.255 -0.300 6.555 0.980 ;
        RECT 7.495 -0.300 7.795 0.595 ;
        RECT 8.595 -0.300 8.895 0.595 ;
        RECT 9.625 -0.300 9.925 0.715 ;
        RECT 10.665 -0.300 10.965 0.715 ;
        RECT 0.000 -0.300 11.070 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.530 2.745 2.035 3.180 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.915 0.895 3.990 ;
        RECT 2.240 2.910 2.440 3.990 ;
        RECT 6.090 2.540 6.395 3.990 ;
        RECT 7.435 2.635 7.735 3.990 ;
        RECT 8.540 2.230 8.710 3.990 ;
        RECT 9.625 2.295 9.925 3.990 ;
        RECT 10.665 2.635 10.965 3.990 ;
        RECT 0.000 3.390 11.070 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 0.275 2.565 ;
        RECT 0.105 1.125 0.405 1.295 ;
        RECT 0.105 2.345 0.405 2.565 ;
        RECT 1.075 2.395 1.245 2.950 ;
        RECT 0.105 2.395 2.790 2.565 ;
        RECT 2.620 2.395 2.790 3.080 ;
        RECT 2.620 2.910 3.795 3.080 ;
        RECT 3.495 2.910 3.795 3.190 ;
        RECT 3.845 1.230 4.145 1.400 ;
        RECT 3.975 1.230 4.145 2.320 ;
        RECT 3.360 2.150 4.145 2.320 ;
        RECT 1.210 0.775 1.380 2.215 ;
        RECT 1.145 2.045 1.445 2.215 ;
        RECT 1.210 0.775 2.035 0.945 ;
        RECT 2.230 0.880 4.325 1.050 ;
        RECT 4.735 2.670 5.085 2.840 ;
        RECT 4.655 2.600 4.665 2.840 ;
        RECT 4.665 2.610 4.675 2.840 ;
        RECT 4.675 2.620 4.685 2.840 ;
        RECT 4.685 2.630 4.695 2.840 ;
        RECT 4.695 2.640 4.705 2.840 ;
        RECT 4.705 2.650 4.715 2.840 ;
        RECT 4.715 2.660 4.725 2.840 ;
        RECT 4.725 2.670 4.735 2.840 ;
        RECT 4.495 2.440 4.505 2.680 ;
        RECT 4.505 2.450 4.515 2.690 ;
        RECT 4.515 2.460 4.525 2.700 ;
        RECT 4.525 2.470 4.535 2.710 ;
        RECT 4.535 2.480 4.545 2.720 ;
        RECT 4.545 2.490 4.555 2.730 ;
        RECT 4.555 2.500 4.565 2.740 ;
        RECT 4.565 2.510 4.575 2.750 ;
        RECT 4.575 2.520 4.585 2.760 ;
        RECT 4.585 2.530 4.595 2.770 ;
        RECT 4.595 2.540 4.605 2.780 ;
        RECT 4.605 2.550 4.615 2.790 ;
        RECT 4.615 2.560 4.625 2.800 ;
        RECT 4.625 2.570 4.635 2.810 ;
        RECT 4.635 2.580 4.645 2.820 ;
        RECT 4.645 2.590 4.655 2.830 ;
        RECT 4.325 0.880 4.335 2.510 ;
        RECT 4.335 0.880 4.345 2.520 ;
        RECT 4.345 0.880 4.355 2.530 ;
        RECT 4.355 0.880 4.365 2.540 ;
        RECT 4.365 0.880 4.375 2.550 ;
        RECT 4.375 0.880 4.385 2.560 ;
        RECT 4.385 0.880 4.395 2.570 ;
        RECT 4.395 0.880 4.405 2.580 ;
        RECT 4.405 0.880 4.415 2.590 ;
        RECT 4.415 0.880 4.425 2.600 ;
        RECT 4.425 0.880 4.435 2.610 ;
        RECT 4.435 0.880 4.445 2.620 ;
        RECT 4.445 0.880 4.455 2.630 ;
        RECT 4.455 0.880 4.465 2.640 ;
        RECT 4.465 0.880 4.475 2.650 ;
        RECT 4.475 0.880 4.485 2.660 ;
        RECT 4.485 0.880 4.495 2.670 ;
        RECT 2.140 0.800 2.150 1.050 ;
        RECT 2.150 0.810 2.160 1.050 ;
        RECT 2.160 0.820 2.170 1.050 ;
        RECT 2.170 0.830 2.180 1.050 ;
        RECT 2.180 0.840 2.190 1.050 ;
        RECT 2.190 0.850 2.200 1.050 ;
        RECT 2.200 0.860 2.210 1.050 ;
        RECT 2.210 0.870 2.220 1.050 ;
        RECT 2.220 0.880 2.230 1.050 ;
        RECT 2.125 0.785 2.135 1.035 ;
        RECT 2.135 0.790 2.141 1.044 ;
        RECT 2.035 0.775 2.045 0.945 ;
        RECT 2.045 0.775 2.055 0.955 ;
        RECT 2.055 0.775 2.065 0.965 ;
        RECT 2.065 0.775 2.075 0.975 ;
        RECT 2.075 0.775 2.085 0.985 ;
        RECT 2.085 0.775 2.095 0.995 ;
        RECT 2.095 0.775 2.105 1.005 ;
        RECT 2.105 0.775 2.115 1.015 ;
        RECT 2.115 0.775 2.125 1.025 ;
        RECT 1.655 1.125 1.955 1.295 ;
        RECT 1.785 1.125 1.955 2.215 ;
        RECT 2.450 1.610 2.620 2.215 ;
        RECT 1.655 2.045 3.140 2.215 ;
        RECT 2.970 2.045 3.140 2.730 ;
        RECT 2.970 2.560 3.945 2.730 ;
        RECT 4.240 2.850 4.325 3.020 ;
        RECT 5.225 2.995 5.395 3.190 ;
        RECT 4.575 3.020 5.395 3.190 ;
        RECT 5.225 2.995 5.565 3.165 ;
        RECT 4.495 2.950 4.505 3.190 ;
        RECT 4.505 2.960 4.515 3.190 ;
        RECT 4.515 2.970 4.525 3.190 ;
        RECT 4.525 2.980 4.535 3.190 ;
        RECT 4.535 2.990 4.545 3.190 ;
        RECT 4.545 3.000 4.555 3.190 ;
        RECT 4.555 3.010 4.565 3.190 ;
        RECT 4.565 3.020 4.575 3.190 ;
        RECT 4.405 2.860 4.415 3.100 ;
        RECT 4.415 2.870 4.425 3.110 ;
        RECT 4.425 2.880 4.435 3.120 ;
        RECT 4.435 2.890 4.445 3.130 ;
        RECT 4.445 2.900 4.455 3.140 ;
        RECT 4.455 2.910 4.465 3.150 ;
        RECT 4.465 2.920 4.475 3.160 ;
        RECT 4.475 2.930 4.485 3.170 ;
        RECT 4.485 2.940 4.495 3.180 ;
        RECT 4.325 2.850 4.335 3.020 ;
        RECT 4.335 2.850 4.345 3.030 ;
        RECT 4.345 2.850 4.355 3.040 ;
        RECT 4.355 2.850 4.365 3.050 ;
        RECT 4.365 2.850 4.375 3.060 ;
        RECT 4.375 2.850 4.385 3.070 ;
        RECT 4.385 2.850 4.395 3.080 ;
        RECT 4.395 2.850 4.405 3.090 ;
        RECT 4.070 2.580 4.080 3.020 ;
        RECT 4.080 2.590 4.090 3.020 ;
        RECT 4.090 2.600 4.100 3.020 ;
        RECT 4.100 2.610 4.110 3.020 ;
        RECT 4.110 2.620 4.120 3.020 ;
        RECT 4.120 2.630 4.130 3.020 ;
        RECT 4.130 2.640 4.140 3.020 ;
        RECT 4.140 2.650 4.150 3.020 ;
        RECT 4.150 2.660 4.160 3.020 ;
        RECT 4.160 2.670 4.170 3.020 ;
        RECT 4.170 2.680 4.180 3.020 ;
        RECT 4.180 2.690 4.190 3.020 ;
        RECT 4.190 2.700 4.200 3.020 ;
        RECT 4.200 2.710 4.210 3.020 ;
        RECT 4.210 2.720 4.220 3.020 ;
        RECT 4.220 2.730 4.230 3.020 ;
        RECT 4.230 2.740 4.240 3.020 ;
        RECT 4.060 2.570 4.070 2.844 ;
        RECT 3.945 2.560 3.955 2.730 ;
        RECT 3.955 2.560 3.965 2.740 ;
        RECT 3.965 2.560 3.975 2.750 ;
        RECT 3.975 2.560 3.985 2.760 ;
        RECT 3.985 2.560 3.995 2.770 ;
        RECT 3.995 2.560 4.005 2.780 ;
        RECT 4.005 2.560 4.015 2.790 ;
        RECT 4.015 2.560 4.025 2.800 ;
        RECT 4.025 2.560 4.035 2.810 ;
        RECT 4.035 2.560 4.045 2.820 ;
        RECT 4.045 2.560 4.055 2.830 ;
        RECT 4.055 2.560 4.061 2.840 ;
        RECT 6.870 1.610 7.040 1.970 ;
        RECT 5.845 1.795 7.040 1.970 ;
        RECT 6.825 0.810 7.495 1.065 ;
        RECT 4.675 0.890 4.845 2.350 ;
        RECT 4.675 0.890 4.975 1.400 ;
        RECT 7.015 2.160 7.525 2.350 ;
        RECT 7.355 1.630 7.525 2.350 ;
        RECT 4.675 2.180 7.525 2.350 ;
        RECT 7.355 1.630 7.995 1.800 ;
        RECT 5.430 1.245 5.600 1.825 ;
        RECT 7.695 0.775 7.865 1.430 ;
        RECT 5.430 1.245 7.865 1.430 ;
        RECT 7.695 0.775 9.380 0.945 ;
        RECT 9.210 0.775 9.380 2.555 ;
        RECT 9.025 2.045 9.380 2.555 ;
        RECT 9.210 1.580 10.605 1.750 ;
  END 
END LATSRHD2XHT

MACRO LATSRHD1XHT
  CLASS  CORE ;
  FOREIGN LATSRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.430 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.205 1.125 7.375 3.145 ;
        RECT 6.970 2.470 7.375 3.145 ;
        RECT 7.105 1.125 7.405 1.295 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.090 0.715 9.330 3.100 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.970 1.185 3.180 1.910 ;
        RECT 2.970 1.610 3.370 1.910 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.565 0.965 2.055 ;
    END
  END G
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.020 0.480 5.230 1.235 ;
        RECT 5.020 0.480 5.705 0.650 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 2.265 -0.300 2.565 0.595 ;
        RECT 5.885 -0.300 6.055 1.085 ;
        RECT 7.770 -0.300 8.070 0.715 ;
        RECT 8.505 -0.300 8.805 0.715 ;
        RECT 0.000 -0.300 9.430 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.580 2.745 2.035 3.180 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.905 0.895 3.990 ;
        RECT 2.270 2.745 2.440 3.990 ;
        RECT 5.630 2.430 5.930 3.990 ;
        RECT 7.555 2.230 7.725 3.990 ;
        RECT 8.505 2.630 8.805 3.990 ;
        RECT 0.000 3.390 9.430 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.655 1.125 1.955 1.295 ;
        RECT 1.785 1.125 1.955 2.215 ;
        RECT 1.655 2.045 1.955 2.215 ;
        RECT 1.785 1.675 2.550 1.845 ;
        RECT 2.380 1.610 2.550 1.910 ;
        RECT 3.420 1.060 3.720 1.360 ;
        RECT 3.550 1.060 3.720 2.290 ;
        RECT 3.315 2.120 3.720 2.290 ;
        RECT 1.210 0.775 1.380 2.215 ;
        RECT 1.145 2.045 1.445 2.215 ;
        RECT 2.975 0.605 3.145 0.945 ;
        RECT 1.210 0.775 3.145 0.945 ;
        RECT 2.975 0.605 3.960 0.775 ;
        RECT 0.105 1.125 0.275 2.565 ;
        RECT 0.105 1.125 0.405 1.295 ;
        RECT 0.105 2.345 0.405 2.565 ;
        RECT 1.075 2.395 1.245 2.950 ;
        RECT 2.665 2.395 2.890 2.710 ;
        RECT 0.105 2.395 2.890 2.565 ;
        RECT 2.665 2.505 3.900 2.710 ;
        RECT 3.760 2.505 3.900 2.860 ;
        RECT 4.540 0.605 4.840 1.020 ;
        RECT 4.265 0.820 4.840 1.020 ;
        RECT 4.180 0.820 4.190 1.094 ;
        RECT 4.190 0.820 4.200 1.084 ;
        RECT 4.200 0.820 4.210 1.074 ;
        RECT 4.210 0.820 4.220 1.064 ;
        RECT 4.220 0.820 4.230 1.054 ;
        RECT 4.230 0.820 4.240 1.044 ;
        RECT 4.240 0.820 4.250 1.034 ;
        RECT 4.250 0.820 4.260 1.024 ;
        RECT 4.260 0.820 4.266 1.020 ;
        RECT 4.070 0.930 4.080 1.204 ;
        RECT 4.080 0.920 4.090 1.194 ;
        RECT 4.090 0.910 4.100 1.184 ;
        RECT 4.100 0.900 4.110 1.174 ;
        RECT 4.110 0.890 4.120 1.164 ;
        RECT 4.120 0.880 4.130 1.154 ;
        RECT 4.130 0.870 4.140 1.144 ;
        RECT 4.140 0.860 4.150 1.134 ;
        RECT 4.150 0.850 4.160 1.124 ;
        RECT 4.160 0.840 4.170 1.114 ;
        RECT 4.170 0.830 4.180 1.104 ;
        RECT 3.900 1.100 3.910 2.860 ;
        RECT 3.910 1.090 3.920 2.860 ;
        RECT 3.920 1.080 3.930 2.860 ;
        RECT 3.930 1.070 3.940 2.860 ;
        RECT 3.940 1.060 3.950 2.860 ;
        RECT 3.950 1.050 3.960 2.860 ;
        RECT 3.960 1.040 3.970 2.860 ;
        RECT 3.970 1.030 3.980 2.860 ;
        RECT 3.980 1.020 3.990 2.860 ;
        RECT 3.990 1.010 4.000 2.860 ;
        RECT 4.000 1.000 4.010 2.860 ;
        RECT 4.010 0.990 4.020 2.860 ;
        RECT 4.020 0.980 4.030 2.860 ;
        RECT 4.030 0.970 4.040 2.860 ;
        RECT 4.040 0.960 4.050 2.860 ;
        RECT 4.050 0.950 4.060 2.860 ;
        RECT 4.060 0.940 4.070 2.860 ;
        RECT 2.640 2.910 2.810 3.210 ;
        RECT 2.640 2.910 3.470 3.080 ;
        RECT 4.250 2.910 4.420 3.210 ;
        RECT 3.680 3.040 4.420 3.210 ;
        RECT 4.250 2.910 5.130 3.080 ;
        RECT 4.830 2.910 5.130 3.210 ;
        RECT 3.600 2.970 3.610 3.210 ;
        RECT 3.610 2.980 3.620 3.210 ;
        RECT 3.620 2.990 3.630 3.210 ;
        RECT 3.630 3.000 3.640 3.210 ;
        RECT 3.640 3.010 3.650 3.210 ;
        RECT 3.650 3.020 3.660 3.210 ;
        RECT 3.660 3.030 3.670 3.210 ;
        RECT 3.670 3.040 3.680 3.210 ;
        RECT 3.550 2.920 3.560 3.160 ;
        RECT 3.560 2.930 3.570 3.170 ;
        RECT 3.570 2.940 3.580 3.180 ;
        RECT 3.580 2.950 3.590 3.190 ;
        RECT 3.590 2.960 3.600 3.200 ;
        RECT 3.470 2.910 3.480 3.080 ;
        RECT 3.480 2.910 3.490 3.090 ;
        RECT 3.490 2.910 3.500 3.100 ;
        RECT 3.500 2.910 3.510 3.110 ;
        RECT 3.510 2.910 3.520 3.120 ;
        RECT 3.520 2.910 3.530 3.130 ;
        RECT 3.530 2.910 3.540 3.140 ;
        RECT 3.540 2.910 3.550 3.150 ;
        RECT 6.405 0.480 6.575 1.085 ;
        RECT 6.405 0.480 6.810 0.650 ;
        RECT 4.345 1.200 4.515 2.435 ;
        RECT 4.345 1.200 4.645 1.370 ;
        RECT 6.690 1.630 6.860 2.240 ;
        RECT 4.345 2.070 6.860 2.240 ;
        RECT 6.690 1.630 7.025 1.800 ;
        RECT 6.180 1.265 6.350 1.845 ;
        RECT 4.970 1.675 6.350 1.845 ;
        RECT 6.180 1.265 6.755 1.450 ;
        RECT 7.025 0.775 7.485 0.945 ;
        RECT 7.755 0.960 8.320 1.130 ;
        RECT 8.150 0.960 8.320 2.280 ;
        RECT 8.110 1.980 8.320 2.280 ;
        RECT 8.150 1.515 8.910 1.815 ;
        RECT 7.670 0.885 7.680 1.129 ;
        RECT 7.680 0.895 7.690 1.129 ;
        RECT 7.690 0.905 7.700 1.129 ;
        RECT 7.700 0.915 7.710 1.129 ;
        RECT 7.710 0.925 7.720 1.129 ;
        RECT 7.720 0.935 7.730 1.129 ;
        RECT 7.730 0.945 7.740 1.129 ;
        RECT 7.740 0.955 7.750 1.129 ;
        RECT 7.750 0.960 7.756 1.130 ;
        RECT 7.570 0.785 7.580 1.029 ;
        RECT 7.580 0.795 7.590 1.039 ;
        RECT 7.590 0.805 7.600 1.049 ;
        RECT 7.600 0.815 7.610 1.059 ;
        RECT 7.610 0.825 7.620 1.069 ;
        RECT 7.620 0.835 7.630 1.079 ;
        RECT 7.630 0.845 7.640 1.089 ;
        RECT 7.640 0.855 7.650 1.099 ;
        RECT 7.650 0.865 7.660 1.109 ;
        RECT 7.660 0.875 7.670 1.119 ;
        RECT 7.485 0.775 7.495 0.945 ;
        RECT 7.495 0.775 7.505 0.955 ;
        RECT 7.505 0.775 7.515 0.965 ;
        RECT 7.515 0.775 7.525 0.975 ;
        RECT 7.525 0.775 7.535 0.985 ;
        RECT 7.535 0.775 7.545 0.995 ;
        RECT 7.545 0.775 7.555 1.005 ;
        RECT 7.555 0.775 7.565 1.015 ;
        RECT 7.565 0.775 7.571 1.025 ;
        RECT 6.945 0.775 6.955 1.015 ;
        RECT 6.955 0.775 6.965 1.005 ;
        RECT 6.965 0.775 6.975 0.995 ;
        RECT 6.975 0.775 6.985 0.985 ;
        RECT 6.985 0.775 6.995 0.975 ;
        RECT 6.995 0.775 7.005 0.965 ;
        RECT 7.005 0.775 7.015 0.955 ;
        RECT 7.015 0.775 7.025 0.945 ;
        RECT 6.925 0.795 6.935 1.035 ;
        RECT 6.935 0.785 6.945 1.025 ;
        RECT 6.755 0.965 6.765 1.449 ;
        RECT 6.765 0.955 6.775 1.449 ;
        RECT 6.775 0.945 6.785 1.449 ;
        RECT 6.785 0.935 6.795 1.449 ;
        RECT 6.795 0.925 6.805 1.449 ;
        RECT 6.805 0.915 6.815 1.449 ;
        RECT 6.815 0.905 6.825 1.449 ;
        RECT 6.825 0.895 6.835 1.449 ;
        RECT 6.835 0.885 6.845 1.449 ;
        RECT 6.845 0.875 6.855 1.449 ;
        RECT 6.855 0.865 6.865 1.449 ;
        RECT 6.865 0.855 6.875 1.449 ;
        RECT 6.875 0.845 6.885 1.449 ;
        RECT 6.885 0.835 6.895 1.449 ;
        RECT 6.895 0.825 6.905 1.449 ;
        RECT 6.905 0.815 6.915 1.449 ;
        RECT 6.915 0.805 6.925 1.449 ;
  END 
END LATSRHD1XHT

MACRO LATSHDMXHT
  CLASS  CORE ;
  FOREIGN LATSHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.790 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 6.410 1.060 6.580 2.280 ;
        RECT 6.410 1.660 6.895 2.025 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.450 1.060 7.645 2.280 ;
        RECT 7.450 1.630 7.690 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.340 2.480 4.640 3.210 ;
        RECT 4.340 2.480 4.825 2.840 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.520 3.000 ;
    END
  END G
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.540 -0.300 0.840 0.745 ;
        RECT 2.255 -0.300 2.425 1.060 ;
        RECT 4.415 -0.300 4.715 0.595 ;
        RECT 5.375 -0.300 5.675 0.720 ;
        RECT 6.865 -0.300 7.165 1.145 ;
        RECT 0.000 -0.300 7.790 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.620 0.510 2.045 0.895 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.730 2.840 0.900 3.990 ;
        RECT 2.060 3.095 2.360 3.990 ;
        RECT 5.190 2.405 5.490 3.990 ;
        RECT 6.835 2.925 7.135 3.990 ;
        RECT 0.000 3.390 7.790 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 3.045 1.060 3.215 2.215 ;
        RECT 2.980 2.045 3.280 2.215 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.520 0.835 1.755 ;
        RECT 1.250 2.745 3.630 2.915 ;
        RECT 1.080 2.450 1.090 2.914 ;
        RECT 1.090 2.460 1.100 2.914 ;
        RECT 1.100 2.470 1.110 2.914 ;
        RECT 1.110 2.480 1.120 2.914 ;
        RECT 1.120 2.490 1.130 2.914 ;
        RECT 1.130 2.500 1.140 2.914 ;
        RECT 1.140 2.510 1.150 2.914 ;
        RECT 1.150 2.520 1.160 2.914 ;
        RECT 1.160 2.530 1.170 2.914 ;
        RECT 1.170 2.540 1.180 2.914 ;
        RECT 1.180 2.550 1.190 2.914 ;
        RECT 1.190 2.560 1.200 2.914 ;
        RECT 1.200 2.570 1.210 2.914 ;
        RECT 1.210 2.580 1.220 2.914 ;
        RECT 1.220 2.590 1.230 2.914 ;
        RECT 1.230 2.600 1.240 2.914 ;
        RECT 1.240 2.610 1.250 2.914 ;
        RECT 1.005 2.375 1.015 2.625 ;
        RECT 1.015 2.385 1.025 2.635 ;
        RECT 1.025 2.395 1.035 2.645 ;
        RECT 1.035 2.405 1.045 2.655 ;
        RECT 1.045 2.415 1.055 2.665 ;
        RECT 1.055 2.425 1.065 2.675 ;
        RECT 1.065 2.435 1.075 2.685 ;
        RECT 1.075 2.440 1.081 2.694 ;
        RECT 0.835 1.520 0.845 2.454 ;
        RECT 0.845 1.520 0.855 2.464 ;
        RECT 0.855 1.520 0.865 2.474 ;
        RECT 0.865 1.520 0.875 2.484 ;
        RECT 0.875 1.520 0.885 2.494 ;
        RECT 0.885 1.520 0.895 2.504 ;
        RECT 0.895 1.520 0.905 2.514 ;
        RECT 0.905 1.520 0.915 2.524 ;
        RECT 0.915 1.520 0.925 2.534 ;
        RECT 0.925 1.520 0.935 2.544 ;
        RECT 0.935 1.520 0.945 2.554 ;
        RECT 0.945 1.520 0.955 2.564 ;
        RECT 0.955 1.520 0.965 2.574 ;
        RECT 0.965 1.520 0.975 2.584 ;
        RECT 0.975 1.520 0.985 2.594 ;
        RECT 0.985 1.520 0.995 2.604 ;
        RECT 0.995 1.520 1.005 2.614 ;
        RECT 1.550 2.395 4.095 2.565 ;
        RECT 3.925 2.395 4.095 2.950 ;
        RECT 1.465 2.320 1.475 2.564 ;
        RECT 1.475 2.330 1.485 2.564 ;
        RECT 1.485 2.340 1.495 2.564 ;
        RECT 1.495 2.350 1.505 2.564 ;
        RECT 1.505 2.360 1.515 2.564 ;
        RECT 1.515 2.370 1.525 2.564 ;
        RECT 1.525 2.380 1.535 2.564 ;
        RECT 1.535 2.390 1.545 2.564 ;
        RECT 1.545 2.395 1.551 2.565 ;
        RECT 1.360 2.215 1.370 2.459 ;
        RECT 1.370 2.225 1.380 2.469 ;
        RECT 1.380 2.235 1.390 2.479 ;
        RECT 1.390 2.245 1.400 2.489 ;
        RECT 1.400 2.255 1.410 2.499 ;
        RECT 1.410 2.265 1.420 2.509 ;
        RECT 1.420 2.275 1.430 2.519 ;
        RECT 1.430 2.285 1.440 2.529 ;
        RECT 1.440 2.295 1.450 2.539 ;
        RECT 1.450 2.305 1.460 2.549 ;
        RECT 1.460 2.310 1.466 2.560 ;
        RECT 1.185 1.060 1.195 2.284 ;
        RECT 1.195 1.060 1.205 2.294 ;
        RECT 1.205 1.060 1.215 2.304 ;
        RECT 1.215 1.060 1.225 2.314 ;
        RECT 1.225 1.060 1.235 2.324 ;
        RECT 1.235 1.060 1.245 2.334 ;
        RECT 1.245 1.060 1.255 2.344 ;
        RECT 1.255 1.060 1.265 2.354 ;
        RECT 1.265 1.060 1.275 2.364 ;
        RECT 1.275 1.060 1.285 2.374 ;
        RECT 1.285 1.060 1.295 2.384 ;
        RECT 1.295 1.060 1.305 2.394 ;
        RECT 1.305 1.060 1.315 2.404 ;
        RECT 1.315 1.060 1.325 2.414 ;
        RECT 1.325 1.060 1.335 2.424 ;
        RECT 1.335 1.060 1.345 2.434 ;
        RECT 1.345 1.060 1.355 2.444 ;
        RECT 1.355 1.060 1.361 2.454 ;
        RECT 1.630 1.125 1.930 1.295 ;
        RECT 1.760 1.125 1.930 2.215 ;
        RECT 1.630 2.045 1.930 2.215 ;
        RECT 2.615 0.620 2.785 1.845 ;
        RECT 1.760 1.675 2.785 1.845 ;
        RECT 3.745 0.620 3.945 0.945 ;
        RECT 2.615 0.620 3.945 0.790 ;
        RECT 4.905 0.500 5.075 0.945 ;
        RECT 3.745 0.775 5.075 0.945 ;
        RECT 3.540 1.125 3.710 2.215 ;
        RECT 3.540 2.045 3.905 2.215 ;
        RECT 3.540 1.125 5.840 1.295 ;
        RECT 5.960 0.485 6.195 0.785 ;
        RECT 4.325 1.495 6.195 1.665 ;
        RECT 5.830 2.045 6.195 2.215 ;
        RECT 6.025 0.485 6.195 2.630 ;
        RECT 7.100 1.520 7.270 2.630 ;
        RECT 6.025 2.460 7.270 2.630 ;
  END 
END LATSHDMXHT

MACRO LATSHDLXHT
  CLASS  CORE ;
  FOREIGN LATSHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.790 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 6.410 1.060 6.580 2.280 ;
        RECT 6.410 1.660 6.895 2.025 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.450 1.060 7.620 2.430 ;
        RECT 7.450 2.045 7.690 2.430 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.315 2.480 4.615 3.095 ;
        RECT 4.315 2.480 4.820 2.840 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.520 3.000 ;
    END
  END G
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.825 ;
        RECT 2.385 -0.300 2.555 1.160 ;
        RECT 4.400 -0.300 4.700 0.595 ;
        RECT 5.375 -0.300 5.675 0.805 ;
        RECT 6.865 -0.300 7.165 1.295 ;
        RECT 0.000 -0.300 7.790 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.645 0.510 2.070 0.940 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.755 2.785 0.925 3.990 ;
        RECT 2.085 3.095 2.385 3.990 ;
        RECT 5.255 2.315 5.555 3.990 ;
        RECT 6.835 2.810 7.135 3.990 ;
        RECT 0.000 3.390 7.790 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 3.085 1.060 3.255 2.215 ;
        RECT 3.070 2.045 3.370 2.215 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.520 0.860 1.690 ;
        RECT 2.685 2.745 2.855 2.985 ;
        RECT 1.275 2.745 2.855 2.915 ;
        RECT 2.685 2.815 3.650 2.985 ;
        RECT 1.105 2.455 1.115 2.915 ;
        RECT 1.115 2.465 1.125 2.915 ;
        RECT 1.125 2.475 1.135 2.915 ;
        RECT 1.135 2.485 1.145 2.915 ;
        RECT 1.145 2.495 1.155 2.915 ;
        RECT 1.155 2.505 1.165 2.915 ;
        RECT 1.165 2.515 1.175 2.915 ;
        RECT 1.175 2.525 1.185 2.915 ;
        RECT 1.185 2.535 1.195 2.915 ;
        RECT 1.195 2.545 1.205 2.915 ;
        RECT 1.205 2.555 1.215 2.915 ;
        RECT 1.215 2.565 1.225 2.915 ;
        RECT 1.225 2.575 1.235 2.915 ;
        RECT 1.235 2.585 1.245 2.915 ;
        RECT 1.245 2.595 1.255 2.915 ;
        RECT 1.255 2.605 1.265 2.915 ;
        RECT 1.265 2.615 1.275 2.915 ;
        RECT 1.030 2.380 1.040 2.634 ;
        RECT 1.040 2.390 1.050 2.644 ;
        RECT 1.050 2.400 1.060 2.654 ;
        RECT 1.060 2.410 1.070 2.664 ;
        RECT 1.070 2.420 1.080 2.674 ;
        RECT 1.080 2.430 1.090 2.684 ;
        RECT 1.090 2.440 1.100 2.694 ;
        RECT 1.100 2.445 1.106 2.705 ;
        RECT 0.860 1.520 0.870 2.464 ;
        RECT 0.870 1.520 0.880 2.474 ;
        RECT 0.880 1.520 0.890 2.484 ;
        RECT 0.890 1.520 0.900 2.494 ;
        RECT 0.900 1.520 0.910 2.504 ;
        RECT 0.910 1.520 0.920 2.514 ;
        RECT 0.920 1.520 0.930 2.524 ;
        RECT 0.930 1.520 0.940 2.534 ;
        RECT 0.940 1.520 0.950 2.544 ;
        RECT 0.950 1.520 0.960 2.554 ;
        RECT 0.960 1.520 0.970 2.564 ;
        RECT 0.970 1.520 0.980 2.574 ;
        RECT 0.980 1.520 0.990 2.584 ;
        RECT 0.990 1.520 1.000 2.594 ;
        RECT 1.000 1.520 1.010 2.604 ;
        RECT 1.010 1.520 1.020 2.614 ;
        RECT 1.020 1.520 1.030 2.624 ;
        RECT 3.175 2.395 3.345 2.635 ;
        RECT 1.570 2.395 3.345 2.565 ;
        RECT 3.175 2.465 4.065 2.635 ;
        RECT 3.895 2.465 4.065 2.790 ;
        RECT 1.495 2.330 1.505 2.564 ;
        RECT 1.505 2.340 1.515 2.564 ;
        RECT 1.515 2.350 1.525 2.564 ;
        RECT 1.525 2.360 1.535 2.564 ;
        RECT 1.535 2.370 1.545 2.564 ;
        RECT 1.545 2.380 1.555 2.564 ;
        RECT 1.555 2.390 1.565 2.564 ;
        RECT 1.565 2.395 1.571 2.565 ;
        RECT 1.385 2.220 1.395 2.454 ;
        RECT 1.395 2.230 1.405 2.464 ;
        RECT 1.405 2.240 1.415 2.474 ;
        RECT 1.415 2.250 1.425 2.484 ;
        RECT 1.425 2.260 1.435 2.494 ;
        RECT 1.435 2.270 1.445 2.504 ;
        RECT 1.445 2.280 1.455 2.514 ;
        RECT 1.455 2.290 1.465 2.524 ;
        RECT 1.465 2.300 1.475 2.534 ;
        RECT 1.475 2.310 1.485 2.544 ;
        RECT 1.485 2.320 1.495 2.554 ;
        RECT 1.210 1.050 1.220 2.280 ;
        RECT 1.220 1.050 1.230 2.290 ;
        RECT 1.230 1.050 1.240 2.300 ;
        RECT 1.240 1.050 1.250 2.310 ;
        RECT 1.250 1.050 1.260 2.320 ;
        RECT 1.260 1.050 1.270 2.330 ;
        RECT 1.270 1.050 1.280 2.340 ;
        RECT 1.280 1.050 1.290 2.350 ;
        RECT 1.290 1.050 1.300 2.360 ;
        RECT 1.300 1.050 1.310 2.370 ;
        RECT 1.310 1.050 1.320 2.380 ;
        RECT 1.320 1.050 1.330 2.390 ;
        RECT 1.330 1.050 1.340 2.400 ;
        RECT 1.340 1.050 1.350 2.410 ;
        RECT 1.350 1.050 1.360 2.420 ;
        RECT 1.360 1.050 1.370 2.430 ;
        RECT 1.370 1.050 1.380 2.440 ;
        RECT 1.380 1.050 1.386 2.450 ;
        RECT 1.655 1.125 1.955 1.295 ;
        RECT 1.785 1.125 1.955 2.215 ;
        RECT 1.655 2.045 1.955 2.215 ;
        RECT 2.735 0.710 2.905 1.835 ;
        RECT 1.785 1.665 2.905 1.835 ;
        RECT 3.695 0.710 3.930 0.945 ;
        RECT 2.735 0.710 3.930 0.880 ;
        RECT 4.905 0.500 5.075 0.945 ;
        RECT 3.695 0.775 5.075 0.945 ;
        RECT 3.605 1.125 3.775 2.280 ;
        RECT 3.605 1.980 3.825 2.280 ;
        RECT 3.540 1.125 5.840 1.295 ;
        RECT 5.960 0.570 6.190 0.870 ;
        RECT 4.265 1.585 6.190 1.755 ;
        RECT 5.830 2.045 6.190 2.215 ;
        RECT 6.020 0.570 6.190 2.630 ;
        RECT 7.100 1.520 7.270 2.630 ;
        RECT 6.020 2.460 7.270 2.630 ;
  END 
END LATSHDLXHT

MACRO LATSHD2XHT
  CLASS  CORE ;
  FOREIGN LATSHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.020 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.010 0.720 7.180 2.280 ;
        RECT 7.010 1.670 7.280 2.020 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.050 0.720 8.220 2.960 ;
        RECT 8.050 1.260 8.510 1.610 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.815 1.610 3.180 2.020 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.520 3.040 ;
    END
  END G
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.745 ;
        RECT 2.315 -0.300 2.485 1.020 ;
        RECT 4.575 -0.300 4.875 0.595 ;
        RECT 6.420 -0.300 6.720 0.715 ;
        RECT 7.465 -0.300 7.765 1.120 ;
        RECT 8.505 -0.300 8.805 1.055 ;
        RECT 0.000 -0.300 9.020 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.645 0.510 2.070 0.895 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.775 3.095 1.075 3.990 ;
        RECT 2.025 3.095 2.325 3.990 ;
        RECT 5.025 2.295 5.665 3.990 ;
        RECT 6.425 2.975 6.725 3.990 ;
        RECT 7.465 2.975 7.765 3.990 ;
        RECT 8.505 2.295 8.805 3.990 ;
        RECT 0.000 3.390 9.020 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 3.015 1.125 3.240 1.295 ;
        RECT 2.975 2.205 3.360 2.375 ;
        RECT 3.360 1.180 3.370 2.374 ;
        RECT 3.370 1.190 3.380 2.374 ;
        RECT 3.380 1.200 3.390 2.374 ;
        RECT 3.390 1.210 3.400 2.374 ;
        RECT 3.400 1.220 3.410 2.374 ;
        RECT 3.410 1.230 3.420 2.374 ;
        RECT 3.420 1.240 3.430 2.374 ;
        RECT 3.430 1.250 3.440 2.374 ;
        RECT 3.440 1.260 3.450 2.374 ;
        RECT 3.450 1.270 3.460 2.374 ;
        RECT 3.460 1.280 3.470 2.374 ;
        RECT 3.470 1.290 3.480 2.374 ;
        RECT 3.480 1.300 3.490 2.374 ;
        RECT 3.490 1.310 3.500 2.374 ;
        RECT 3.500 1.320 3.510 2.374 ;
        RECT 3.510 1.330 3.520 2.374 ;
        RECT 3.520 1.340 3.530 2.374 ;
        RECT 3.315 1.135 3.325 1.369 ;
        RECT 3.325 1.145 3.335 1.379 ;
        RECT 3.335 1.155 3.345 1.389 ;
        RECT 3.345 1.165 3.355 1.399 ;
        RECT 3.355 1.170 3.361 1.410 ;
        RECT 3.240 1.125 3.250 1.295 ;
        RECT 3.250 1.125 3.260 1.305 ;
        RECT 3.260 1.125 3.270 1.315 ;
        RECT 3.270 1.125 3.280 1.325 ;
        RECT 3.280 1.125 3.290 1.335 ;
        RECT 3.290 1.125 3.300 1.345 ;
        RECT 3.300 1.125 3.310 1.355 ;
        RECT 3.310 1.125 3.316 1.365 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.520 1.030 1.755 ;
        RECT 0.785 1.520 0.955 2.915 ;
        RECT 0.785 1.520 1.030 1.820 ;
        RECT 0.785 2.745 2.420 2.915 ;
        RECT 2.700 2.950 3.555 3.120 ;
        RECT 2.625 2.885 2.635 3.119 ;
        RECT 2.635 2.895 2.645 3.119 ;
        RECT 2.645 2.905 2.655 3.119 ;
        RECT 2.655 2.915 2.665 3.119 ;
        RECT 2.665 2.925 2.675 3.119 ;
        RECT 2.675 2.935 2.685 3.119 ;
        RECT 2.685 2.945 2.695 3.119 ;
        RECT 2.695 2.950 2.701 3.120 ;
        RECT 2.495 2.755 2.505 2.989 ;
        RECT 2.505 2.765 2.515 2.999 ;
        RECT 2.515 2.775 2.525 3.009 ;
        RECT 2.525 2.785 2.535 3.019 ;
        RECT 2.535 2.795 2.545 3.029 ;
        RECT 2.545 2.805 2.555 3.039 ;
        RECT 2.555 2.815 2.565 3.049 ;
        RECT 2.565 2.825 2.575 3.059 ;
        RECT 2.575 2.835 2.585 3.069 ;
        RECT 2.585 2.845 2.595 3.079 ;
        RECT 2.595 2.855 2.605 3.089 ;
        RECT 2.605 2.865 2.615 3.099 ;
        RECT 2.615 2.875 2.625 3.109 ;
        RECT 2.420 2.745 2.430 2.915 ;
        RECT 2.430 2.745 2.440 2.925 ;
        RECT 2.440 2.745 2.450 2.935 ;
        RECT 2.450 2.745 2.460 2.945 ;
        RECT 2.460 2.745 2.470 2.955 ;
        RECT 2.470 2.745 2.480 2.965 ;
        RECT 2.480 2.745 2.490 2.975 ;
        RECT 2.490 2.745 2.496 2.985 ;
        RECT 1.210 0.480 1.385 2.280 ;
        RECT 1.150 1.980 1.385 2.280 ;
        RECT 1.215 0.480 1.385 2.565 ;
        RECT 1.210 0.480 1.435 0.780 ;
        RECT 1.215 2.395 2.585 2.565 ;
        RECT 2.865 2.600 4.155 2.770 ;
        RECT 3.855 2.600 4.155 2.855 ;
        RECT 2.790 2.535 2.800 2.769 ;
        RECT 2.800 2.545 2.810 2.769 ;
        RECT 2.810 2.555 2.820 2.769 ;
        RECT 2.820 2.565 2.830 2.769 ;
        RECT 2.830 2.575 2.840 2.769 ;
        RECT 2.840 2.585 2.850 2.769 ;
        RECT 2.850 2.595 2.860 2.769 ;
        RECT 2.860 2.600 2.866 2.770 ;
        RECT 2.660 2.405 2.670 2.639 ;
        RECT 2.670 2.415 2.680 2.649 ;
        RECT 2.680 2.425 2.690 2.659 ;
        RECT 2.690 2.435 2.700 2.669 ;
        RECT 2.700 2.445 2.710 2.679 ;
        RECT 2.710 2.455 2.720 2.689 ;
        RECT 2.720 2.465 2.730 2.699 ;
        RECT 2.730 2.475 2.740 2.709 ;
        RECT 2.740 2.485 2.750 2.719 ;
        RECT 2.750 2.495 2.760 2.729 ;
        RECT 2.760 2.505 2.770 2.739 ;
        RECT 2.770 2.515 2.780 2.749 ;
        RECT 2.780 2.525 2.790 2.759 ;
        RECT 2.585 2.395 2.595 2.565 ;
        RECT 2.595 2.395 2.605 2.575 ;
        RECT 2.605 2.395 2.615 2.585 ;
        RECT 2.615 2.395 2.625 2.595 ;
        RECT 2.625 2.395 2.635 2.605 ;
        RECT 2.635 2.395 2.645 2.615 ;
        RECT 2.645 2.395 2.655 2.625 ;
        RECT 2.655 2.395 2.661 2.635 ;
        RECT 1.655 1.125 1.955 1.295 ;
        RECT 1.785 1.125 1.955 2.215 ;
        RECT 1.595 2.045 1.955 2.215 ;
        RECT 2.445 1.240 2.615 1.845 ;
        RECT 1.785 1.675 2.615 1.845 ;
        RECT 2.665 0.545 2.835 1.410 ;
        RECT 2.445 1.240 2.835 1.410 ;
        RECT 2.665 0.545 4.360 0.715 ;
        RECT 4.175 0.545 4.360 0.945 ;
        RECT 5.565 0.585 5.735 0.945 ;
        RECT 4.175 0.775 5.735 0.945 ;
        RECT 3.540 0.900 3.910 1.070 ;
        RECT 3.740 0.900 3.910 2.280 ;
        RECT 3.740 1.125 5.515 1.295 ;
        RECT 5.345 1.125 5.515 1.710 ;
        RECT 5.345 1.540 6.375 1.710 ;
        RECT 4.430 1.550 4.600 2.095 ;
        RECT 5.980 1.925 6.150 2.630 ;
        RECT 5.870 1.125 6.785 1.295 ;
        RECT 6.615 1.125 6.785 2.095 ;
        RECT 4.430 1.925 6.785 2.095 ;
        RECT 7.670 1.520 7.840 2.630 ;
        RECT 5.980 2.460 7.840 2.630 ;
  END 
END LATSHD2XHT

MACRO LATSHD1XHT
  CLASS  CORE ;
  FOREIGN LATSHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.790 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 6.410 1.060 6.580 2.280 ;
        RECT 6.410 1.660 6.895 2.025 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.450 0.720 7.645 2.960 ;
        RECT 7.450 2.455 7.690 2.960 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.445 2.480 4.615 3.210 ;
        RECT 4.315 3.040 4.615 3.210 ;
        RECT 4.445 2.480 4.820 2.840 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.545 3.000 ;
    END
  END G
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.745 ;
        RECT 2.385 -0.300 2.555 1.020 ;
        RECT 4.400 -0.300 4.700 0.595 ;
        RECT 5.375 -0.300 5.675 0.795 ;
        RECT 6.865 -0.300 7.165 1.055 ;
        RECT 0.000 -0.300 7.790 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.645 0.510 2.070 0.895 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.775 3.095 1.075 3.990 ;
        RECT 2.085 3.095 2.385 3.990 ;
        RECT 5.190 2.405 5.490 3.990 ;
        RECT 6.865 2.975 7.165 3.990 ;
        RECT 0.000 3.390 7.790 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 3.085 1.060 3.255 2.215 ;
        RECT 3.070 2.045 3.370 2.215 ;
        RECT 0.195 1.060 0.365 2.280 ;
        RECT 0.195 1.585 1.030 1.755 ;
        RECT 0.860 1.520 1.030 2.915 ;
        RECT 2.710 2.745 2.880 3.035 ;
        RECT 0.860 2.745 2.880 2.915 ;
        RECT 2.710 2.865 3.650 3.035 ;
        RECT 1.210 1.060 1.385 2.565 ;
        RECT 1.210 2.395 4.065 2.565 ;
        RECT 3.895 2.395 4.065 2.920 ;
        RECT 1.655 1.125 1.955 1.295 ;
        RECT 1.785 1.125 1.955 2.215 ;
        RECT 1.655 2.045 1.955 2.215 ;
        RECT 2.735 0.620 2.905 1.665 ;
        RECT 1.785 1.495 2.905 1.665 ;
        RECT 3.765 0.620 3.935 0.945 ;
        RECT 2.735 0.620 3.935 0.790 ;
        RECT 4.905 0.500 5.075 0.945 ;
        RECT 3.765 0.775 5.075 0.945 ;
        RECT 3.540 1.125 3.775 1.360 ;
        RECT 3.590 1.125 3.775 2.215 ;
        RECT 3.590 1.980 3.890 2.215 ;
        RECT 3.540 1.125 5.840 1.295 ;
        RECT 5.960 0.560 6.190 0.860 ;
        RECT 4.265 1.585 6.190 1.755 ;
        RECT 5.830 2.045 6.190 2.215 ;
        RECT 6.020 0.560 6.190 2.630 ;
        RECT 7.100 1.520 7.270 2.630 ;
        RECT 6.020 2.460 7.270 2.630 ;
  END 
END LATSHD1XHT

MACRO LATRHDMXHT
  CLASS  CORE ;
  FOREIGN LATRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.380 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.840 0.840 6.170 1.200 ;
        RECT 6.000 0.840 6.170 2.280 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.040 1.060 7.210 2.280 ;
        RECT 7.040 1.260 7.280 1.610 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.595 2.150 2.135 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.465 0.585 2.885 ;
    END
  END G
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.360 0.645 1.530 0.945 ;
        RECT 2.080 0.545 2.250 0.945 ;
        RECT 1.360 0.775 2.250 0.945 ;
        RECT 4.085 0.500 4.645 0.715 ;
        RECT 2.080 0.545 4.645 0.715 ;
        RECT 4.095 0.500 4.645 0.720 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.745 ;
        RECT 1.730 -0.300 1.900 0.575 ;
        RECT 4.840 -0.300 5.010 1.090 ;
        RECT 4.710 0.920 5.010 1.090 ;
        RECT 6.455 -0.300 6.755 1.145 ;
        RECT 0.000 -0.300 7.380 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.590 3.095 0.890 3.990 ;
        RECT 1.625 3.095 1.925 3.990 ;
        RECT 4.010 2.455 4.310 3.990 ;
        RECT 4.990 2.745 5.290 3.990 ;
        RECT 6.485 2.925 6.785 3.990 ;
        RECT 0.000 3.390 7.380 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.030 1.755 ;
        RECT 0.860 1.520 1.030 2.915 ;
        RECT 0.860 2.745 2.005 2.915 ;
        RECT 2.355 3.020 2.835 3.190 ;
        RECT 2.280 2.955 2.290 3.189 ;
        RECT 2.290 2.965 2.300 3.189 ;
        RECT 2.300 2.975 2.310 3.189 ;
        RECT 2.310 2.985 2.320 3.189 ;
        RECT 2.320 2.995 2.330 3.189 ;
        RECT 2.330 3.005 2.340 3.189 ;
        RECT 2.340 3.015 2.350 3.189 ;
        RECT 2.350 3.020 2.356 3.190 ;
        RECT 2.080 2.755 2.090 2.989 ;
        RECT 2.090 2.765 2.100 2.999 ;
        RECT 2.100 2.775 2.110 3.009 ;
        RECT 2.110 2.785 2.120 3.019 ;
        RECT 2.120 2.795 2.130 3.029 ;
        RECT 2.130 2.805 2.140 3.039 ;
        RECT 2.140 2.815 2.150 3.049 ;
        RECT 2.150 2.825 2.160 3.059 ;
        RECT 2.160 2.835 2.170 3.069 ;
        RECT 2.170 2.845 2.180 3.079 ;
        RECT 2.180 2.855 2.190 3.089 ;
        RECT 2.190 2.865 2.200 3.099 ;
        RECT 2.200 2.875 2.210 3.109 ;
        RECT 2.210 2.885 2.220 3.119 ;
        RECT 2.220 2.895 2.230 3.129 ;
        RECT 2.230 2.905 2.240 3.139 ;
        RECT 2.240 2.915 2.250 3.149 ;
        RECT 2.250 2.925 2.260 3.159 ;
        RECT 2.260 2.935 2.270 3.169 ;
        RECT 2.270 2.945 2.280 3.179 ;
        RECT 2.005 2.745 2.015 2.915 ;
        RECT 2.015 2.745 2.025 2.925 ;
        RECT 2.025 2.745 2.035 2.935 ;
        RECT 2.035 2.745 2.045 2.945 ;
        RECT 2.045 2.745 2.055 2.955 ;
        RECT 2.055 2.745 2.065 2.965 ;
        RECT 2.065 2.745 2.075 2.975 ;
        RECT 2.075 2.745 2.081 2.985 ;
        RECT 2.430 0.895 2.600 2.280 ;
        RECT 2.380 1.980 2.600 2.280 ;
        RECT 2.430 0.895 2.945 1.065 ;
        RECT 1.080 1.125 1.385 1.295 ;
        RECT 1.210 1.125 1.385 2.565 ;
        RECT 1.210 2.395 2.165 2.565 ;
        RECT 2.805 1.290 2.920 2.840 ;
        RECT 2.515 2.670 2.920 2.840 ;
        RECT 2.975 1.290 3.225 1.460 ;
        RECT 3.150 2.825 3.570 2.995 ;
        RECT 3.075 2.760 3.085 2.994 ;
        RECT 3.085 2.770 3.095 2.994 ;
        RECT 3.095 2.780 3.105 2.994 ;
        RECT 3.105 2.790 3.115 2.994 ;
        RECT 3.115 2.800 3.125 2.994 ;
        RECT 3.125 2.810 3.135 2.994 ;
        RECT 3.135 2.820 3.145 2.994 ;
        RECT 3.145 2.825 3.151 2.995 ;
        RECT 2.995 2.680 3.005 2.914 ;
        RECT 3.005 2.690 3.015 2.924 ;
        RECT 3.015 2.700 3.025 2.934 ;
        RECT 3.025 2.710 3.035 2.944 ;
        RECT 3.035 2.720 3.045 2.954 ;
        RECT 3.045 2.730 3.055 2.964 ;
        RECT 3.055 2.740 3.065 2.974 ;
        RECT 3.065 2.750 3.075 2.984 ;
        RECT 2.975 2.670 2.985 2.894 ;
        RECT 2.985 2.670 2.995 2.904 ;
        RECT 2.920 1.290 2.930 2.840 ;
        RECT 2.930 1.290 2.940 2.850 ;
        RECT 2.940 1.290 2.950 2.860 ;
        RECT 2.950 1.290 2.960 2.870 ;
        RECT 2.960 1.290 2.970 2.880 ;
        RECT 2.970 1.290 2.976 2.890 ;
        RECT 2.440 2.605 2.450 2.839 ;
        RECT 2.450 2.615 2.460 2.839 ;
        RECT 2.460 2.625 2.470 2.839 ;
        RECT 2.470 2.635 2.480 2.839 ;
        RECT 2.480 2.645 2.490 2.839 ;
        RECT 2.490 2.655 2.500 2.839 ;
        RECT 2.500 2.665 2.510 2.839 ;
        RECT 2.510 2.670 2.516 2.840 ;
        RECT 2.240 2.405 2.250 2.639 ;
        RECT 2.250 2.415 2.260 2.649 ;
        RECT 2.260 2.425 2.270 2.659 ;
        RECT 2.270 2.435 2.280 2.669 ;
        RECT 2.280 2.445 2.290 2.679 ;
        RECT 2.290 2.455 2.300 2.689 ;
        RECT 2.300 2.465 2.310 2.699 ;
        RECT 2.310 2.475 2.320 2.709 ;
        RECT 2.320 2.485 2.330 2.719 ;
        RECT 2.330 2.495 2.340 2.729 ;
        RECT 2.340 2.505 2.350 2.739 ;
        RECT 2.350 2.515 2.360 2.749 ;
        RECT 2.360 2.525 2.370 2.759 ;
        RECT 2.370 2.535 2.380 2.769 ;
        RECT 2.380 2.545 2.390 2.779 ;
        RECT 2.390 2.555 2.400 2.789 ;
        RECT 2.400 2.565 2.410 2.799 ;
        RECT 2.410 2.575 2.420 2.809 ;
        RECT 2.420 2.585 2.430 2.819 ;
        RECT 2.430 2.595 2.440 2.829 ;
        RECT 2.165 2.395 2.175 2.565 ;
        RECT 2.175 2.395 2.185 2.575 ;
        RECT 2.185 2.395 2.195 2.585 ;
        RECT 2.195 2.395 2.205 2.595 ;
        RECT 2.205 2.395 2.215 2.605 ;
        RECT 2.215 2.395 2.225 2.615 ;
        RECT 2.225 2.395 2.235 2.625 ;
        RECT 2.235 2.395 2.241 2.635 ;
        RECT 3.155 2.040 3.330 2.570 ;
        RECT 3.165 0.895 3.590 1.065 ;
        RECT 3.420 0.895 3.590 2.215 ;
        RECT 4.560 2.040 4.860 2.325 ;
        RECT 3.155 2.040 5.360 2.215 ;
        RECT 5.355 0.855 5.525 1.860 ;
        RECT 3.855 1.690 5.745 1.860 ;
        RECT 5.575 1.690 5.745 2.860 ;
        RECT 6.660 1.540 6.830 2.630 ;
        RECT 5.575 2.460 6.830 2.630 ;
  END 
END LATRHDMXHT

MACRO LATRHDLXHT
  CLASS  CORE ;
  FOREIGN LATRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.380 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.840 0.835 6.170 1.225 ;
        RECT 6.000 0.835 6.170 2.280 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.040 1.060 7.210 2.280 ;
        RECT 7.040 1.060 7.280 1.610 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.735 1.595 2.205 2.135 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.460 0.550 2.840 ;
    END
  END G
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.010 0.550 4.655 0.670 ;
        RECT 2.160 0.500 2.310 0.720 ;
        RECT 2.010 0.500 2.310 0.670 ;
        RECT 4.085 0.500 4.655 0.720 ;
        RECT 2.160 0.550 4.655 0.720 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.825 ;
        RECT 1.660 -0.300 1.830 1.040 ;
        RECT 1.660 0.870 1.995 1.040 ;
        RECT 4.840 -0.300 5.010 1.140 ;
        RECT 4.710 0.970 5.010 1.140 ;
        RECT 6.455 -0.300 6.755 1.295 ;
        RECT 0.000 -0.300 7.380 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.750 2.730 0.920 3.990 ;
        RECT 1.650 3.095 1.950 3.990 ;
        RECT 4.025 2.440 4.325 3.990 ;
        RECT 4.995 2.670 5.295 3.990 ;
        RECT 6.485 2.815 6.785 3.990 ;
        RECT 0.000 3.390 7.380 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 0.885 1.755 ;
        RECT 1.270 2.745 2.035 2.915 ;
        RECT 2.325 2.960 2.790 3.130 ;
        RECT 2.250 2.895 2.260 3.129 ;
        RECT 2.260 2.905 2.270 3.129 ;
        RECT 2.270 2.915 2.280 3.129 ;
        RECT 2.280 2.925 2.290 3.129 ;
        RECT 2.290 2.935 2.300 3.129 ;
        RECT 2.300 2.945 2.310 3.129 ;
        RECT 2.310 2.955 2.320 3.129 ;
        RECT 2.320 2.960 2.326 3.130 ;
        RECT 2.110 2.755 2.120 2.989 ;
        RECT 2.120 2.765 2.130 2.999 ;
        RECT 2.130 2.775 2.140 3.009 ;
        RECT 2.140 2.785 2.150 3.019 ;
        RECT 2.150 2.795 2.160 3.029 ;
        RECT 2.160 2.805 2.170 3.039 ;
        RECT 2.170 2.815 2.180 3.049 ;
        RECT 2.180 2.825 2.190 3.059 ;
        RECT 2.190 2.835 2.200 3.069 ;
        RECT 2.200 2.845 2.210 3.079 ;
        RECT 2.210 2.855 2.220 3.089 ;
        RECT 2.220 2.865 2.230 3.099 ;
        RECT 2.230 2.875 2.240 3.109 ;
        RECT 2.240 2.885 2.250 3.119 ;
        RECT 2.035 2.745 2.045 2.915 ;
        RECT 2.045 2.745 2.055 2.925 ;
        RECT 2.055 2.745 2.065 2.935 ;
        RECT 2.065 2.745 2.075 2.945 ;
        RECT 2.075 2.745 2.085 2.955 ;
        RECT 2.085 2.745 2.095 2.965 ;
        RECT 2.095 2.745 2.105 2.975 ;
        RECT 2.105 2.745 2.111 2.985 ;
        RECT 1.100 2.415 1.110 2.915 ;
        RECT 1.110 2.425 1.120 2.915 ;
        RECT 1.120 2.435 1.130 2.915 ;
        RECT 1.130 2.445 1.140 2.915 ;
        RECT 1.140 2.455 1.150 2.915 ;
        RECT 1.150 2.465 1.160 2.915 ;
        RECT 1.160 2.475 1.170 2.915 ;
        RECT 1.170 2.485 1.180 2.915 ;
        RECT 1.180 2.495 1.190 2.915 ;
        RECT 1.190 2.505 1.200 2.915 ;
        RECT 1.200 2.515 1.210 2.915 ;
        RECT 1.210 2.525 1.220 2.915 ;
        RECT 1.220 2.535 1.230 2.915 ;
        RECT 1.230 2.545 1.240 2.915 ;
        RECT 1.240 2.555 1.250 2.915 ;
        RECT 1.250 2.565 1.260 2.915 ;
        RECT 1.260 2.575 1.270 2.915 ;
        RECT 1.055 2.370 1.065 2.610 ;
        RECT 1.065 2.380 1.075 2.620 ;
        RECT 1.075 2.390 1.085 2.630 ;
        RECT 1.085 2.400 1.095 2.640 ;
        RECT 1.095 2.405 1.101 2.649 ;
        RECT 0.885 1.520 0.895 2.440 ;
        RECT 0.895 1.520 0.905 2.450 ;
        RECT 0.905 1.520 0.915 2.460 ;
        RECT 0.915 1.520 0.925 2.470 ;
        RECT 0.925 1.520 0.935 2.480 ;
        RECT 0.935 1.520 0.945 2.490 ;
        RECT 0.945 1.520 0.955 2.500 ;
        RECT 0.955 1.520 0.965 2.510 ;
        RECT 0.965 1.520 0.975 2.520 ;
        RECT 0.975 1.520 0.985 2.530 ;
        RECT 0.985 1.520 0.995 2.540 ;
        RECT 0.995 1.520 1.005 2.550 ;
        RECT 1.005 1.520 1.015 2.560 ;
        RECT 1.015 1.520 1.025 2.570 ;
        RECT 1.025 1.520 1.035 2.580 ;
        RECT 1.035 1.520 1.045 2.590 ;
        RECT 1.045 1.520 1.055 2.600 ;
        RECT 2.405 0.970 2.575 2.280 ;
        RECT 2.405 0.970 2.970 1.140 ;
        RECT 1.115 1.125 1.235 1.295 ;
        RECT 1.605 2.395 2.190 2.565 ;
        RECT 2.820 1.340 2.885 2.770 ;
        RECT 2.470 2.600 2.885 2.770 ;
        RECT 2.990 1.340 3.260 1.510 ;
        RECT 3.095 2.735 3.585 2.905 ;
        RECT 3.020 2.670 3.030 2.904 ;
        RECT 3.030 2.680 3.040 2.904 ;
        RECT 3.040 2.690 3.050 2.904 ;
        RECT 3.050 2.700 3.060 2.904 ;
        RECT 3.060 2.710 3.070 2.904 ;
        RECT 3.070 2.720 3.080 2.904 ;
        RECT 3.080 2.730 3.090 2.904 ;
        RECT 3.090 2.735 3.096 2.905 ;
        RECT 2.990 2.640 3.000 2.874 ;
        RECT 3.000 2.650 3.010 2.884 ;
        RECT 3.010 2.660 3.020 2.894 ;
        RECT 2.885 1.340 2.895 2.770 ;
        RECT 2.895 1.340 2.905 2.780 ;
        RECT 2.905 1.340 2.915 2.790 ;
        RECT 2.915 1.340 2.925 2.800 ;
        RECT 2.925 1.340 2.935 2.810 ;
        RECT 2.935 1.340 2.945 2.820 ;
        RECT 2.945 1.340 2.955 2.830 ;
        RECT 2.955 1.340 2.965 2.840 ;
        RECT 2.965 1.340 2.975 2.850 ;
        RECT 2.975 1.340 2.985 2.860 ;
        RECT 2.985 1.340 2.991 2.870 ;
        RECT 2.395 2.535 2.405 2.769 ;
        RECT 2.405 2.545 2.415 2.769 ;
        RECT 2.415 2.555 2.425 2.769 ;
        RECT 2.425 2.565 2.435 2.769 ;
        RECT 2.435 2.575 2.445 2.769 ;
        RECT 2.445 2.585 2.455 2.769 ;
        RECT 2.455 2.595 2.465 2.769 ;
        RECT 2.465 2.600 2.471 2.770 ;
        RECT 2.265 2.405 2.275 2.639 ;
        RECT 2.275 2.415 2.285 2.649 ;
        RECT 2.285 2.425 2.295 2.659 ;
        RECT 2.295 2.435 2.305 2.669 ;
        RECT 2.305 2.445 2.315 2.679 ;
        RECT 2.315 2.455 2.325 2.689 ;
        RECT 2.325 2.465 2.335 2.699 ;
        RECT 2.335 2.475 2.345 2.709 ;
        RECT 2.345 2.485 2.355 2.719 ;
        RECT 2.355 2.495 2.365 2.729 ;
        RECT 2.365 2.505 2.375 2.739 ;
        RECT 2.375 2.515 2.385 2.749 ;
        RECT 2.385 2.525 2.395 2.759 ;
        RECT 2.190 2.395 2.200 2.565 ;
        RECT 2.200 2.395 2.210 2.575 ;
        RECT 2.210 2.395 2.220 2.585 ;
        RECT 2.220 2.395 2.230 2.595 ;
        RECT 2.230 2.395 2.240 2.605 ;
        RECT 2.240 2.395 2.250 2.615 ;
        RECT 2.250 2.395 2.260 2.625 ;
        RECT 2.260 2.395 2.266 2.635 ;
        RECT 1.520 2.320 1.530 2.564 ;
        RECT 1.530 2.330 1.540 2.564 ;
        RECT 1.540 2.340 1.550 2.564 ;
        RECT 1.550 2.350 1.560 2.564 ;
        RECT 1.560 2.360 1.570 2.564 ;
        RECT 1.570 2.370 1.580 2.564 ;
        RECT 1.580 2.380 1.590 2.564 ;
        RECT 1.590 2.390 1.600 2.564 ;
        RECT 1.600 2.395 1.606 2.565 ;
        RECT 1.415 2.215 1.425 2.459 ;
        RECT 1.425 2.225 1.435 2.469 ;
        RECT 1.435 2.235 1.445 2.479 ;
        RECT 1.445 2.245 1.455 2.489 ;
        RECT 1.455 2.255 1.465 2.499 ;
        RECT 1.465 2.265 1.475 2.509 ;
        RECT 1.475 2.275 1.485 2.519 ;
        RECT 1.485 2.285 1.495 2.529 ;
        RECT 1.495 2.295 1.505 2.539 ;
        RECT 1.505 2.305 1.515 2.549 ;
        RECT 1.515 2.310 1.521 2.560 ;
        RECT 1.235 1.125 1.245 2.279 ;
        RECT 1.245 1.125 1.255 2.289 ;
        RECT 1.255 1.125 1.265 2.299 ;
        RECT 1.265 1.125 1.275 2.309 ;
        RECT 1.275 1.125 1.285 2.319 ;
        RECT 1.285 1.125 1.295 2.329 ;
        RECT 1.295 1.125 1.305 2.339 ;
        RECT 1.305 1.125 1.315 2.349 ;
        RECT 1.315 1.125 1.325 2.359 ;
        RECT 1.325 1.125 1.335 2.369 ;
        RECT 1.335 1.125 1.345 2.379 ;
        RECT 1.345 1.125 1.355 2.389 ;
        RECT 1.355 1.125 1.365 2.399 ;
        RECT 1.365 1.125 1.375 2.409 ;
        RECT 1.375 1.125 1.385 2.419 ;
        RECT 1.385 1.125 1.395 2.429 ;
        RECT 1.395 1.125 1.405 2.439 ;
        RECT 1.405 1.125 1.415 2.449 ;
        RECT 3.170 2.045 3.340 2.555 ;
        RECT 3.190 0.970 3.655 1.140 ;
        RECT 3.485 0.970 3.655 2.215 ;
        RECT 3.170 2.045 5.380 2.215 ;
        RECT 4.005 1.315 4.175 1.745 ;
        RECT 5.370 0.905 5.540 1.745 ;
        RECT 4.005 1.575 5.750 1.745 ;
        RECT 5.580 1.575 5.750 2.785 ;
        RECT 6.660 1.540 6.830 2.635 ;
        RECT 5.580 2.465 6.830 2.635 ;
  END 
END LATRHDLXHT

MACRO LATRHD2XHT
  CLASS  CORE ;
  FOREIGN LATRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.610 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 6.660 0.845 6.880 1.195 ;
        RECT 6.710 0.720 6.880 2.280 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.750 0.720 7.920 2.960 ;
        RECT 7.750 1.635 8.100 2.035 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.595 2.110 2.120 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.585 2.885 ;
    END
  END G
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.365 0.645 1.540 0.945 ;
        RECT 2.100 0.550 2.270 0.945 ;
        RECT 1.365 0.775 2.270 0.945 ;
        RECT 4.115 0.510 4.610 0.720 ;
        RECT 2.100 0.550 4.610 0.720 ;
        RECT 4.440 0.510 4.610 1.665 ;
        RECT 4.375 1.495 4.675 1.665 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.715 ;
        RECT 1.740 -0.300 1.910 0.575 ;
        RECT 4.840 -0.300 5.140 0.995 ;
        RECT 6.125 -0.300 6.425 1.055 ;
        RECT 7.165 -0.300 7.465 1.055 ;
        RECT 8.200 -0.300 8.505 1.055 ;
        RECT 0.000 -0.300 8.610 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.590 3.095 0.890 3.990 ;
        RECT 1.515 3.095 1.815 3.990 ;
        RECT 4.035 2.975 4.335 3.990 ;
        RECT 5.095 2.585 5.395 3.990 ;
        RECT 6.125 2.975 6.425 3.990 ;
        RECT 7.165 2.975 7.465 3.990 ;
        RECT 8.205 2.295 8.505 3.990 ;
        RECT 0.000 3.390 8.610 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.030 1.755 ;
        RECT 0.860 1.520 1.030 2.915 ;
        RECT 0.860 2.745 1.890 2.915 ;
        RECT 2.265 3.040 2.680 3.210 ;
        RECT 2.185 2.970 2.195 3.210 ;
        RECT 2.195 2.980 2.205 3.210 ;
        RECT 2.205 2.990 2.215 3.210 ;
        RECT 2.215 3.000 2.225 3.210 ;
        RECT 2.225 3.010 2.235 3.210 ;
        RECT 2.235 3.020 2.245 3.210 ;
        RECT 2.245 3.030 2.255 3.210 ;
        RECT 2.255 3.040 2.265 3.210 ;
        RECT 1.970 2.755 1.980 2.995 ;
        RECT 1.980 2.765 1.990 3.005 ;
        RECT 1.990 2.775 2.000 3.015 ;
        RECT 2.000 2.785 2.010 3.025 ;
        RECT 2.010 2.795 2.020 3.035 ;
        RECT 2.020 2.805 2.030 3.045 ;
        RECT 2.030 2.815 2.040 3.055 ;
        RECT 2.040 2.825 2.050 3.065 ;
        RECT 2.050 2.835 2.060 3.075 ;
        RECT 2.060 2.845 2.070 3.085 ;
        RECT 2.070 2.855 2.080 3.095 ;
        RECT 2.080 2.865 2.090 3.105 ;
        RECT 2.090 2.875 2.100 3.115 ;
        RECT 2.100 2.885 2.110 3.125 ;
        RECT 2.110 2.895 2.120 3.135 ;
        RECT 2.120 2.905 2.130 3.145 ;
        RECT 2.130 2.915 2.140 3.155 ;
        RECT 2.140 2.925 2.150 3.165 ;
        RECT 2.150 2.935 2.160 3.175 ;
        RECT 2.160 2.945 2.170 3.185 ;
        RECT 2.170 2.955 2.180 3.195 ;
        RECT 2.180 2.960 2.186 3.204 ;
        RECT 1.890 2.745 1.900 2.915 ;
        RECT 1.900 2.745 1.910 2.925 ;
        RECT 1.910 2.745 1.920 2.935 ;
        RECT 1.920 2.745 1.930 2.945 ;
        RECT 1.930 2.745 1.940 2.955 ;
        RECT 1.940 2.745 1.950 2.965 ;
        RECT 1.950 2.745 1.960 2.975 ;
        RECT 1.960 2.745 1.970 2.985 ;
        RECT 2.450 1.045 2.620 2.450 ;
        RECT 2.445 2.150 2.620 2.450 ;
        RECT 2.450 1.045 2.965 1.215 ;
        RECT 1.070 1.125 1.405 1.295 ;
        RECT 1.210 1.125 1.405 2.565 ;
        RECT 1.210 2.395 2.045 2.565 ;
        RECT 2.800 1.415 2.810 2.860 ;
        RECT 2.415 2.690 2.810 2.860 ;
        RECT 2.970 1.415 3.245 1.585 ;
        RECT 3.175 2.980 3.565 3.150 ;
        RECT 3.100 2.915 3.110 3.149 ;
        RECT 3.110 2.925 3.120 3.149 ;
        RECT 3.120 2.935 3.130 3.149 ;
        RECT 3.130 2.945 3.140 3.149 ;
        RECT 3.140 2.955 3.150 3.149 ;
        RECT 3.150 2.965 3.160 3.149 ;
        RECT 3.160 2.975 3.170 3.149 ;
        RECT 3.170 2.980 3.176 3.150 ;
        RECT 2.970 2.785 2.980 3.019 ;
        RECT 2.980 2.795 2.990 3.029 ;
        RECT 2.990 2.805 3.000 3.039 ;
        RECT 3.000 2.815 3.010 3.049 ;
        RECT 3.010 2.825 3.020 3.059 ;
        RECT 3.020 2.835 3.030 3.069 ;
        RECT 3.030 2.845 3.040 3.079 ;
        RECT 3.040 2.855 3.050 3.089 ;
        RECT 3.050 2.865 3.060 3.099 ;
        RECT 3.060 2.875 3.070 3.109 ;
        RECT 3.070 2.885 3.080 3.119 ;
        RECT 3.080 2.895 3.090 3.129 ;
        RECT 3.090 2.905 3.100 3.139 ;
        RECT 2.810 1.415 2.820 2.859 ;
        RECT 2.820 1.415 2.830 2.869 ;
        RECT 2.830 1.415 2.840 2.879 ;
        RECT 2.840 1.415 2.850 2.889 ;
        RECT 2.850 1.415 2.860 2.899 ;
        RECT 2.860 1.415 2.870 2.909 ;
        RECT 2.870 1.415 2.880 2.919 ;
        RECT 2.880 1.415 2.890 2.929 ;
        RECT 2.890 1.415 2.900 2.939 ;
        RECT 2.900 1.415 2.910 2.949 ;
        RECT 2.910 1.415 2.920 2.959 ;
        RECT 2.920 1.415 2.930 2.969 ;
        RECT 2.930 1.415 2.940 2.979 ;
        RECT 2.940 1.415 2.950 2.989 ;
        RECT 2.950 1.415 2.960 2.999 ;
        RECT 2.960 1.415 2.970 3.009 ;
        RECT 2.340 2.625 2.350 2.859 ;
        RECT 2.350 2.635 2.360 2.859 ;
        RECT 2.360 2.645 2.370 2.859 ;
        RECT 2.370 2.655 2.380 2.859 ;
        RECT 2.380 2.665 2.390 2.859 ;
        RECT 2.390 2.675 2.400 2.859 ;
        RECT 2.400 2.685 2.410 2.859 ;
        RECT 2.410 2.690 2.416 2.860 ;
        RECT 2.120 2.405 2.130 2.639 ;
        RECT 2.130 2.415 2.140 2.649 ;
        RECT 2.140 2.425 2.150 2.659 ;
        RECT 2.150 2.435 2.160 2.669 ;
        RECT 2.160 2.445 2.170 2.679 ;
        RECT 2.170 2.455 2.180 2.689 ;
        RECT 2.180 2.465 2.190 2.699 ;
        RECT 2.190 2.475 2.200 2.709 ;
        RECT 2.200 2.485 2.210 2.719 ;
        RECT 2.210 2.495 2.220 2.729 ;
        RECT 2.220 2.505 2.230 2.739 ;
        RECT 2.230 2.515 2.240 2.749 ;
        RECT 2.240 2.525 2.250 2.759 ;
        RECT 2.250 2.535 2.260 2.769 ;
        RECT 2.260 2.545 2.270 2.779 ;
        RECT 2.270 2.555 2.280 2.789 ;
        RECT 2.280 2.565 2.290 2.799 ;
        RECT 2.290 2.575 2.300 2.809 ;
        RECT 2.300 2.585 2.310 2.819 ;
        RECT 2.310 2.595 2.320 2.829 ;
        RECT 2.320 2.605 2.330 2.839 ;
        RECT 2.330 2.615 2.340 2.849 ;
        RECT 2.045 2.395 2.055 2.565 ;
        RECT 2.055 2.395 2.065 2.575 ;
        RECT 2.065 2.395 2.075 2.585 ;
        RECT 2.075 2.395 2.085 2.595 ;
        RECT 2.085 2.395 2.095 2.605 ;
        RECT 2.095 2.395 2.105 2.615 ;
        RECT 2.105 2.395 2.115 2.625 ;
        RECT 2.115 2.395 2.121 2.635 ;
        RECT 3.150 2.395 3.325 2.695 ;
        RECT 3.180 1.045 3.665 1.215 ;
        RECT 3.495 1.045 3.665 2.630 ;
        RECT 3.150 2.395 3.665 2.630 ;
        RECT 3.150 2.455 4.885 2.630 ;
        RECT 4.585 2.195 4.885 3.045 ;
        RECT 5.330 1.595 5.500 2.370 ;
        RECT 4.585 2.195 5.500 2.370 ;
        RECT 3.960 1.605 4.130 2.015 ;
        RECT 4.895 1.245 5.065 2.015 ;
        RECT 3.960 1.845 5.065 2.015 ;
        RECT 5.425 1.060 5.595 1.415 ;
        RECT 4.895 1.245 5.850 1.415 ;
        RECT 5.680 1.245 5.850 2.640 ;
        RECT 7.400 1.540 7.570 2.640 ;
        RECT 5.680 2.460 7.570 2.640 ;
  END 
END LATRHD2XHT

MACRO LATRHD1XHT
  CLASS  CORE ;
  FOREIGN LATRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.380 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.840 0.720 6.170 1.200 ;
        RECT 6.000 0.720 6.170 2.280 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.040 0.720 7.210 2.960 ;
        RECT 7.040 1.260 7.280 1.610 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.595 2.090 2.135 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.460 0.520 2.840 ;
    END
  END G
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.355 0.645 1.525 0.945 ;
        RECT 2.080 0.575 2.250 0.945 ;
        RECT 1.355 0.775 2.250 0.945 ;
        RECT 4.120 0.500 4.635 0.745 ;
        RECT 2.080 0.575 4.635 0.745 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.715 ;
        RECT 1.725 -0.300 1.895 0.575 ;
        RECT 4.830 -0.300 5.000 1.155 ;
        RECT 4.700 0.985 5.000 1.155 ;
        RECT 6.455 -0.300 6.755 1.055 ;
        RECT 0.000 -0.300 7.380 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.730 2.740 0.900 3.990 ;
        RECT 1.595 3.095 1.895 3.990 ;
        RECT 4.010 2.505 4.310 3.990 ;
        RECT 4.980 2.650 5.280 3.990 ;
        RECT 6.455 2.975 6.755 3.990 ;
        RECT 0.000 3.390 7.380 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 0.860 1.755 ;
        RECT 1.250 2.745 1.975 2.915 ;
        RECT 2.285 2.975 2.825 3.145 ;
        RECT 2.205 2.905 2.215 3.145 ;
        RECT 2.215 2.915 2.225 3.145 ;
        RECT 2.225 2.925 2.235 3.145 ;
        RECT 2.235 2.935 2.245 3.145 ;
        RECT 2.245 2.945 2.255 3.145 ;
        RECT 2.255 2.955 2.265 3.145 ;
        RECT 2.265 2.965 2.275 3.145 ;
        RECT 2.275 2.975 2.285 3.145 ;
        RECT 2.055 2.755 2.065 2.995 ;
        RECT 2.065 2.765 2.075 3.005 ;
        RECT 2.075 2.775 2.085 3.015 ;
        RECT 2.085 2.785 2.095 3.025 ;
        RECT 2.095 2.795 2.105 3.035 ;
        RECT 2.105 2.805 2.115 3.045 ;
        RECT 2.115 2.815 2.125 3.055 ;
        RECT 2.125 2.825 2.135 3.065 ;
        RECT 2.135 2.835 2.145 3.075 ;
        RECT 2.145 2.845 2.155 3.085 ;
        RECT 2.155 2.855 2.165 3.095 ;
        RECT 2.165 2.865 2.175 3.105 ;
        RECT 2.175 2.875 2.185 3.115 ;
        RECT 2.185 2.885 2.195 3.125 ;
        RECT 2.195 2.895 2.205 3.135 ;
        RECT 1.975 2.745 1.985 2.915 ;
        RECT 1.985 2.745 1.995 2.925 ;
        RECT 1.995 2.745 2.005 2.935 ;
        RECT 2.005 2.745 2.015 2.945 ;
        RECT 2.015 2.745 2.025 2.955 ;
        RECT 2.025 2.745 2.035 2.965 ;
        RECT 2.035 2.745 2.045 2.975 ;
        RECT 2.045 2.745 2.055 2.985 ;
        RECT 1.080 2.420 1.090 2.914 ;
        RECT 1.090 2.430 1.100 2.914 ;
        RECT 1.100 2.440 1.110 2.914 ;
        RECT 1.110 2.450 1.120 2.914 ;
        RECT 1.120 2.460 1.130 2.914 ;
        RECT 1.130 2.470 1.140 2.914 ;
        RECT 1.140 2.480 1.150 2.914 ;
        RECT 1.150 2.490 1.160 2.914 ;
        RECT 1.160 2.500 1.170 2.914 ;
        RECT 1.170 2.510 1.180 2.914 ;
        RECT 1.180 2.520 1.190 2.914 ;
        RECT 1.190 2.530 1.200 2.914 ;
        RECT 1.200 2.540 1.210 2.914 ;
        RECT 1.210 2.550 1.220 2.914 ;
        RECT 1.220 2.560 1.230 2.914 ;
        RECT 1.230 2.570 1.240 2.914 ;
        RECT 1.240 2.580 1.250 2.914 ;
        RECT 1.030 2.370 1.040 2.604 ;
        RECT 1.040 2.380 1.050 2.614 ;
        RECT 1.050 2.390 1.060 2.624 ;
        RECT 1.060 2.400 1.070 2.634 ;
        RECT 1.070 2.410 1.080 2.644 ;
        RECT 0.860 1.520 0.870 2.434 ;
        RECT 0.870 1.520 0.880 2.444 ;
        RECT 0.880 1.520 0.890 2.454 ;
        RECT 0.890 1.520 0.900 2.464 ;
        RECT 0.900 1.520 0.910 2.474 ;
        RECT 0.910 1.520 0.920 2.484 ;
        RECT 0.920 1.520 0.930 2.494 ;
        RECT 0.930 1.520 0.940 2.504 ;
        RECT 0.940 1.520 0.950 2.514 ;
        RECT 0.950 1.520 0.960 2.524 ;
        RECT 0.960 1.520 0.970 2.534 ;
        RECT 0.970 1.520 0.980 2.544 ;
        RECT 0.980 1.520 0.990 2.554 ;
        RECT 0.990 1.520 1.000 2.564 ;
        RECT 1.000 1.520 1.010 2.574 ;
        RECT 1.010 1.520 1.020 2.584 ;
        RECT 1.020 1.520 1.030 2.594 ;
        RECT 2.445 0.925 2.615 2.235 ;
        RECT 2.300 2.065 2.615 2.235 ;
        RECT 2.445 0.925 2.945 1.095 ;
        RECT 1.085 1.125 1.210 1.295 ;
        RECT 1.585 2.395 2.135 2.565 ;
        RECT 2.805 1.295 2.900 2.795 ;
        RECT 2.445 2.625 2.900 2.795 ;
        RECT 2.975 1.295 3.225 1.465 ;
        RECT 3.125 2.775 3.570 2.945 ;
        RECT 3.050 2.710 3.060 2.944 ;
        RECT 3.060 2.720 3.070 2.944 ;
        RECT 3.070 2.730 3.080 2.944 ;
        RECT 3.080 2.740 3.090 2.944 ;
        RECT 3.090 2.750 3.100 2.944 ;
        RECT 3.100 2.760 3.110 2.944 ;
        RECT 3.110 2.770 3.120 2.944 ;
        RECT 3.120 2.775 3.126 2.945 ;
        RECT 2.975 2.635 2.985 2.869 ;
        RECT 2.985 2.645 2.995 2.879 ;
        RECT 2.995 2.655 3.005 2.889 ;
        RECT 3.005 2.665 3.015 2.899 ;
        RECT 3.015 2.675 3.025 2.909 ;
        RECT 3.025 2.685 3.035 2.919 ;
        RECT 3.035 2.695 3.045 2.929 ;
        RECT 3.045 2.700 3.051 2.940 ;
        RECT 2.900 1.295 2.910 2.795 ;
        RECT 2.910 1.295 2.920 2.805 ;
        RECT 2.920 1.295 2.930 2.815 ;
        RECT 2.930 1.295 2.940 2.825 ;
        RECT 2.940 1.295 2.950 2.835 ;
        RECT 2.950 1.295 2.960 2.845 ;
        RECT 2.960 1.295 2.970 2.855 ;
        RECT 2.970 1.295 2.976 2.865 ;
        RECT 2.365 2.555 2.375 2.795 ;
        RECT 2.375 2.565 2.385 2.795 ;
        RECT 2.385 2.575 2.395 2.795 ;
        RECT 2.395 2.585 2.405 2.795 ;
        RECT 2.405 2.595 2.415 2.795 ;
        RECT 2.415 2.605 2.425 2.795 ;
        RECT 2.425 2.615 2.435 2.795 ;
        RECT 2.435 2.625 2.445 2.795 ;
        RECT 2.215 2.405 2.225 2.645 ;
        RECT 2.225 2.415 2.235 2.655 ;
        RECT 2.235 2.425 2.245 2.665 ;
        RECT 2.245 2.435 2.255 2.675 ;
        RECT 2.255 2.445 2.265 2.685 ;
        RECT 2.265 2.455 2.275 2.695 ;
        RECT 2.275 2.465 2.285 2.705 ;
        RECT 2.285 2.475 2.295 2.715 ;
        RECT 2.295 2.485 2.305 2.725 ;
        RECT 2.305 2.495 2.315 2.735 ;
        RECT 2.315 2.505 2.325 2.745 ;
        RECT 2.325 2.515 2.335 2.755 ;
        RECT 2.335 2.525 2.345 2.765 ;
        RECT 2.345 2.535 2.355 2.775 ;
        RECT 2.355 2.545 2.365 2.785 ;
        RECT 2.135 2.395 2.145 2.565 ;
        RECT 2.145 2.395 2.155 2.575 ;
        RECT 2.155 2.395 2.165 2.585 ;
        RECT 2.165 2.395 2.175 2.595 ;
        RECT 2.175 2.395 2.185 2.605 ;
        RECT 2.185 2.395 2.195 2.615 ;
        RECT 2.195 2.395 2.205 2.625 ;
        RECT 2.205 2.395 2.215 2.635 ;
        RECT 1.495 2.315 1.505 2.565 ;
        RECT 1.505 2.325 1.515 2.565 ;
        RECT 1.515 2.335 1.525 2.565 ;
        RECT 1.525 2.345 1.535 2.565 ;
        RECT 1.535 2.355 1.545 2.565 ;
        RECT 1.545 2.365 1.555 2.565 ;
        RECT 1.555 2.375 1.565 2.565 ;
        RECT 1.565 2.385 1.575 2.565 ;
        RECT 1.575 2.395 1.585 2.565 ;
        RECT 1.405 2.225 1.415 2.475 ;
        RECT 1.415 2.235 1.425 2.485 ;
        RECT 1.425 2.245 1.435 2.495 ;
        RECT 1.435 2.255 1.445 2.505 ;
        RECT 1.445 2.265 1.455 2.515 ;
        RECT 1.455 2.275 1.465 2.525 ;
        RECT 1.465 2.285 1.475 2.535 ;
        RECT 1.475 2.295 1.485 2.545 ;
        RECT 1.485 2.305 1.495 2.555 ;
        RECT 1.210 1.125 1.220 2.279 ;
        RECT 1.220 1.125 1.230 2.289 ;
        RECT 1.230 1.125 1.240 2.299 ;
        RECT 1.240 1.125 1.250 2.309 ;
        RECT 1.250 1.125 1.260 2.319 ;
        RECT 1.260 1.125 1.270 2.329 ;
        RECT 1.270 1.125 1.280 2.339 ;
        RECT 1.280 1.125 1.290 2.349 ;
        RECT 1.290 1.125 1.300 2.359 ;
        RECT 1.300 1.125 1.310 2.369 ;
        RECT 1.310 1.125 1.320 2.379 ;
        RECT 1.320 1.125 1.330 2.389 ;
        RECT 1.330 1.125 1.340 2.399 ;
        RECT 1.340 1.125 1.350 2.409 ;
        RECT 1.350 1.125 1.360 2.419 ;
        RECT 1.360 1.125 1.370 2.429 ;
        RECT 1.370 1.125 1.380 2.439 ;
        RECT 1.380 1.125 1.390 2.449 ;
        RECT 1.390 1.125 1.400 2.459 ;
        RECT 1.400 1.125 1.406 2.469 ;
        RECT 3.155 2.045 3.325 2.520 ;
        RECT 3.165 0.925 3.705 1.095 ;
        RECT 3.535 0.925 3.705 2.215 ;
        RECT 5.060 1.980 5.360 2.215 ;
        RECT 3.155 2.045 5.360 2.215 ;
        RECT 5.345 0.920 5.515 1.685 ;
        RECT 3.900 1.515 5.735 1.685 ;
        RECT 5.565 1.515 5.735 2.765 ;
        RECT 6.660 1.540 6.830 2.630 ;
        RECT 5.565 2.460 6.830 2.630 ;
  END 
END LATRHD1XHT

MACRO LATHD1XSPGHT
  CLASS  CORE ;
  FOREIGN LATHD1XSPGHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.150 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 5.265 0.300 5.805 3.075 ;
      LAYER V7 ;
        RECT 5.355 1.665 5.715 2.025 ;
      LAYER M7 ;
        RECT 5.025 1.655 5.805 2.035 ;
      LAYER V6 ;
        RECT 5.440 1.750 5.630 1.940 ;
      LAYER M4 ;
        RECT 5.435 1.365 5.635 2.170 ;
      LAYER V3 ;
        RECT 5.440 1.750 5.630 1.940 ;
      LAYER M3 ;
        RECT 5.205 1.745 6.045 1.945 ;
        RECT 5.845 1.670 6.045 2.010 ;
      LAYER V2 ;
        RECT 5.850 1.750 6.040 1.940 ;
      LAYER M2 ;
        RECT 5.845 1.670 6.045 2.425 ;
      LAYER V1 ;
        RECT 5.850 2.160 6.040 2.350 ;
      LAYER M1 ;
        RECT 5.770 0.720 5.940 2.960 ;
        RECT 5.770 2.090 6.050 2.425 ;
      LAYER M6 ;
        RECT 5.435 1.060 5.635 2.475 ;
      LAYER V5 ;
        RECT 5.440 1.750 5.630 1.940 ;
      LAYER M5 ;
        RECT 5.025 1.745 5.805 1.945 ;
      LAYER V4 ;
        RECT 5.440 1.750 5.630 1.940 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 4.035 0.300 4.575 3.075 ;
      LAYER V7 ;
        RECT 4.125 0.845 4.485 1.205 ;
      LAYER M7 ;
        RECT 4.035 0.835 4.815 1.215 ;
      LAYER V6 ;
        RECT 4.210 0.930 4.400 1.120 ;
      LAYER M4 ;
        RECT 4.615 0.590 4.815 1.420 ;
      LAYER V3 ;
        RECT 4.620 0.930 4.810 1.120 ;
      LAYER M3 ;
        RECT 4.255 0.925 5.180 1.125 ;
      LAYER V2 ;
        RECT 4.620 0.930 4.810 1.120 ;
      LAYER M2 ;
        RECT 4.615 0.565 4.815 1.435 ;
      LAYER V1 ;
        RECT 4.620 0.930 4.810 1.120 ;
      LAYER M1 ;
        RECT 4.610 0.850 4.900 1.205 ;
        RECT 4.730 0.720 4.900 2.280 ;
      LAYER M6 ;
        RECT 4.205 0.510 4.405 2.475 ;
      LAYER V5 ;
        RECT 4.210 0.930 4.400 1.120 ;
      LAYER M5 ;
        RECT 4.035 0.925 4.915 1.125 ;
      LAYER V4 ;
        RECT 4.620 0.930 4.810 1.120 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 1.575 0.300 2.115 3.075 ;
      LAYER V7 ;
        RECT 1.665 1.255 2.025 1.615 ;
      LAYER M7 ;
        RECT 1.515 1.245 2.250 1.625 ;
      LAYER V6 ;
        RECT 1.750 1.340 1.940 1.530 ;
      LAYER M4 ;
        RECT 1.745 1.095 1.945 1.915 ;
      LAYER V3 ;
        RECT 1.750 1.340 1.940 1.530 ;
      LAYER M3 ;
        RECT 1.485 1.335 2.300 1.535 ;
      LAYER V2 ;
        RECT 1.750 1.340 1.940 1.530 ;
      LAYER M2 ;
        RECT 1.745 1.215 1.945 2.025 ;
      LAYER V1 ;
        RECT 1.750 1.750 1.940 1.940 ;
      LAYER M1 ;
        RECT 1.680 1.585 2.135 1.950 ;
      LAYER M6 ;
        RECT 1.745 1.055 1.945 3.075 ;
      LAYER V5 ;
        RECT 1.750 1.340 1.940 1.530 ;
      LAYER M5 ;
        RECT 1.515 1.335 2.250 1.535 ;
      LAYER V4 ;
        RECT 1.750 1.340 1.940 1.530 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 0.345 0.300 0.885 3.075 ;
      LAYER V7 ;
        RECT 0.435 2.075 0.795 2.435 ;
      LAYER M7 ;
        RECT 0.315 2.065 1.050 2.445 ;
      LAYER V6 ;
        RECT 0.520 2.160 0.710 2.350 ;
      LAYER M4 ;
        RECT 0.515 1.845 0.715 2.600 ;
      LAYER V3 ;
        RECT 0.520 2.160 0.710 2.350 ;
      LAYER M3 ;
        RECT 0.105 2.060 0.305 2.425 ;
        RECT 0.105 2.155 0.885 2.355 ;
      LAYER V2 ;
        RECT 0.110 2.160 0.300 2.350 ;
      LAYER M2 ;
        RECT 0.105 2.060 0.305 2.865 ;
      LAYER V1 ;
        RECT 0.110 2.570 0.300 2.760 ;
      LAYER M1 ;
        RECT 0.100 2.495 0.510 2.955 ;
      LAYER M6 ;
        RECT 0.515 1.055 0.715 3.075 ;
      LAYER V5 ;
        RECT 0.520 2.160 0.710 2.350 ;
      LAYER M5 ;
        RECT 0.315 2.155 1.050 2.355 ;
      LAYER V4 ;
        RECT 0.520 2.160 0.710 2.350 ;
    END
  END G
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 1.625 -0.300 1.925 0.780 ;
        RECT 3.435 -0.300 3.735 1.295 ;
        RECT 5.185 -0.300 5.485 1.055 ;
        RECT 0.000 -0.300 6.150 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.280 0.860 3.990 ;
        RECT 1.655 2.545 1.955 3.990 ;
        RECT 3.405 2.995 3.705 3.990 ;
        RECT 5.185 2.975 5.485 3.990 ;
        RECT 0.000 3.390 6.150 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.520 1.030 1.820 ;
        RECT 1.210 1.060 1.380 2.300 ;
        RECT 1.210 2.130 2.375 2.300 ;
        RECT 2.205 2.130 2.375 3.095 ;
        RECT 2.260 0.605 2.430 1.230 ;
        RECT 1.210 1.060 2.430 1.230 ;
        RECT 2.260 0.605 2.665 0.775 ;
        RECT 2.205 2.925 3.025 3.095 ;
        RECT 3.255 1.850 3.555 2.020 ;
        RECT 3.385 1.850 3.555 2.395 ;
        RECT 3.955 1.125 4.430 1.295 ;
        RECT 4.260 1.125 4.430 2.395 ;
        RECT 3.385 2.225 4.430 2.395 ;
        RECT 4.260 1.520 4.550 1.820 ;
        RECT 2.610 1.060 2.780 2.745 ;
        RECT 2.610 1.500 4.075 1.670 ;
        RECT 5.420 1.520 5.590 2.745 ;
        RECT 2.610 2.575 5.590 2.745 ;
  END 
END LATHD1XSPGHT

MACRO INVTSHD16XHT
  CLASS  CORE ;
  FOREIGN INVTSHD16XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.270 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 17.865 1.325 18.525 1.780 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.675 0.535 2.045 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.055 ;
        RECT 1.665 -0.300 1.965 1.055 ;
        RECT 5.865 -0.300 6.165 1.055 ;
        RECT 6.905 -0.300 7.205 1.055 ;
        RECT 7.945 -0.300 8.245 1.055 ;
        RECT 8.985 -0.300 9.285 1.055 ;
        RECT 10.025 -0.300 10.325 1.055 ;
        RECT 11.065 -0.300 11.365 1.055 ;
        RECT 12.105 -0.300 12.405 1.055 ;
        RECT 13.145 -0.300 13.445 1.055 ;
        RECT 14.405 -0.300 14.705 0.715 ;
        RECT 15.445 -0.300 15.745 0.715 ;
        RECT 16.485 -0.300 16.785 0.715 ;
        RECT 17.525 -0.300 17.825 0.715 ;
        RECT 18.565 -0.300 18.865 1.055 ;
        RECT 0.000 -0.300 19.270 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 5.410 0.720 5.580 2.960 ;
        RECT 6.445 0.785 6.625 2.965 ;
        RECT 6.385 0.785 6.685 1.980 ;
        RECT 7.485 0.785 7.665 2.960 ;
        RECT 7.425 0.785 7.725 1.980 ;
        RECT 8.530 0.785 8.700 2.965 ;
        RECT 8.465 0.785 8.765 1.980 ;
        RECT 9.570 0.785 9.740 2.965 ;
        RECT 9.505 0.785 9.805 1.980 ;
        RECT 10.610 0.785 10.780 2.960 ;
        RECT 10.545 0.785 10.845 1.980 ;
        RECT 11.650 0.785 11.820 2.960 ;
        RECT 11.585 0.785 11.885 1.980 ;
        RECT 12.690 0.760 12.860 2.960 ;
        RECT 12.625 0.760 12.925 1.980 ;
        RECT 5.410 1.360 13.900 1.980 ;
        RECT 13.720 0.720 13.900 2.965 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.595 0.925 3.990 ;
        RECT 1.665 2.975 1.965 3.990 ;
        RECT 5.865 2.295 6.165 3.990 ;
        RECT 6.905 2.295 7.205 3.990 ;
        RECT 7.945 2.295 8.245 3.990 ;
        RECT 8.985 2.295 9.285 3.990 ;
        RECT 10.025 2.295 10.325 3.990 ;
        RECT 11.065 2.295 11.365 3.990 ;
        RECT 12.105 2.295 12.405 3.990 ;
        RECT 13.145 2.295 13.445 3.990 ;
        RECT 14.405 2.570 14.705 3.990 ;
        RECT 15.445 2.295 15.745 3.990 ;
        RECT 16.485 2.295 16.785 3.990 ;
        RECT 17.525 2.635 17.825 3.990 ;
        RECT 18.565 2.295 18.865 3.990 ;
        RECT 0.000 3.390 19.270 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.160 0.610 0.350 1.440 ;
        RECT 0.160 2.225 0.350 3.205 ;
        RECT 0.160 1.250 1.015 1.440 ;
        RECT 0.825 1.250 1.015 2.415 ;
        RECT 0.160 2.225 1.015 2.415 ;
        RECT 0.825 1.770 3.610 2.070 ;
        RECT 1.200 0.720 1.400 1.515 ;
        RECT 2.240 0.720 2.420 1.515 ;
        RECT 2.750 0.720 2.930 1.515 ;
        RECT 1.200 1.315 3.990 1.515 ;
        RECT 3.790 1.040 3.990 2.420 ;
        RECT 2.695 2.250 4.035 2.420 ;
        RECT 3.790 1.160 4.860 1.460 ;
        RECT 1.205 2.265 1.385 2.905 ;
        RECT 1.205 2.265 2.485 2.465 ;
        RECT 2.185 2.265 2.485 2.885 ;
        RECT 3.215 0.560 3.515 1.135 ;
        RECT 4.255 2.245 4.555 2.885 ;
        RECT 2.185 2.705 4.555 2.885 ;
        RECT 3.215 0.560 5.210 0.860 ;
        RECT 5.040 0.560 5.210 2.465 ;
        RECT 4.255 2.245 5.210 2.465 ;
        RECT 14.095 1.180 14.275 1.570 ;
        RECT 14.990 0.720 15.160 1.360 ;
        RECT 16.030 0.720 16.200 1.360 ;
        RECT 17.060 0.720 17.240 1.360 ;
        RECT 14.095 1.180 17.240 1.360 ;
        RECT 14.095 1.770 14.275 2.105 ;
        RECT 14.970 1.925 15.170 2.960 ;
        RECT 16.015 1.925 16.215 2.960 ;
        RECT 14.095 1.925 17.245 2.105 ;
        RECT 17.065 1.925 17.245 2.960 ;
        RECT 14.910 1.575 17.620 1.745 ;
        RECT 17.430 0.930 17.620 2.390 ;
        RECT 17.430 2.200 18.285 2.390 ;
        RECT 18.095 2.200 18.285 3.180 ;
        RECT 18.100 0.480 18.290 1.120 ;
        RECT 17.430 0.930 18.290 1.120 ;
  END 
END INVTSHD16XHT

MACRO LATNSRHD1XHT
  CLASS  CORE ;
  FOREIGN LATNSRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.430 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.205 1.125 7.375 3.145 ;
        RECT 6.970 2.470 7.375 3.145 ;
        RECT 7.105 1.125 7.405 1.295 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.565 0.965 2.055 ;
        RECT 0.510 1.565 1.040 1.865 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.090 0.715 9.330 2.960 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.970 1.185 3.180 1.910 ;
        RECT 2.970 1.610 3.370 1.910 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.020 0.480 5.230 1.235 ;
        RECT 5.020 0.480 5.705 0.650 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 2.265 -0.300 2.565 0.595 ;
        RECT 5.885 -0.300 6.055 1.085 ;
        RECT 7.770 -0.300 8.070 0.715 ;
        RECT 8.505 -0.300 8.805 0.715 ;
        RECT 0.000 -0.300 9.430 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.355 2.745 2.035 3.180 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.905 0.895 3.990 ;
        RECT 2.270 2.745 2.440 3.990 ;
        RECT 5.630 2.430 5.930 3.990 ;
        RECT 7.555 2.230 7.725 3.990 ;
        RECT 8.505 2.630 8.825 3.990 ;
        RECT 0.000 3.390 9.430 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.655 1.125 1.955 1.295 ;
        RECT 1.785 1.125 1.955 2.215 ;
        RECT 1.655 2.045 1.955 2.215 ;
        RECT 1.785 1.610 2.550 1.910 ;
        RECT 3.420 1.125 3.720 1.295 ;
        RECT 3.550 1.125 3.720 2.325 ;
        RECT 3.235 2.155 3.720 2.325 ;
        RECT 1.210 0.625 1.445 1.360 ;
        RECT 1.275 0.625 1.445 2.215 ;
        RECT 1.145 2.045 1.445 2.215 ;
        RECT 1.210 0.625 1.585 0.945 ;
        RECT 2.975 0.605 3.145 0.945 ;
        RECT 1.210 0.775 3.145 0.945 ;
        RECT 2.975 0.605 3.960 0.775 ;
        RECT 0.105 1.060 0.275 2.565 ;
        RECT 0.105 1.060 0.340 1.360 ;
        RECT 0.105 2.345 0.405 2.565 ;
        RECT 2.665 2.395 2.890 2.710 ;
        RECT 0.105 2.395 2.890 2.565 ;
        RECT 2.665 2.505 3.900 2.710 ;
        RECT 3.760 2.505 3.900 2.860 ;
        RECT 4.540 0.605 4.840 1.020 ;
        RECT 4.265 0.820 4.840 1.020 ;
        RECT 4.180 0.820 4.190 1.094 ;
        RECT 4.190 0.820 4.200 1.084 ;
        RECT 4.200 0.820 4.210 1.074 ;
        RECT 4.210 0.820 4.220 1.064 ;
        RECT 4.220 0.820 4.230 1.054 ;
        RECT 4.230 0.820 4.240 1.044 ;
        RECT 4.240 0.820 4.250 1.034 ;
        RECT 4.250 0.820 4.260 1.024 ;
        RECT 4.260 0.820 4.266 1.020 ;
        RECT 4.070 0.930 4.080 1.204 ;
        RECT 4.080 0.920 4.090 1.194 ;
        RECT 4.090 0.910 4.100 1.184 ;
        RECT 4.100 0.900 4.110 1.174 ;
        RECT 4.110 0.890 4.120 1.164 ;
        RECT 4.120 0.880 4.130 1.154 ;
        RECT 4.130 0.870 4.140 1.144 ;
        RECT 4.140 0.860 4.150 1.134 ;
        RECT 4.150 0.850 4.160 1.124 ;
        RECT 4.160 0.840 4.170 1.114 ;
        RECT 4.170 0.830 4.180 1.104 ;
        RECT 3.900 1.100 3.910 2.860 ;
        RECT 3.910 1.090 3.920 2.860 ;
        RECT 3.920 1.080 3.930 2.860 ;
        RECT 3.930 1.070 3.940 2.860 ;
        RECT 3.940 1.060 3.950 2.860 ;
        RECT 3.950 1.050 3.960 2.860 ;
        RECT 3.960 1.040 3.970 2.860 ;
        RECT 3.970 1.030 3.980 2.860 ;
        RECT 3.980 1.020 3.990 2.860 ;
        RECT 3.990 1.010 4.000 2.860 ;
        RECT 4.000 1.000 4.010 2.860 ;
        RECT 4.010 0.990 4.020 2.860 ;
        RECT 4.020 0.980 4.030 2.860 ;
        RECT 4.030 0.970 4.040 2.860 ;
        RECT 4.040 0.960 4.050 2.860 ;
        RECT 4.050 0.950 4.060 2.860 ;
        RECT 4.060 0.940 4.070 2.860 ;
        RECT 2.640 2.910 2.810 3.210 ;
        RECT 3.395 2.910 3.580 3.210 ;
        RECT 2.640 2.910 3.580 3.090 ;
        RECT 4.215 3.000 4.385 3.210 ;
        RECT 3.395 3.040 4.385 3.210 ;
        RECT 4.215 3.000 5.130 3.170 ;
        RECT 6.405 0.480 6.575 1.085 ;
        RECT 6.405 0.480 6.810 0.650 ;
        RECT 4.345 1.200 4.520 2.355 ;
        RECT 4.345 1.200 4.645 1.370 ;
        RECT 6.690 1.630 6.860 2.240 ;
        RECT 4.345 2.070 6.860 2.240 ;
        RECT 6.690 1.630 7.025 1.800 ;
        RECT 6.180 1.265 6.400 1.845 ;
        RECT 4.970 1.675 6.400 1.845 ;
        RECT 6.180 1.265 6.755 1.450 ;
        RECT 7.025 0.775 7.485 0.945 ;
        RECT 7.755 0.960 8.320 1.130 ;
        RECT 8.150 0.960 8.320 2.280 ;
        RECT 8.110 1.980 8.320 2.280 ;
        RECT 8.150 1.515 8.910 1.815 ;
        RECT 7.670 0.885 7.680 1.129 ;
        RECT 7.680 0.895 7.690 1.129 ;
        RECT 7.690 0.905 7.700 1.129 ;
        RECT 7.700 0.915 7.710 1.129 ;
        RECT 7.710 0.925 7.720 1.129 ;
        RECT 7.720 0.935 7.730 1.129 ;
        RECT 7.730 0.945 7.740 1.129 ;
        RECT 7.740 0.955 7.750 1.129 ;
        RECT 7.750 0.960 7.756 1.130 ;
        RECT 7.570 0.785 7.580 1.029 ;
        RECT 7.580 0.795 7.590 1.039 ;
        RECT 7.590 0.805 7.600 1.049 ;
        RECT 7.600 0.815 7.610 1.059 ;
        RECT 7.610 0.825 7.620 1.069 ;
        RECT 7.620 0.835 7.630 1.079 ;
        RECT 7.630 0.845 7.640 1.089 ;
        RECT 7.640 0.855 7.650 1.099 ;
        RECT 7.650 0.865 7.660 1.109 ;
        RECT 7.660 0.875 7.670 1.119 ;
        RECT 7.485 0.775 7.495 0.945 ;
        RECT 7.495 0.775 7.505 0.955 ;
        RECT 7.505 0.775 7.515 0.965 ;
        RECT 7.515 0.775 7.525 0.975 ;
        RECT 7.525 0.775 7.535 0.985 ;
        RECT 7.535 0.775 7.545 0.995 ;
        RECT 7.545 0.775 7.555 1.005 ;
        RECT 7.555 0.775 7.565 1.015 ;
        RECT 7.565 0.775 7.571 1.025 ;
        RECT 6.945 0.775 6.955 1.015 ;
        RECT 6.955 0.775 6.965 1.005 ;
        RECT 6.965 0.775 6.975 0.995 ;
        RECT 6.975 0.775 6.985 0.985 ;
        RECT 6.985 0.775 6.995 0.975 ;
        RECT 6.995 0.775 7.005 0.965 ;
        RECT 7.005 0.775 7.015 0.955 ;
        RECT 7.015 0.775 7.025 0.945 ;
        RECT 6.925 0.795 6.935 1.035 ;
        RECT 6.935 0.785 6.945 1.025 ;
        RECT 6.755 0.965 6.765 1.449 ;
        RECT 6.765 0.955 6.775 1.449 ;
        RECT 6.775 0.945 6.785 1.449 ;
        RECT 6.785 0.935 6.795 1.449 ;
        RECT 6.795 0.925 6.805 1.449 ;
        RECT 6.805 0.915 6.815 1.449 ;
        RECT 6.815 0.905 6.825 1.449 ;
        RECT 6.825 0.895 6.835 1.449 ;
        RECT 6.835 0.885 6.845 1.449 ;
        RECT 6.845 0.875 6.855 1.449 ;
        RECT 6.855 0.865 6.865 1.449 ;
        RECT 6.865 0.855 6.875 1.449 ;
        RECT 6.875 0.845 6.885 1.449 ;
        RECT 6.885 0.835 6.895 1.449 ;
        RECT 6.895 0.825 6.905 1.449 ;
        RECT 6.905 0.815 6.915 1.449 ;
        RECT 6.915 0.805 6.925 1.449 ;
  END 
END LATNSRHD1XHT

MACRO LATNSHDMXHT
  CLASS  CORE ;
  FOREIGN LATNSHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.790 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 6.410 1.060 6.580 2.280 ;
        RECT 6.410 1.660 6.895 2.025 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.520 3.000 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.450 1.060 7.645 2.280 ;
        RECT 7.450 1.245 7.690 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.340 2.480 4.640 3.210 ;
        RECT 4.340 2.480 4.825 2.840 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.540 -0.300 0.840 0.715 ;
        RECT 2.255 -0.300 2.425 1.060 ;
        RECT 4.415 -0.300 4.715 0.595 ;
        RECT 5.375 -0.300 5.675 0.720 ;
        RECT 6.865 -0.300 7.165 1.145 ;
        RECT 0.000 -0.300 7.790 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.620 0.510 2.045 0.945 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.730 2.855 0.900 3.990 ;
        RECT 2.060 3.095 2.360 3.990 ;
        RECT 5.245 2.405 5.545 3.990 ;
        RECT 6.835 2.925 7.135 3.990 ;
        RECT 0.000 3.390 7.790 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 3.045 1.060 3.215 2.390 ;
        RECT 1.525 2.395 2.715 2.565 ;
        RECT 3.395 1.720 3.565 2.740 ;
        RECT 2.970 2.570 3.565 2.740 ;
        RECT 2.890 2.500 2.900 2.740 ;
        RECT 2.900 2.510 2.910 2.740 ;
        RECT 2.910 2.520 2.920 2.740 ;
        RECT 2.920 2.530 2.930 2.740 ;
        RECT 2.930 2.540 2.940 2.740 ;
        RECT 2.940 2.550 2.950 2.740 ;
        RECT 2.950 2.560 2.960 2.740 ;
        RECT 2.960 2.570 2.970 2.740 ;
        RECT 2.795 2.405 2.805 2.645 ;
        RECT 2.805 2.415 2.815 2.655 ;
        RECT 2.815 2.425 2.825 2.665 ;
        RECT 2.825 2.435 2.835 2.675 ;
        RECT 2.835 2.445 2.845 2.685 ;
        RECT 2.845 2.455 2.855 2.695 ;
        RECT 2.855 2.465 2.865 2.705 ;
        RECT 2.865 2.475 2.875 2.715 ;
        RECT 2.875 2.485 2.885 2.725 ;
        RECT 2.885 2.490 2.891 2.734 ;
        RECT 2.715 2.395 2.725 2.565 ;
        RECT 2.725 2.395 2.735 2.575 ;
        RECT 2.735 2.395 2.745 2.585 ;
        RECT 2.745 2.395 2.755 2.595 ;
        RECT 2.755 2.395 2.765 2.605 ;
        RECT 2.765 2.395 2.775 2.615 ;
        RECT 2.775 2.395 2.785 2.625 ;
        RECT 2.785 2.395 2.795 2.635 ;
        RECT 1.450 2.330 1.460 2.564 ;
        RECT 1.460 2.340 1.470 2.564 ;
        RECT 1.470 2.350 1.480 2.564 ;
        RECT 1.480 2.360 1.490 2.564 ;
        RECT 1.490 2.370 1.500 2.564 ;
        RECT 1.500 2.380 1.510 2.564 ;
        RECT 1.510 2.390 1.520 2.564 ;
        RECT 1.520 2.395 1.526 2.565 ;
        RECT 1.360 2.240 1.370 2.474 ;
        RECT 1.370 2.250 1.380 2.484 ;
        RECT 1.380 2.260 1.390 2.494 ;
        RECT 1.390 2.270 1.400 2.504 ;
        RECT 1.400 2.280 1.410 2.514 ;
        RECT 1.410 2.290 1.420 2.524 ;
        RECT 1.420 2.300 1.430 2.534 ;
        RECT 1.430 2.310 1.440 2.544 ;
        RECT 1.440 2.320 1.450 2.554 ;
        RECT 1.185 1.060 1.195 2.300 ;
        RECT 1.195 1.060 1.205 2.310 ;
        RECT 1.205 1.060 1.215 2.320 ;
        RECT 1.215 1.060 1.225 2.330 ;
        RECT 1.225 1.060 1.235 2.340 ;
        RECT 1.235 1.060 1.245 2.350 ;
        RECT 1.245 1.060 1.255 2.360 ;
        RECT 1.255 1.060 1.265 2.370 ;
        RECT 1.265 1.060 1.275 2.380 ;
        RECT 1.275 1.060 1.285 2.390 ;
        RECT 1.285 1.060 1.295 2.400 ;
        RECT 1.295 1.060 1.305 2.410 ;
        RECT 1.305 1.060 1.315 2.420 ;
        RECT 1.315 1.060 1.325 2.430 ;
        RECT 1.325 1.060 1.335 2.440 ;
        RECT 1.335 1.060 1.345 2.450 ;
        RECT 1.345 1.060 1.355 2.460 ;
        RECT 1.355 1.060 1.361 2.470 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.520 0.835 1.755 ;
        RECT 1.250 2.745 2.545 2.915 ;
        RECT 3.895 2.760 4.065 3.145 ;
        RECT 2.850 2.975 4.065 3.145 ;
        RECT 2.775 2.910 2.785 3.144 ;
        RECT 2.785 2.920 2.795 3.144 ;
        RECT 2.795 2.930 2.805 3.144 ;
        RECT 2.805 2.940 2.815 3.144 ;
        RECT 2.815 2.950 2.825 3.144 ;
        RECT 2.825 2.960 2.835 3.144 ;
        RECT 2.835 2.970 2.845 3.144 ;
        RECT 2.845 2.975 2.851 3.145 ;
        RECT 2.620 2.755 2.630 2.989 ;
        RECT 2.630 2.765 2.640 2.999 ;
        RECT 2.640 2.775 2.650 3.009 ;
        RECT 2.650 2.785 2.660 3.019 ;
        RECT 2.660 2.795 2.670 3.029 ;
        RECT 2.670 2.805 2.680 3.039 ;
        RECT 2.680 2.815 2.690 3.049 ;
        RECT 2.690 2.825 2.700 3.059 ;
        RECT 2.700 2.835 2.710 3.069 ;
        RECT 2.710 2.845 2.720 3.079 ;
        RECT 2.720 2.855 2.730 3.089 ;
        RECT 2.730 2.865 2.740 3.099 ;
        RECT 2.740 2.875 2.750 3.109 ;
        RECT 2.750 2.885 2.760 3.119 ;
        RECT 2.760 2.895 2.770 3.129 ;
        RECT 2.770 2.900 2.776 3.140 ;
        RECT 2.545 2.745 2.555 2.915 ;
        RECT 2.555 2.745 2.565 2.925 ;
        RECT 2.565 2.745 2.575 2.935 ;
        RECT 2.575 2.745 2.585 2.945 ;
        RECT 2.585 2.745 2.595 2.955 ;
        RECT 2.595 2.745 2.605 2.965 ;
        RECT 2.605 2.745 2.615 2.975 ;
        RECT 2.615 2.745 2.621 2.985 ;
        RECT 1.080 2.460 1.090 2.914 ;
        RECT 1.090 2.470 1.100 2.914 ;
        RECT 1.100 2.480 1.110 2.914 ;
        RECT 1.110 2.490 1.120 2.914 ;
        RECT 1.120 2.500 1.130 2.914 ;
        RECT 1.130 2.510 1.140 2.914 ;
        RECT 1.140 2.520 1.150 2.914 ;
        RECT 1.150 2.530 1.160 2.914 ;
        RECT 1.160 2.540 1.170 2.914 ;
        RECT 1.170 2.550 1.180 2.914 ;
        RECT 1.180 2.560 1.190 2.914 ;
        RECT 1.190 2.570 1.200 2.914 ;
        RECT 1.200 2.580 1.210 2.914 ;
        RECT 1.210 2.590 1.220 2.914 ;
        RECT 1.220 2.600 1.230 2.914 ;
        RECT 1.230 2.610 1.240 2.914 ;
        RECT 1.240 2.620 1.250 2.914 ;
        RECT 1.005 2.385 1.015 2.625 ;
        RECT 1.015 2.395 1.025 2.635 ;
        RECT 1.025 2.405 1.035 2.645 ;
        RECT 1.035 2.415 1.045 2.655 ;
        RECT 1.045 2.425 1.055 2.665 ;
        RECT 1.055 2.435 1.065 2.675 ;
        RECT 1.065 2.445 1.075 2.685 ;
        RECT 1.075 2.450 1.081 2.694 ;
        RECT 0.835 1.520 0.845 2.454 ;
        RECT 0.845 1.520 0.855 2.464 ;
        RECT 0.855 1.520 0.865 2.474 ;
        RECT 0.865 1.520 0.875 2.484 ;
        RECT 0.875 1.520 0.885 2.494 ;
        RECT 0.885 1.520 0.895 2.504 ;
        RECT 0.895 1.520 0.905 2.514 ;
        RECT 0.905 1.520 0.915 2.524 ;
        RECT 0.915 1.520 0.925 2.534 ;
        RECT 0.925 1.520 0.935 2.544 ;
        RECT 0.935 1.520 0.945 2.554 ;
        RECT 0.945 1.520 0.955 2.564 ;
        RECT 0.955 1.520 0.965 2.574 ;
        RECT 0.965 1.520 0.975 2.584 ;
        RECT 0.975 1.520 0.985 2.594 ;
        RECT 0.985 1.520 0.995 2.604 ;
        RECT 0.995 1.520 1.005 2.614 ;
        RECT 1.630 1.125 1.930 1.295 ;
        RECT 1.760 1.125 1.930 2.215 ;
        RECT 1.630 2.045 1.930 2.215 ;
        RECT 2.615 0.620 2.785 1.810 ;
        RECT 1.760 1.640 2.785 1.810 ;
        RECT 3.745 0.620 3.945 0.945 ;
        RECT 2.615 0.620 3.945 0.790 ;
        RECT 4.905 0.500 5.075 0.945 ;
        RECT 3.745 0.775 5.075 0.945 ;
        RECT 3.745 1.125 3.915 2.390 ;
        RECT 3.540 1.125 5.840 1.295 ;
        RECT 5.960 0.485 6.195 0.785 ;
        RECT 4.325 1.495 6.195 1.665 ;
        RECT 5.830 2.045 6.195 2.215 ;
        RECT 6.025 0.485 6.195 2.630 ;
        RECT 7.100 1.520 7.270 2.630 ;
        RECT 6.025 2.460 7.270 2.630 ;
  END 
END LATNSHDMXHT

MACRO LATNSHDLXHT
  CLASS  CORE ;
  FOREIGN LATNSHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.790 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 6.410 1.060 6.580 2.280 ;
        RECT 6.410 1.660 6.895 2.025 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.520 3.000 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.450 1.060 7.620 2.430 ;
        RECT 7.450 2.045 7.690 2.430 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.315 2.480 4.615 3.095 ;
        RECT 4.315 2.480 4.820 2.840 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.570 -0.300 0.870 0.825 ;
        RECT 2.385 -0.300 2.555 1.160 ;
        RECT 4.400 -0.300 4.700 0.595 ;
        RECT 5.375 -0.300 5.675 0.805 ;
        RECT 6.865 -0.300 7.165 1.295 ;
        RECT 0.000 -0.300 7.790 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.645 0.510 2.070 0.940 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.755 2.765 0.925 3.990 ;
        RECT 2.085 3.095 2.385 3.990 ;
        RECT 5.190 2.315 5.490 3.990 ;
        RECT 6.835 2.810 7.135 3.990 ;
        RECT 0.000 3.390 7.790 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 3.085 1.060 3.255 2.215 ;
        RECT 3.070 2.045 3.370 2.215 ;
        RECT 1.385 0.480 1.460 0.780 ;
        RECT 1.575 2.395 3.055 2.565 ;
        RECT 3.295 2.560 3.650 2.730 ;
        RECT 3.220 2.495 3.230 2.729 ;
        RECT 3.230 2.505 3.240 2.729 ;
        RECT 3.240 2.515 3.250 2.729 ;
        RECT 3.250 2.525 3.260 2.729 ;
        RECT 3.260 2.535 3.270 2.729 ;
        RECT 3.270 2.545 3.280 2.729 ;
        RECT 3.280 2.555 3.290 2.729 ;
        RECT 3.290 2.560 3.296 2.730 ;
        RECT 3.130 2.405 3.140 2.639 ;
        RECT 3.140 2.415 3.150 2.649 ;
        RECT 3.150 2.425 3.160 2.659 ;
        RECT 3.160 2.435 3.170 2.669 ;
        RECT 3.170 2.445 3.180 2.679 ;
        RECT 3.180 2.455 3.190 2.689 ;
        RECT 3.190 2.465 3.200 2.699 ;
        RECT 3.200 2.475 3.210 2.709 ;
        RECT 3.210 2.485 3.220 2.719 ;
        RECT 3.055 2.395 3.065 2.565 ;
        RECT 3.065 2.395 3.075 2.575 ;
        RECT 3.075 2.395 3.085 2.585 ;
        RECT 3.085 2.395 3.095 2.595 ;
        RECT 3.095 2.395 3.105 2.605 ;
        RECT 3.105 2.395 3.115 2.615 ;
        RECT 3.115 2.395 3.125 2.625 ;
        RECT 3.125 2.395 3.131 2.635 ;
        RECT 1.495 2.325 1.505 2.565 ;
        RECT 1.505 2.335 1.515 2.565 ;
        RECT 1.515 2.345 1.525 2.565 ;
        RECT 1.525 2.355 1.535 2.565 ;
        RECT 1.535 2.365 1.545 2.565 ;
        RECT 1.545 2.375 1.555 2.565 ;
        RECT 1.555 2.385 1.565 2.565 ;
        RECT 1.565 2.395 1.575 2.565 ;
        RECT 1.385 2.215 1.395 2.455 ;
        RECT 1.395 2.225 1.405 2.465 ;
        RECT 1.405 2.235 1.415 2.475 ;
        RECT 1.415 2.245 1.425 2.485 ;
        RECT 1.425 2.255 1.435 2.495 ;
        RECT 1.435 2.265 1.445 2.505 ;
        RECT 1.445 2.275 1.455 2.515 ;
        RECT 1.455 2.285 1.465 2.525 ;
        RECT 1.465 2.295 1.475 2.535 ;
        RECT 1.475 2.305 1.485 2.545 ;
        RECT 1.485 2.315 1.495 2.555 ;
        RECT 1.210 0.480 1.220 2.280 ;
        RECT 1.220 0.480 1.230 2.290 ;
        RECT 1.230 0.480 1.240 2.300 ;
        RECT 1.240 0.480 1.250 2.310 ;
        RECT 1.250 0.480 1.260 2.320 ;
        RECT 1.260 0.480 1.270 2.330 ;
        RECT 1.270 0.480 1.280 2.340 ;
        RECT 1.280 0.480 1.290 2.350 ;
        RECT 1.290 0.480 1.300 2.360 ;
        RECT 1.300 0.480 1.310 2.370 ;
        RECT 1.310 0.480 1.320 2.380 ;
        RECT 1.320 0.480 1.330 2.390 ;
        RECT 1.330 0.480 1.340 2.400 ;
        RECT 1.340 0.480 1.350 2.410 ;
        RECT 1.350 0.480 1.360 2.420 ;
        RECT 1.360 0.480 1.370 2.430 ;
        RECT 1.370 0.480 1.380 2.440 ;
        RECT 1.380 0.480 1.386 2.450 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.520 0.860 1.690 ;
        RECT 2.685 2.745 2.855 3.080 ;
        RECT 1.275 2.745 2.855 2.915 ;
        RECT 3.895 2.540 4.065 3.080 ;
        RECT 2.685 2.910 4.065 3.080 ;
        RECT 1.105 2.445 1.115 2.915 ;
        RECT 1.115 2.455 1.125 2.915 ;
        RECT 1.125 2.465 1.135 2.915 ;
        RECT 1.135 2.475 1.145 2.915 ;
        RECT 1.145 2.485 1.155 2.915 ;
        RECT 1.155 2.495 1.165 2.915 ;
        RECT 1.165 2.505 1.175 2.915 ;
        RECT 1.175 2.515 1.185 2.915 ;
        RECT 1.185 2.525 1.195 2.915 ;
        RECT 1.195 2.535 1.205 2.915 ;
        RECT 1.205 2.545 1.215 2.915 ;
        RECT 1.215 2.555 1.225 2.915 ;
        RECT 1.225 2.565 1.235 2.915 ;
        RECT 1.235 2.575 1.245 2.915 ;
        RECT 1.245 2.585 1.255 2.915 ;
        RECT 1.255 2.595 1.265 2.915 ;
        RECT 1.265 2.605 1.275 2.915 ;
        RECT 1.030 2.370 1.040 2.610 ;
        RECT 1.040 2.380 1.050 2.620 ;
        RECT 1.050 2.390 1.060 2.630 ;
        RECT 1.060 2.400 1.070 2.640 ;
        RECT 1.070 2.410 1.080 2.650 ;
        RECT 1.080 2.420 1.090 2.660 ;
        RECT 1.090 2.430 1.100 2.670 ;
        RECT 1.100 2.435 1.106 2.679 ;
        RECT 0.860 1.520 0.870 2.440 ;
        RECT 0.870 1.520 0.880 2.450 ;
        RECT 0.880 1.520 0.890 2.460 ;
        RECT 0.890 1.520 0.900 2.470 ;
        RECT 0.900 1.520 0.910 2.480 ;
        RECT 0.910 1.520 0.920 2.490 ;
        RECT 0.920 1.520 0.930 2.500 ;
        RECT 0.930 1.520 0.940 2.510 ;
        RECT 0.940 1.520 0.950 2.520 ;
        RECT 0.950 1.520 0.960 2.530 ;
        RECT 0.960 1.520 0.970 2.540 ;
        RECT 0.970 1.520 0.980 2.550 ;
        RECT 0.980 1.520 0.990 2.560 ;
        RECT 0.990 1.520 1.000 2.570 ;
        RECT 1.000 1.520 1.010 2.580 ;
        RECT 1.010 1.520 1.020 2.590 ;
        RECT 1.020 1.520 1.030 2.600 ;
        RECT 1.655 1.125 1.955 1.295 ;
        RECT 1.785 1.125 1.955 2.215 ;
        RECT 1.655 2.045 1.955 2.215 ;
        RECT 2.735 0.710 2.905 1.795 ;
        RECT 1.785 1.625 2.905 1.795 ;
        RECT 3.695 0.710 3.930 0.945 ;
        RECT 2.735 0.710 3.930 0.880 ;
        RECT 4.905 0.500 5.075 0.945 ;
        RECT 3.695 0.775 5.075 0.945 ;
        RECT 3.605 1.125 3.775 2.280 ;
        RECT 3.605 1.980 3.825 2.280 ;
        RECT 3.540 1.125 5.840 1.295 ;
        RECT 5.960 0.570 6.190 0.870 ;
        RECT 4.265 1.585 6.190 1.755 ;
        RECT 5.830 2.045 6.190 2.215 ;
        RECT 6.020 0.570 6.190 2.630 ;
        RECT 7.100 1.520 7.270 2.630 ;
        RECT 6.020 2.460 7.270 2.630 ;
  END 
END LATNSHDLXHT

MACRO LATNSHD2XHT
  CLASS  CORE ;
  FOREIGN LATNSHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.020 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.010 0.720 7.180 2.280 ;
        RECT 7.010 1.670 7.280 2.020 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.520 3.040 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.050 0.720 8.220 2.960 ;
        RECT 8.050 1.260 8.510 1.610 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.350 2.950 4.890 3.210 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.715 ;
        RECT 2.315 -0.300 2.485 1.360 ;
        RECT 4.585 -0.300 4.885 0.595 ;
        RECT 6.420 -0.300 6.720 1.055 ;
        RECT 7.465 -0.300 7.765 1.060 ;
        RECT 8.505 -0.300 8.805 1.055 ;
        RECT 0.000 -0.300 9.020 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.645 0.510 2.070 0.895 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 2.820 0.890 3.990 ;
        RECT 2.025 3.095 2.325 3.990 ;
        RECT 5.150 2.295 5.450 3.990 ;
        RECT 6.425 2.975 6.725 3.990 ;
        RECT 7.465 2.975 7.765 3.990 ;
        RECT 8.505 2.295 8.805 3.990 ;
        RECT 0.000 3.390 9.020 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 3.040 1.060 3.210 2.420 ;
        RECT 1.500 2.395 2.560 2.565 ;
        RECT 3.390 1.750 3.560 2.775 ;
        RECT 2.845 2.605 3.560 2.775 ;
        RECT 2.770 2.540 2.780 2.774 ;
        RECT 2.780 2.550 2.790 2.774 ;
        RECT 2.790 2.560 2.800 2.774 ;
        RECT 2.800 2.570 2.810 2.774 ;
        RECT 2.810 2.580 2.820 2.774 ;
        RECT 2.820 2.590 2.830 2.774 ;
        RECT 2.830 2.600 2.840 2.774 ;
        RECT 2.840 2.605 2.846 2.775 ;
        RECT 2.635 2.405 2.645 2.639 ;
        RECT 2.645 2.415 2.655 2.649 ;
        RECT 2.655 2.425 2.665 2.659 ;
        RECT 2.665 2.435 2.675 2.669 ;
        RECT 2.675 2.445 2.685 2.679 ;
        RECT 2.685 2.455 2.695 2.689 ;
        RECT 2.695 2.465 2.705 2.699 ;
        RECT 2.705 2.475 2.715 2.709 ;
        RECT 2.715 2.485 2.725 2.719 ;
        RECT 2.725 2.495 2.735 2.729 ;
        RECT 2.735 2.505 2.745 2.739 ;
        RECT 2.745 2.515 2.755 2.749 ;
        RECT 2.755 2.525 2.765 2.759 ;
        RECT 2.765 2.530 2.771 2.770 ;
        RECT 2.560 2.395 2.570 2.565 ;
        RECT 2.570 2.395 2.580 2.575 ;
        RECT 2.580 2.395 2.590 2.585 ;
        RECT 2.590 2.395 2.600 2.595 ;
        RECT 2.600 2.395 2.610 2.605 ;
        RECT 2.610 2.395 2.620 2.615 ;
        RECT 2.620 2.395 2.630 2.625 ;
        RECT 2.630 2.395 2.636 2.635 ;
        RECT 1.420 2.325 1.430 2.565 ;
        RECT 1.430 2.335 1.440 2.565 ;
        RECT 1.440 2.345 1.450 2.565 ;
        RECT 1.450 2.355 1.460 2.565 ;
        RECT 1.460 2.365 1.470 2.565 ;
        RECT 1.470 2.375 1.480 2.565 ;
        RECT 1.480 2.385 1.490 2.565 ;
        RECT 1.490 2.395 1.500 2.565 ;
        RECT 1.385 2.290 1.395 2.530 ;
        RECT 1.395 2.300 1.405 2.540 ;
        RECT 1.405 2.310 1.415 2.550 ;
        RECT 1.415 2.315 1.421 2.559 ;
        RECT 1.210 1.060 1.220 2.354 ;
        RECT 1.220 1.060 1.230 2.364 ;
        RECT 1.230 1.060 1.240 2.374 ;
        RECT 1.240 1.060 1.250 2.384 ;
        RECT 1.250 1.060 1.260 2.394 ;
        RECT 1.260 1.060 1.270 2.404 ;
        RECT 1.270 1.060 1.280 2.414 ;
        RECT 1.280 1.060 1.290 2.424 ;
        RECT 1.290 1.060 1.300 2.434 ;
        RECT 1.300 1.060 1.310 2.444 ;
        RECT 1.310 1.060 1.320 2.454 ;
        RECT 1.320 1.060 1.330 2.464 ;
        RECT 1.330 1.060 1.340 2.474 ;
        RECT 1.340 1.060 1.350 2.484 ;
        RECT 1.350 1.060 1.360 2.494 ;
        RECT 1.360 1.060 1.370 2.504 ;
        RECT 1.370 1.060 1.380 2.514 ;
        RECT 1.380 1.060 1.386 2.524 ;
        RECT 1.150 1.980 1.160 2.294 ;
        RECT 1.160 1.980 1.170 2.304 ;
        RECT 1.170 1.980 1.180 2.314 ;
        RECT 1.180 1.980 1.190 2.324 ;
        RECT 1.190 1.980 1.200 2.334 ;
        RECT 1.200 1.980 1.210 2.344 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.520 0.800 1.690 ;
        RECT 0.970 1.520 1.030 1.820 ;
        RECT 1.240 2.745 2.405 2.915 ;
        RECT 3.935 2.685 4.105 3.125 ;
        RECT 2.690 2.955 4.105 3.125 ;
        RECT 2.615 2.890 2.625 3.124 ;
        RECT 2.625 2.900 2.635 3.124 ;
        RECT 2.635 2.910 2.645 3.124 ;
        RECT 2.645 2.920 2.655 3.124 ;
        RECT 2.655 2.930 2.665 3.124 ;
        RECT 2.665 2.940 2.675 3.124 ;
        RECT 2.675 2.950 2.685 3.124 ;
        RECT 2.685 2.955 2.691 3.125 ;
        RECT 2.480 2.755 2.490 2.989 ;
        RECT 2.490 2.765 2.500 2.999 ;
        RECT 2.500 2.775 2.510 3.009 ;
        RECT 2.510 2.785 2.520 3.019 ;
        RECT 2.520 2.795 2.530 3.029 ;
        RECT 2.530 2.805 2.540 3.039 ;
        RECT 2.540 2.815 2.550 3.049 ;
        RECT 2.550 2.825 2.560 3.059 ;
        RECT 2.560 2.835 2.570 3.069 ;
        RECT 2.570 2.845 2.580 3.079 ;
        RECT 2.580 2.855 2.590 3.089 ;
        RECT 2.590 2.865 2.600 3.099 ;
        RECT 2.600 2.875 2.610 3.109 ;
        RECT 2.610 2.880 2.616 3.120 ;
        RECT 2.405 2.745 2.415 2.915 ;
        RECT 2.415 2.745 2.425 2.925 ;
        RECT 2.425 2.745 2.435 2.935 ;
        RECT 2.435 2.745 2.445 2.945 ;
        RECT 2.445 2.745 2.455 2.955 ;
        RECT 2.455 2.745 2.465 2.965 ;
        RECT 2.465 2.745 2.475 2.975 ;
        RECT 2.475 2.745 2.481 2.985 ;
        RECT 1.070 2.480 1.080 2.914 ;
        RECT 1.080 2.490 1.090 2.914 ;
        RECT 1.090 2.500 1.100 2.914 ;
        RECT 1.100 2.510 1.110 2.914 ;
        RECT 1.110 2.520 1.120 2.914 ;
        RECT 1.120 2.530 1.130 2.914 ;
        RECT 1.130 2.540 1.140 2.914 ;
        RECT 1.140 2.550 1.150 2.914 ;
        RECT 1.150 2.560 1.160 2.914 ;
        RECT 1.160 2.570 1.170 2.914 ;
        RECT 1.170 2.580 1.180 2.914 ;
        RECT 1.180 2.590 1.190 2.914 ;
        RECT 1.190 2.600 1.200 2.914 ;
        RECT 1.200 2.610 1.210 2.914 ;
        RECT 1.210 2.620 1.220 2.914 ;
        RECT 1.220 2.630 1.230 2.914 ;
        RECT 1.230 2.640 1.240 2.914 ;
        RECT 0.970 2.380 0.980 2.630 ;
        RECT 0.980 2.390 0.990 2.640 ;
        RECT 0.990 2.400 1.000 2.650 ;
        RECT 1.000 2.410 1.010 2.660 ;
        RECT 1.010 2.420 1.020 2.670 ;
        RECT 1.020 2.430 1.030 2.680 ;
        RECT 1.030 2.440 1.040 2.690 ;
        RECT 1.040 2.450 1.050 2.700 ;
        RECT 1.050 2.460 1.060 2.710 ;
        RECT 1.060 2.470 1.070 2.720 ;
        RECT 0.800 1.520 0.810 2.460 ;
        RECT 0.810 1.520 0.820 2.470 ;
        RECT 0.820 1.520 0.830 2.480 ;
        RECT 0.830 1.520 0.840 2.490 ;
        RECT 0.840 1.520 0.850 2.500 ;
        RECT 0.850 1.520 0.860 2.510 ;
        RECT 0.860 1.520 0.870 2.520 ;
        RECT 0.870 1.520 0.880 2.530 ;
        RECT 0.880 1.520 0.890 2.540 ;
        RECT 0.890 1.520 0.900 2.550 ;
        RECT 0.900 1.520 0.910 2.560 ;
        RECT 0.910 1.520 0.920 2.570 ;
        RECT 0.920 1.520 0.930 2.580 ;
        RECT 0.930 1.520 0.940 2.590 ;
        RECT 0.940 1.520 0.950 2.600 ;
        RECT 0.950 1.520 0.960 2.610 ;
        RECT 0.960 1.520 0.970 2.620 ;
        RECT 1.655 1.125 1.955 1.295 ;
        RECT 1.785 1.125 1.955 2.215 ;
        RECT 1.595 2.045 1.955 2.215 ;
        RECT 2.665 0.710 2.835 1.805 ;
        RECT 1.785 1.635 2.835 1.805 ;
        RECT 3.780 0.710 3.960 0.945 ;
        RECT 2.665 0.710 3.960 0.880 ;
        RECT 5.495 0.585 5.665 0.945 ;
        RECT 3.780 0.775 5.665 0.945 ;
        RECT 3.540 1.125 3.910 1.300 ;
        RECT 3.740 1.125 3.910 2.420 ;
        RECT 3.540 1.125 5.515 1.295 ;
        RECT 5.345 1.125 5.515 1.665 ;
        RECT 5.345 1.495 5.800 1.665 ;
        RECT 4.400 1.520 4.570 2.015 ;
        RECT 5.935 1.060 6.150 1.360 ;
        RECT 4.400 1.845 6.150 2.015 ;
        RECT 5.980 1.060 6.150 2.630 ;
        RECT 7.670 1.520 7.840 2.630 ;
        RECT 5.980 2.460 7.840 2.630 ;
  END 
END LATNSHD2XHT

MACRO LATNSHD1XHT
  CLASS  CORE ;
  FOREIGN LATNSHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.790 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 6.410 1.060 6.580 2.280 ;
        RECT 6.410 1.660 6.895 2.025 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.545 3.000 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.450 0.720 7.645 2.960 ;
        RECT 7.450 2.455 7.690 2.960 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.445 2.480 4.615 3.210 ;
        RECT 4.315 3.040 4.615 3.210 ;
        RECT 4.445 2.480 4.820 2.840 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.715 ;
        RECT 2.385 -0.300 2.555 1.020 ;
        RECT 4.400 -0.300 4.700 0.595 ;
        RECT 5.375 -0.300 5.675 0.720 ;
        RECT 6.865 -0.300 7.165 1.055 ;
        RECT 0.000 -0.300 7.790 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.645 0.510 2.135 0.895 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.755 2.855 0.925 3.990 ;
        RECT 2.085 3.095 2.385 3.990 ;
        RECT 5.235 2.405 5.535 3.990 ;
        RECT 6.865 2.975 7.165 3.990 ;
        RECT 0.000 3.390 7.790 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 3.085 1.060 3.255 2.215 ;
        RECT 3.070 2.045 3.370 2.215 ;
        RECT 1.385 0.480 1.460 0.780 ;
        RECT 1.525 2.395 3.475 2.565 ;
        RECT 3.305 2.395 3.475 2.840 ;
        RECT 3.305 2.670 3.650 2.840 ;
        RECT 1.445 2.325 1.455 2.565 ;
        RECT 1.455 2.335 1.465 2.565 ;
        RECT 1.465 2.345 1.475 2.565 ;
        RECT 1.475 2.355 1.485 2.565 ;
        RECT 1.485 2.365 1.495 2.565 ;
        RECT 1.495 2.375 1.505 2.565 ;
        RECT 1.505 2.385 1.515 2.565 ;
        RECT 1.515 2.395 1.525 2.565 ;
        RECT 1.385 2.265 1.395 2.505 ;
        RECT 1.395 2.275 1.405 2.515 ;
        RECT 1.405 2.285 1.415 2.525 ;
        RECT 1.415 2.295 1.425 2.535 ;
        RECT 1.425 2.305 1.435 2.545 ;
        RECT 1.435 2.315 1.445 2.555 ;
        RECT 1.210 0.480 1.220 2.330 ;
        RECT 1.220 0.480 1.230 2.340 ;
        RECT 1.230 0.480 1.240 2.350 ;
        RECT 1.240 0.480 1.250 2.360 ;
        RECT 1.250 0.480 1.260 2.370 ;
        RECT 1.260 0.480 1.270 2.380 ;
        RECT 1.270 0.480 1.280 2.390 ;
        RECT 1.280 0.480 1.290 2.400 ;
        RECT 1.290 0.480 1.300 2.410 ;
        RECT 1.300 0.480 1.310 2.420 ;
        RECT 1.310 0.480 1.320 2.430 ;
        RECT 1.320 0.480 1.330 2.440 ;
        RECT 1.330 0.480 1.340 2.450 ;
        RECT 1.340 0.480 1.350 2.460 ;
        RECT 1.350 0.480 1.360 2.470 ;
        RECT 1.360 0.480 1.370 2.480 ;
        RECT 1.370 0.480 1.380 2.490 ;
        RECT 1.380 0.480 1.386 2.500 ;
        RECT 0.195 1.060 0.365 2.280 ;
        RECT 0.195 1.520 0.860 1.690 ;
        RECT 1.275 2.745 2.955 2.915 ;
        RECT 3.830 2.685 4.000 3.190 ;
        RECT 3.230 3.020 4.000 3.190 ;
        RECT 3.830 2.685 4.130 2.855 ;
        RECT 3.145 2.945 3.155 3.189 ;
        RECT 3.155 2.955 3.165 3.189 ;
        RECT 3.165 2.965 3.175 3.189 ;
        RECT 3.175 2.975 3.185 3.189 ;
        RECT 3.185 2.985 3.195 3.189 ;
        RECT 3.195 2.995 3.205 3.189 ;
        RECT 3.205 3.005 3.215 3.189 ;
        RECT 3.215 3.015 3.225 3.189 ;
        RECT 3.225 3.020 3.231 3.190 ;
        RECT 3.125 2.925 3.135 3.169 ;
        RECT 3.135 2.935 3.145 3.179 ;
        RECT 2.955 2.745 2.965 2.999 ;
        RECT 2.965 2.745 2.975 3.009 ;
        RECT 2.975 2.745 2.985 3.019 ;
        RECT 2.985 2.745 2.995 3.029 ;
        RECT 2.995 2.745 3.005 3.039 ;
        RECT 3.005 2.745 3.015 3.049 ;
        RECT 3.015 2.745 3.025 3.059 ;
        RECT 3.025 2.745 3.035 3.069 ;
        RECT 3.035 2.745 3.045 3.079 ;
        RECT 3.045 2.745 3.055 3.089 ;
        RECT 3.055 2.745 3.065 3.099 ;
        RECT 3.065 2.745 3.075 3.109 ;
        RECT 3.075 2.745 3.085 3.119 ;
        RECT 3.085 2.745 3.095 3.129 ;
        RECT 3.095 2.745 3.105 3.139 ;
        RECT 3.105 2.745 3.115 3.149 ;
        RECT 3.115 2.745 3.125 3.159 ;
        RECT 1.105 2.490 1.115 2.914 ;
        RECT 1.115 2.500 1.125 2.914 ;
        RECT 1.125 2.510 1.135 2.914 ;
        RECT 1.135 2.520 1.145 2.914 ;
        RECT 1.145 2.530 1.155 2.914 ;
        RECT 1.155 2.540 1.165 2.914 ;
        RECT 1.165 2.550 1.175 2.914 ;
        RECT 1.175 2.560 1.185 2.914 ;
        RECT 1.185 2.570 1.195 2.914 ;
        RECT 1.195 2.580 1.205 2.914 ;
        RECT 1.205 2.590 1.215 2.914 ;
        RECT 1.215 2.600 1.225 2.914 ;
        RECT 1.225 2.610 1.235 2.914 ;
        RECT 1.235 2.620 1.245 2.914 ;
        RECT 1.245 2.630 1.255 2.914 ;
        RECT 1.255 2.640 1.265 2.914 ;
        RECT 1.265 2.650 1.275 2.914 ;
        RECT 1.030 2.415 1.040 2.649 ;
        RECT 1.040 2.425 1.050 2.659 ;
        RECT 1.050 2.435 1.060 2.669 ;
        RECT 1.060 2.445 1.070 2.679 ;
        RECT 1.070 2.455 1.080 2.689 ;
        RECT 1.080 2.465 1.090 2.699 ;
        RECT 1.090 2.475 1.100 2.709 ;
        RECT 1.100 2.480 1.106 2.720 ;
        RECT 0.860 1.520 0.870 2.480 ;
        RECT 0.870 1.520 0.880 2.490 ;
        RECT 0.880 1.520 0.890 2.500 ;
        RECT 0.890 1.520 0.900 2.510 ;
        RECT 0.900 1.520 0.910 2.520 ;
        RECT 0.910 1.520 0.920 2.530 ;
        RECT 0.920 1.520 0.930 2.540 ;
        RECT 0.930 1.520 0.940 2.550 ;
        RECT 0.940 1.520 0.950 2.560 ;
        RECT 0.950 1.520 0.960 2.570 ;
        RECT 0.960 1.520 0.970 2.580 ;
        RECT 0.970 1.520 0.980 2.590 ;
        RECT 0.980 1.520 0.990 2.600 ;
        RECT 0.990 1.520 1.000 2.610 ;
        RECT 1.000 1.520 1.010 2.620 ;
        RECT 1.010 1.520 1.020 2.630 ;
        RECT 1.020 1.520 1.030 2.640 ;
        RECT 1.655 1.125 1.955 1.295 ;
        RECT 1.785 1.125 1.955 2.215 ;
        RECT 1.655 2.045 1.955 2.215 ;
        RECT 2.735 0.710 2.905 1.835 ;
        RECT 1.785 1.665 2.905 1.835 ;
        RECT 3.765 0.710 4.020 0.945 ;
        RECT 2.735 0.710 4.020 0.880 ;
        RECT 4.905 0.500 5.075 0.945 ;
        RECT 3.765 0.775 5.075 0.945 ;
        RECT 3.655 1.125 3.825 2.280 ;
        RECT 3.540 1.125 5.840 1.295 ;
        RECT 5.960 0.485 6.190 0.785 ;
        RECT 4.265 1.585 6.190 1.755 ;
        RECT 5.830 2.045 6.190 2.215 ;
        RECT 6.020 0.485 6.190 2.630 ;
        RECT 7.100 1.520 7.270 2.630 ;
        RECT 6.020 2.460 7.270 2.630 ;
  END 
END LATNSHD1XHT

MACRO LATNRHDMXHT
  CLASS  CORE ;
  FOREIGN LATNRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.380 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.840 0.840 6.170 1.200 ;
        RECT 6.000 0.840 6.170 2.280 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.465 0.520 2.950 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.040 1.060 7.210 2.280 ;
        RECT 7.040 1.260 7.280 1.610 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.595 2.090 2.135 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.360 0.645 1.530 0.945 ;
        RECT 2.080 0.575 2.250 0.945 ;
        RECT 1.360 0.775 2.250 0.945 ;
        RECT 2.080 0.575 4.570 0.745 ;
        RECT 4.400 0.575 4.570 1.800 ;
        RECT 4.400 1.330 4.615 1.800 ;
        RECT 4.400 1.330 4.900 1.540 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.745 ;
        RECT 1.730 -0.300 1.900 0.575 ;
        RECT 4.750 -0.300 5.050 1.095 ;
        RECT 6.455 -0.300 6.755 1.145 ;
        RECT 0.000 -0.300 7.380 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.730 2.830 0.900 3.990 ;
        RECT 1.625 3.095 1.925 3.990 ;
        RECT 4.010 2.395 4.310 3.990 ;
        RECT 4.980 2.745 5.280 3.990 ;
        RECT 6.485 2.925 6.785 3.990 ;
        RECT 0.000 3.390 7.380 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 0.860 1.755 ;
        RECT 1.250 2.745 2.435 2.915 ;
        RECT 2.265 2.745 2.435 3.205 ;
        RECT 2.265 3.035 2.755 3.205 ;
        RECT 1.080 2.425 1.090 2.915 ;
        RECT 1.090 2.435 1.100 2.915 ;
        RECT 1.100 2.445 1.110 2.915 ;
        RECT 1.110 2.455 1.120 2.915 ;
        RECT 1.120 2.465 1.130 2.915 ;
        RECT 1.130 2.475 1.140 2.915 ;
        RECT 1.140 2.485 1.150 2.915 ;
        RECT 1.150 2.495 1.160 2.915 ;
        RECT 1.160 2.505 1.170 2.915 ;
        RECT 1.170 2.515 1.180 2.915 ;
        RECT 1.180 2.525 1.190 2.915 ;
        RECT 1.190 2.535 1.200 2.915 ;
        RECT 1.200 2.545 1.210 2.915 ;
        RECT 1.210 2.555 1.220 2.915 ;
        RECT 1.220 2.565 1.230 2.915 ;
        RECT 1.230 2.575 1.240 2.915 ;
        RECT 1.240 2.585 1.250 2.915 ;
        RECT 1.030 2.375 1.040 2.619 ;
        RECT 1.040 2.385 1.050 2.629 ;
        RECT 1.050 2.395 1.060 2.639 ;
        RECT 1.060 2.405 1.070 2.649 ;
        RECT 1.070 2.415 1.080 2.659 ;
        RECT 0.860 1.520 0.870 2.450 ;
        RECT 0.870 1.520 0.880 2.460 ;
        RECT 0.880 1.520 0.890 2.470 ;
        RECT 0.890 1.520 0.900 2.480 ;
        RECT 0.900 1.520 0.910 2.490 ;
        RECT 0.910 1.520 0.920 2.500 ;
        RECT 0.920 1.520 0.930 2.510 ;
        RECT 0.930 1.520 0.940 2.520 ;
        RECT 0.940 1.520 0.950 2.530 ;
        RECT 0.950 1.520 0.960 2.540 ;
        RECT 0.960 1.520 0.970 2.550 ;
        RECT 0.970 1.520 0.980 2.560 ;
        RECT 0.980 1.520 0.990 2.570 ;
        RECT 0.990 1.520 1.000 2.580 ;
        RECT 1.000 1.520 1.010 2.590 ;
        RECT 1.010 1.520 1.020 2.600 ;
        RECT 1.020 1.520 1.030 2.610 ;
        RECT 2.445 0.925 2.615 2.215 ;
        RECT 2.315 2.045 2.615 2.215 ;
        RECT 2.445 0.925 2.945 1.095 ;
        RECT 1.085 1.125 1.210 1.295 ;
        RECT 2.805 1.345 2.975 2.715 ;
        RECT 1.565 2.395 2.975 2.565 ;
        RECT 2.805 2.540 3.175 2.715 ;
        RECT 3.005 2.540 3.175 2.950 ;
        RECT 2.805 1.345 3.830 1.515 ;
        RECT 1.490 2.330 1.500 2.564 ;
        RECT 1.500 2.340 1.510 2.564 ;
        RECT 1.510 2.350 1.520 2.564 ;
        RECT 1.520 2.360 1.530 2.564 ;
        RECT 1.530 2.370 1.540 2.564 ;
        RECT 1.540 2.380 1.550 2.564 ;
        RECT 1.550 2.390 1.560 2.564 ;
        RECT 1.560 2.395 1.566 2.565 ;
        RECT 1.385 2.225 1.395 2.459 ;
        RECT 1.395 2.235 1.405 2.469 ;
        RECT 1.405 2.245 1.415 2.479 ;
        RECT 1.415 2.255 1.425 2.489 ;
        RECT 1.425 2.265 1.435 2.499 ;
        RECT 1.435 2.275 1.445 2.509 ;
        RECT 1.445 2.285 1.455 2.519 ;
        RECT 1.455 2.295 1.465 2.529 ;
        RECT 1.465 2.305 1.475 2.539 ;
        RECT 1.475 2.315 1.485 2.549 ;
        RECT 1.485 2.320 1.491 2.560 ;
        RECT 1.210 1.125 1.220 2.285 ;
        RECT 1.220 1.125 1.230 2.295 ;
        RECT 1.230 1.125 1.240 2.305 ;
        RECT 1.240 1.125 1.250 2.315 ;
        RECT 1.250 1.125 1.260 2.325 ;
        RECT 1.260 1.125 1.270 2.335 ;
        RECT 1.270 1.125 1.280 2.345 ;
        RECT 1.280 1.125 1.290 2.355 ;
        RECT 1.290 1.125 1.300 2.365 ;
        RECT 1.300 1.125 1.310 2.375 ;
        RECT 1.310 1.125 1.320 2.385 ;
        RECT 1.320 1.125 1.330 2.395 ;
        RECT 1.330 1.125 1.340 2.405 ;
        RECT 1.340 1.125 1.350 2.415 ;
        RECT 1.350 1.125 1.360 2.425 ;
        RECT 1.360 1.125 1.370 2.435 ;
        RECT 1.370 1.125 1.380 2.445 ;
        RECT 1.380 1.125 1.386 2.455 ;
        RECT 3.155 1.980 3.325 2.280 ;
        RECT 3.155 2.045 3.330 2.280 ;
        RECT 3.165 0.925 4.220 1.095 ;
        RECT 4.050 0.925 4.220 2.215 ;
        RECT 5.060 1.730 5.360 2.215 ;
        RECT 3.155 2.045 5.360 2.215 ;
        RECT 4.630 2.395 4.800 3.175 ;
        RECT 4.500 3.005 4.800 3.175 ;
        RECT 5.345 0.860 5.515 1.550 ;
        RECT 5.345 1.380 5.735 1.550 ;
        RECT 4.630 2.395 5.735 2.565 ;
        RECT 5.565 1.380 5.735 2.860 ;
        RECT 6.660 1.540 6.830 2.630 ;
        RECT 5.565 2.460 6.830 2.630 ;
  END 
END LATNRHDMXHT

MACRO LATNRHDLXHT
  CLASS  CORE ;
  FOREIGN LATNRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.380 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.840 0.800 6.170 1.225 ;
        RECT 6.000 0.800 6.170 2.280 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.465 0.395 2.840 ;
        RECT 0.100 2.465 0.590 2.635 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.040 1.060 7.235 2.280 ;
        RECT 7.040 1.060 7.280 1.610 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.735 1.595 2.115 2.135 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.010 0.550 4.655 0.670 ;
        RECT 2.205 0.500 2.375 0.720 ;
        RECT 2.010 0.500 2.375 0.670 ;
        RECT 4.085 0.500 4.655 0.720 ;
        RECT 2.205 0.550 4.655 0.720 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.780 ;
        RECT 1.660 -0.300 1.830 1.040 ;
        RECT 1.660 0.870 1.995 1.040 ;
        RECT 4.840 -0.300 5.010 1.095 ;
        RECT 4.710 0.925 5.010 1.095 ;
        RECT 6.455 -0.300 6.755 1.295 ;
        RECT 0.000 -0.300 7.380 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.685 2.860 0.985 3.990 ;
        RECT 1.650 3.095 1.950 3.990 ;
        RECT 4.025 2.440 4.325 3.990 ;
        RECT 4.995 2.745 5.295 3.990 ;
        RECT 6.485 2.815 6.785 3.990 ;
        RECT 0.000 3.390 7.380 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.470 0.970 2.640 2.215 ;
        RECT 2.340 2.045 2.640 2.215 ;
        RECT 2.470 0.970 2.970 1.140 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 0.885 1.755 ;
        RECT 2.145 2.745 2.315 3.085 ;
        RECT 1.335 2.745 2.315 2.915 ;
        RECT 3.350 2.480 3.520 3.085 ;
        RECT 2.145 2.915 3.520 3.085 ;
        RECT 1.165 2.485 1.175 2.915 ;
        RECT 1.175 2.495 1.185 2.915 ;
        RECT 1.185 2.505 1.195 2.915 ;
        RECT 1.195 2.515 1.205 2.915 ;
        RECT 1.205 2.525 1.215 2.915 ;
        RECT 1.215 2.535 1.225 2.915 ;
        RECT 1.225 2.545 1.235 2.915 ;
        RECT 1.235 2.555 1.245 2.915 ;
        RECT 1.245 2.565 1.255 2.915 ;
        RECT 1.255 2.575 1.265 2.915 ;
        RECT 1.265 2.585 1.275 2.915 ;
        RECT 1.275 2.595 1.285 2.915 ;
        RECT 1.285 2.605 1.295 2.915 ;
        RECT 1.295 2.615 1.305 2.915 ;
        RECT 1.305 2.625 1.315 2.915 ;
        RECT 1.315 2.635 1.325 2.915 ;
        RECT 1.325 2.645 1.335 2.915 ;
        RECT 1.055 2.375 1.065 2.609 ;
        RECT 1.065 2.385 1.075 2.619 ;
        RECT 1.075 2.395 1.085 2.629 ;
        RECT 1.085 2.405 1.095 2.639 ;
        RECT 1.095 2.415 1.105 2.649 ;
        RECT 1.105 2.425 1.115 2.659 ;
        RECT 1.115 2.435 1.125 2.669 ;
        RECT 1.125 2.445 1.135 2.679 ;
        RECT 1.135 2.455 1.145 2.689 ;
        RECT 1.145 2.465 1.155 2.699 ;
        RECT 1.155 2.475 1.165 2.709 ;
        RECT 0.885 1.520 0.895 2.440 ;
        RECT 0.895 1.520 0.905 2.450 ;
        RECT 0.905 1.520 0.915 2.460 ;
        RECT 0.915 1.520 0.925 2.470 ;
        RECT 0.925 1.520 0.935 2.480 ;
        RECT 0.935 1.520 0.945 2.490 ;
        RECT 0.945 1.520 0.955 2.500 ;
        RECT 0.955 1.520 0.965 2.510 ;
        RECT 0.965 1.520 0.975 2.520 ;
        RECT 0.975 1.520 0.985 2.530 ;
        RECT 0.985 1.520 0.995 2.540 ;
        RECT 0.995 1.520 1.005 2.550 ;
        RECT 1.005 1.520 1.015 2.560 ;
        RECT 1.015 1.520 1.025 2.570 ;
        RECT 1.025 1.520 1.035 2.580 ;
        RECT 1.035 1.520 1.045 2.590 ;
        RECT 1.045 1.520 1.055 2.600 ;
        RECT 1.115 1.125 1.235 1.295 ;
        RECT 1.595 2.395 2.990 2.565 ;
        RECT 2.820 1.345 2.990 2.735 ;
        RECT 2.650 2.395 2.990 2.735 ;
        RECT 2.820 1.345 3.850 1.515 ;
        RECT 1.515 2.325 1.525 2.565 ;
        RECT 1.525 2.335 1.535 2.565 ;
        RECT 1.535 2.345 1.545 2.565 ;
        RECT 1.545 2.355 1.555 2.565 ;
        RECT 1.555 2.365 1.565 2.565 ;
        RECT 1.565 2.375 1.575 2.565 ;
        RECT 1.575 2.385 1.585 2.565 ;
        RECT 1.585 2.395 1.595 2.565 ;
        RECT 1.415 2.225 1.425 2.465 ;
        RECT 1.425 2.235 1.435 2.475 ;
        RECT 1.435 2.245 1.445 2.485 ;
        RECT 1.445 2.255 1.455 2.495 ;
        RECT 1.455 2.265 1.465 2.505 ;
        RECT 1.465 2.275 1.475 2.515 ;
        RECT 1.475 2.285 1.485 2.525 ;
        RECT 1.485 2.295 1.495 2.535 ;
        RECT 1.495 2.305 1.505 2.545 ;
        RECT 1.505 2.315 1.515 2.555 ;
        RECT 1.235 1.125 1.245 2.285 ;
        RECT 1.245 1.125 1.255 2.295 ;
        RECT 1.255 1.125 1.265 2.305 ;
        RECT 1.265 1.125 1.275 2.315 ;
        RECT 1.275 1.125 1.285 2.325 ;
        RECT 1.285 1.125 1.295 2.335 ;
        RECT 1.295 1.125 1.305 2.345 ;
        RECT 1.305 1.125 1.315 2.355 ;
        RECT 1.315 1.125 1.325 2.365 ;
        RECT 1.325 1.125 1.335 2.375 ;
        RECT 1.335 1.125 1.345 2.385 ;
        RECT 1.345 1.125 1.355 2.395 ;
        RECT 1.355 1.125 1.365 2.405 ;
        RECT 1.365 1.125 1.375 2.415 ;
        RECT 1.375 1.125 1.385 2.425 ;
        RECT 1.385 1.125 1.395 2.435 ;
        RECT 1.395 1.125 1.405 2.445 ;
        RECT 1.405 1.125 1.415 2.455 ;
        RECT 3.170 1.980 3.340 2.280 ;
        RECT 3.205 0.970 4.275 1.140 ;
        RECT 4.105 0.970 4.275 2.215 ;
        RECT 5.145 1.795 5.445 2.215 ;
        RECT 3.170 2.045 5.445 2.215 ;
        RECT 4.525 2.395 4.695 3.080 ;
        RECT 5.370 0.860 5.540 1.590 ;
        RECT 5.370 1.420 5.815 1.590 ;
        RECT 5.580 2.395 5.750 2.860 ;
        RECT 5.645 1.420 5.815 2.635 ;
        RECT 4.525 2.395 5.815 2.565 ;
        RECT 6.660 1.540 6.830 2.635 ;
        RECT 5.580 2.465 6.830 2.635 ;
  END 
END LATNRHDLXHT

MACRO LATNRHD2XHT
  CLASS  CORE ;
  FOREIGN LATNRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.610 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 6.660 0.845 6.880 1.195 ;
        RECT 6.710 0.720 6.880 2.280 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.520 2.950 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.750 0.720 7.920 2.960 ;
        RECT 7.750 1.635 8.100 2.035 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.595 2.110 2.120 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.375 0.645 1.545 0.945 ;
        RECT 2.100 0.550 2.270 0.945 ;
        RECT 1.375 0.775 2.270 0.945 ;
        RECT 2.100 0.550 4.610 0.720 ;
        RECT 4.440 0.550 4.610 1.820 ;
        RECT 4.440 1.330 4.925 1.540 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.715 ;
        RECT 1.745 -0.300 1.915 0.595 ;
        RECT 4.840 -0.300 5.010 1.060 ;
        RECT 6.125 -0.300 6.425 1.055 ;
        RECT 7.165 -0.300 7.465 1.055 ;
        RECT 8.205 -0.300 8.505 1.055 ;
        RECT 0.000 -0.300 8.610 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.730 2.830 0.900 3.990 ;
        RECT 1.515 3.050 1.815 3.990 ;
        RECT 4.005 2.975 4.305 3.990 ;
        RECT 5.095 2.755 5.395 3.990 ;
        RECT 6.125 2.975 6.425 3.990 ;
        RECT 7.165 2.975 7.465 3.990 ;
        RECT 8.205 2.295 8.505 3.990 ;
        RECT 0.000 3.390 8.610 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.520 0.860 1.690 ;
        RECT 1.250 2.700 1.895 2.870 ;
        RECT 2.315 3.040 2.665 3.210 ;
        RECT 2.235 2.970 2.245 3.210 ;
        RECT 2.245 2.980 2.255 3.210 ;
        RECT 2.255 2.990 2.265 3.210 ;
        RECT 2.265 3.000 2.275 3.210 ;
        RECT 2.275 3.010 2.285 3.210 ;
        RECT 2.285 3.020 2.295 3.210 ;
        RECT 2.295 3.030 2.305 3.210 ;
        RECT 2.305 3.040 2.315 3.210 ;
        RECT 1.975 2.710 1.985 2.950 ;
        RECT 1.985 2.720 1.995 2.960 ;
        RECT 1.995 2.730 2.005 2.970 ;
        RECT 2.005 2.740 2.015 2.980 ;
        RECT 2.015 2.750 2.025 2.990 ;
        RECT 2.025 2.760 2.035 3.000 ;
        RECT 2.035 2.770 2.045 3.010 ;
        RECT 2.045 2.780 2.055 3.020 ;
        RECT 2.055 2.790 2.065 3.030 ;
        RECT 2.065 2.800 2.075 3.040 ;
        RECT 2.075 2.810 2.085 3.050 ;
        RECT 2.085 2.820 2.095 3.060 ;
        RECT 2.095 2.830 2.105 3.070 ;
        RECT 2.105 2.840 2.115 3.080 ;
        RECT 2.115 2.850 2.125 3.090 ;
        RECT 2.125 2.860 2.135 3.100 ;
        RECT 2.135 2.870 2.145 3.110 ;
        RECT 2.145 2.880 2.155 3.120 ;
        RECT 2.155 2.890 2.165 3.130 ;
        RECT 2.165 2.900 2.175 3.140 ;
        RECT 2.175 2.910 2.185 3.150 ;
        RECT 2.185 2.920 2.195 3.160 ;
        RECT 2.195 2.930 2.205 3.170 ;
        RECT 2.205 2.940 2.215 3.180 ;
        RECT 2.215 2.950 2.225 3.190 ;
        RECT 2.225 2.960 2.235 3.200 ;
        RECT 1.895 2.700 1.905 2.870 ;
        RECT 1.905 2.700 1.915 2.880 ;
        RECT 1.915 2.700 1.925 2.890 ;
        RECT 1.925 2.700 1.935 2.900 ;
        RECT 1.935 2.700 1.945 2.910 ;
        RECT 1.945 2.700 1.955 2.920 ;
        RECT 1.955 2.700 1.965 2.930 ;
        RECT 1.965 2.700 1.975 2.940 ;
        RECT 1.080 2.415 1.090 2.869 ;
        RECT 1.090 2.425 1.100 2.869 ;
        RECT 1.100 2.435 1.110 2.869 ;
        RECT 1.110 2.445 1.120 2.869 ;
        RECT 1.120 2.455 1.130 2.869 ;
        RECT 1.130 2.465 1.140 2.869 ;
        RECT 1.140 2.475 1.150 2.869 ;
        RECT 1.150 2.485 1.160 2.869 ;
        RECT 1.160 2.495 1.170 2.869 ;
        RECT 1.170 2.505 1.180 2.869 ;
        RECT 1.180 2.515 1.190 2.869 ;
        RECT 1.190 2.525 1.200 2.869 ;
        RECT 1.200 2.535 1.210 2.869 ;
        RECT 1.210 2.545 1.220 2.869 ;
        RECT 1.220 2.555 1.230 2.869 ;
        RECT 1.230 2.565 1.240 2.869 ;
        RECT 1.240 2.575 1.250 2.869 ;
        RECT 1.030 2.365 1.040 2.605 ;
        RECT 1.040 2.375 1.050 2.615 ;
        RECT 1.050 2.385 1.060 2.625 ;
        RECT 1.060 2.395 1.070 2.635 ;
        RECT 1.070 2.405 1.080 2.645 ;
        RECT 0.860 1.520 0.870 2.434 ;
        RECT 0.870 1.520 0.880 2.444 ;
        RECT 0.880 1.520 0.890 2.454 ;
        RECT 0.890 1.520 0.900 2.464 ;
        RECT 0.900 1.520 0.910 2.474 ;
        RECT 0.910 1.520 0.920 2.484 ;
        RECT 0.920 1.520 0.930 2.494 ;
        RECT 0.930 1.520 0.940 2.504 ;
        RECT 0.940 1.520 0.950 2.514 ;
        RECT 0.950 1.520 0.960 2.524 ;
        RECT 0.960 1.520 0.970 2.534 ;
        RECT 0.970 1.520 0.980 2.544 ;
        RECT 0.980 1.520 0.990 2.554 ;
        RECT 0.990 1.520 1.000 2.564 ;
        RECT 1.000 1.520 1.010 2.574 ;
        RECT 1.010 1.520 1.020 2.584 ;
        RECT 1.020 1.520 1.030 2.594 ;
        RECT 2.450 0.925 2.620 2.410 ;
        RECT 2.445 2.110 2.620 2.410 ;
        RECT 2.450 0.925 2.965 1.095 ;
        RECT 1.085 1.125 1.210 1.295 ;
        RECT 1.540 2.350 2.050 2.520 ;
        RECT 2.365 2.590 3.135 2.760 ;
        RECT 2.800 1.345 2.970 2.760 ;
        RECT 2.965 2.570 3.135 3.150 ;
        RECT 2.800 1.345 3.875 1.515 ;
        RECT 2.290 2.525 2.300 2.759 ;
        RECT 2.300 2.535 2.310 2.759 ;
        RECT 2.310 2.545 2.320 2.759 ;
        RECT 2.320 2.555 2.330 2.759 ;
        RECT 2.330 2.565 2.340 2.759 ;
        RECT 2.340 2.575 2.350 2.759 ;
        RECT 2.350 2.585 2.360 2.759 ;
        RECT 2.360 2.590 2.366 2.760 ;
        RECT 2.125 2.360 2.135 2.594 ;
        RECT 2.135 2.370 2.145 2.604 ;
        RECT 2.145 2.380 2.155 2.614 ;
        RECT 2.155 2.390 2.165 2.624 ;
        RECT 2.165 2.400 2.175 2.634 ;
        RECT 2.175 2.410 2.185 2.644 ;
        RECT 2.185 2.420 2.195 2.654 ;
        RECT 2.195 2.430 2.205 2.664 ;
        RECT 2.205 2.440 2.215 2.674 ;
        RECT 2.215 2.450 2.225 2.684 ;
        RECT 2.225 2.460 2.235 2.694 ;
        RECT 2.235 2.470 2.245 2.704 ;
        RECT 2.245 2.480 2.255 2.714 ;
        RECT 2.255 2.490 2.265 2.724 ;
        RECT 2.265 2.500 2.275 2.734 ;
        RECT 2.275 2.510 2.285 2.744 ;
        RECT 2.285 2.515 2.291 2.755 ;
        RECT 2.050 2.350 2.060 2.520 ;
        RECT 2.060 2.350 2.070 2.530 ;
        RECT 2.070 2.350 2.080 2.540 ;
        RECT 2.080 2.350 2.090 2.550 ;
        RECT 2.090 2.350 2.100 2.560 ;
        RECT 2.100 2.350 2.110 2.570 ;
        RECT 2.110 2.350 2.120 2.580 ;
        RECT 2.120 2.350 2.126 2.590 ;
        RECT 1.450 2.270 1.460 2.520 ;
        RECT 1.460 2.280 1.470 2.520 ;
        RECT 1.470 2.290 1.480 2.520 ;
        RECT 1.480 2.300 1.490 2.520 ;
        RECT 1.490 2.310 1.500 2.520 ;
        RECT 1.500 2.320 1.510 2.520 ;
        RECT 1.510 2.330 1.520 2.520 ;
        RECT 1.520 2.340 1.530 2.520 ;
        RECT 1.530 2.350 1.540 2.520 ;
        RECT 1.385 2.205 1.395 2.455 ;
        RECT 1.395 2.215 1.405 2.465 ;
        RECT 1.405 2.225 1.415 2.475 ;
        RECT 1.415 2.235 1.425 2.485 ;
        RECT 1.425 2.245 1.435 2.495 ;
        RECT 1.435 2.255 1.445 2.505 ;
        RECT 1.445 2.260 1.451 2.514 ;
        RECT 1.210 1.125 1.220 2.279 ;
        RECT 1.220 1.125 1.230 2.289 ;
        RECT 1.230 1.125 1.240 2.299 ;
        RECT 1.240 1.125 1.250 2.309 ;
        RECT 1.250 1.125 1.260 2.319 ;
        RECT 1.260 1.125 1.270 2.329 ;
        RECT 1.270 1.125 1.280 2.339 ;
        RECT 1.280 1.125 1.290 2.349 ;
        RECT 1.290 1.125 1.300 2.359 ;
        RECT 1.300 1.125 1.310 2.369 ;
        RECT 1.310 1.125 1.320 2.379 ;
        RECT 1.320 1.125 1.330 2.389 ;
        RECT 1.330 1.125 1.340 2.399 ;
        RECT 1.340 1.125 1.350 2.409 ;
        RECT 1.350 1.125 1.360 2.419 ;
        RECT 1.360 1.125 1.370 2.429 ;
        RECT 1.370 1.125 1.380 2.439 ;
        RECT 1.380 1.125 1.386 2.449 ;
        RECT 3.150 2.035 3.325 2.345 ;
        RECT 3.180 0.925 4.230 1.095 ;
        RECT 4.060 0.925 4.230 2.215 ;
        RECT 5.330 1.670 5.500 2.215 ;
        RECT 3.150 2.035 5.500 2.215 ;
        RECT 4.205 2.395 4.375 2.735 ;
        RECT 3.745 2.565 4.375 2.735 ;
        RECT 5.355 1.125 5.850 1.295 ;
        RECT 4.205 2.395 5.850 2.565 ;
        RECT 5.680 1.125 5.850 2.795 ;
        RECT 7.375 1.540 7.545 2.630 ;
        RECT 5.680 2.460 7.545 2.630 ;
  END 
END LATNRHD2XHT

MACRO LATNRHD1XHT
  CLASS  CORE ;
  FOREIGN LATNRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.380 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.840 0.720 6.170 1.200 ;
        RECT 6.000 0.720 6.170 2.280 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.465 0.380 2.840 ;
        RECT 0.100 2.465 0.585 2.635 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.040 0.720 7.210 2.960 ;
        RECT 7.040 2.080 7.280 2.425 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.595 2.090 2.135 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.355 0.645 1.525 0.945 ;
        RECT 2.080 0.575 2.250 0.945 ;
        RECT 1.355 0.775 2.250 0.945 ;
        RECT 2.080 0.575 4.570 0.745 ;
        RECT 4.400 0.575 4.570 1.800 ;
        RECT 4.400 1.330 4.615 1.800 ;
        RECT 4.400 1.330 4.900 1.540 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.715 ;
        RECT 1.725 -0.300 1.895 0.575 ;
        RECT 4.750 -0.300 5.050 1.095 ;
        RECT 6.455 -0.300 6.755 1.055 ;
        RECT 0.000 -0.300 7.380 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.665 2.835 0.965 3.990 ;
        RECT 1.625 3.095 1.925 3.990 ;
        RECT 4.010 2.505 4.310 3.990 ;
        RECT 4.980 2.650 5.280 3.990 ;
        RECT 6.455 2.975 6.755 3.990 ;
        RECT 0.000 3.390 7.380 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.445 0.925 2.615 2.215 ;
        RECT 2.315 2.045 2.615 2.215 ;
        RECT 2.445 0.925 2.945 1.095 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.520 1.030 1.690 ;
        RECT 0.860 1.520 1.030 2.655 ;
        RECT 0.860 2.485 1.080 2.655 ;
        RECT 1.145 2.485 1.155 2.915 ;
        RECT 1.315 2.745 2.290 2.915 ;
        RECT 2.120 2.745 2.290 3.135 ;
        RECT 3.335 2.470 3.505 3.135 ;
        RECT 2.120 2.965 3.505 3.135 ;
        RECT 1.155 2.495 1.165 2.915 ;
        RECT 1.165 2.505 1.175 2.915 ;
        RECT 1.175 2.515 1.185 2.915 ;
        RECT 1.185 2.525 1.195 2.915 ;
        RECT 1.195 2.535 1.205 2.915 ;
        RECT 1.205 2.545 1.215 2.915 ;
        RECT 1.215 2.555 1.225 2.915 ;
        RECT 1.225 2.565 1.235 2.915 ;
        RECT 1.235 2.575 1.245 2.915 ;
        RECT 1.245 2.585 1.255 2.915 ;
        RECT 1.255 2.595 1.265 2.915 ;
        RECT 1.265 2.605 1.275 2.915 ;
        RECT 1.275 2.615 1.285 2.915 ;
        RECT 1.285 2.625 1.295 2.915 ;
        RECT 1.295 2.635 1.305 2.915 ;
        RECT 1.305 2.645 1.315 2.915 ;
        RECT 1.080 2.485 1.090 2.655 ;
        RECT 1.090 2.485 1.100 2.665 ;
        RECT 1.100 2.485 1.110 2.675 ;
        RECT 1.110 2.485 1.120 2.685 ;
        RECT 1.120 2.485 1.130 2.695 ;
        RECT 1.130 2.485 1.140 2.705 ;
        RECT 1.140 2.485 1.146 2.715 ;
        RECT 1.085 1.125 1.210 1.295 ;
        RECT 1.570 2.395 2.975 2.565 ;
        RECT 2.805 1.345 2.975 2.785 ;
        RECT 2.630 2.395 2.975 2.785 ;
        RECT 2.805 1.345 3.830 1.515 ;
        RECT 1.495 2.330 1.505 2.564 ;
        RECT 1.505 2.340 1.515 2.564 ;
        RECT 1.515 2.350 1.525 2.564 ;
        RECT 1.525 2.360 1.535 2.564 ;
        RECT 1.535 2.370 1.545 2.564 ;
        RECT 1.545 2.380 1.555 2.564 ;
        RECT 1.555 2.390 1.565 2.564 ;
        RECT 1.565 2.395 1.571 2.565 ;
        RECT 1.405 2.240 1.415 2.474 ;
        RECT 1.415 2.250 1.425 2.484 ;
        RECT 1.425 2.260 1.435 2.494 ;
        RECT 1.435 2.270 1.445 2.504 ;
        RECT 1.445 2.280 1.455 2.514 ;
        RECT 1.455 2.290 1.465 2.524 ;
        RECT 1.465 2.300 1.475 2.534 ;
        RECT 1.475 2.310 1.485 2.544 ;
        RECT 1.485 2.320 1.495 2.554 ;
        RECT 1.210 1.125 1.220 2.279 ;
        RECT 1.220 1.125 1.230 2.289 ;
        RECT 1.230 1.125 1.240 2.299 ;
        RECT 1.240 1.125 1.250 2.309 ;
        RECT 1.250 1.125 1.260 2.319 ;
        RECT 1.260 1.125 1.270 2.329 ;
        RECT 1.270 1.125 1.280 2.339 ;
        RECT 1.280 1.125 1.290 2.349 ;
        RECT 1.290 1.125 1.300 2.359 ;
        RECT 1.300 1.125 1.310 2.369 ;
        RECT 1.310 1.125 1.320 2.379 ;
        RECT 1.320 1.125 1.330 2.389 ;
        RECT 1.330 1.125 1.340 2.399 ;
        RECT 1.340 1.125 1.350 2.409 ;
        RECT 1.350 1.125 1.360 2.419 ;
        RECT 1.360 1.125 1.370 2.429 ;
        RECT 1.370 1.125 1.380 2.439 ;
        RECT 1.380 1.125 1.390 2.449 ;
        RECT 1.390 1.125 1.400 2.459 ;
        RECT 1.400 1.125 1.406 2.469 ;
        RECT 3.155 1.980 3.325 2.280 ;
        RECT 3.155 2.045 3.330 2.280 ;
        RECT 3.165 0.925 4.220 1.095 ;
        RECT 4.050 0.925 4.220 2.215 ;
        RECT 5.175 1.770 5.345 2.215 ;
        RECT 3.155 2.045 5.345 2.215 ;
        RECT 5.345 0.860 5.515 1.550 ;
        RECT 5.345 1.380 5.735 1.550 ;
        RECT 5.565 1.380 5.735 3.205 ;
        RECT 6.025 2.460 6.195 3.205 ;
        RECT 5.565 3.035 6.195 3.205 ;
        RECT 6.660 1.540 6.830 2.630 ;
        RECT 6.025 2.460 6.830 2.630 ;
  END 
END LATNRHD1XHT

MACRO LATNHDMXHT
  CLASS  CORE ;
  FOREIGN LATNHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.150 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.770 1.060 5.940 2.425 ;
        RECT 5.770 2.080 6.050 2.425 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.495 0.510 2.950 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.610 0.850 4.900 1.210 ;
        RECT 4.730 0.850 4.900 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.670 1.585 2.165 1.950 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 1.655 -0.300 1.955 0.900 ;
        RECT 3.465 -0.300 3.765 1.190 ;
        RECT 5.185 -0.300 5.485 1.145 ;
        RECT 0.000 -0.300 6.150 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.280 0.860 3.990 ;
        RECT 1.655 2.485 1.955 3.990 ;
        RECT 3.495 2.860 3.795 3.990 ;
        RECT 5.155 2.925 5.455 3.990 ;
        RECT 0.000 3.390 6.150 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.520 1.030 1.820 ;
        RECT 1.210 1.060 1.380 2.305 ;
        RECT 1.210 2.135 2.405 2.305 ;
        RECT 2.235 2.135 2.405 3.030 ;
        RECT 2.290 0.605 2.460 1.250 ;
        RECT 1.210 1.080 2.460 1.250 ;
        RECT 2.235 2.860 2.695 3.030 ;
        RECT 2.290 0.605 3.055 0.775 ;
        RECT 3.285 1.790 3.585 1.960 ;
        RECT 3.415 1.790 3.585 2.330 ;
        RECT 3.985 1.020 4.415 1.190 ;
        RECT 4.245 1.020 4.415 2.330 ;
        RECT 3.415 2.160 4.415 2.330 ;
        RECT 4.245 1.520 4.550 1.820 ;
        RECT 2.640 0.955 2.810 2.680 ;
        RECT 2.640 1.440 4.065 1.610 ;
        RECT 5.420 1.520 5.590 2.680 ;
        RECT 2.640 2.510 5.590 2.680 ;
  END 
END LATNHDMXHT

MACRO LATNHDLXHT
  CLASS  CORE ;
  FOREIGN LATNHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.150 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.770 1.060 5.940 2.425 ;
        RECT 5.770 2.085 6.050 2.425 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.475 0.510 2.910 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.610 0.850 4.900 1.200 ;
        RECT 4.730 0.850 4.900 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.655 1.585 2.125 1.950 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.785 ;
        RECT 1.565 -0.300 1.865 0.820 ;
        RECT 3.405 -0.300 3.705 0.745 ;
        RECT 5.185 -0.300 5.485 1.295 ;
        RECT 0.000 -0.300 6.150 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.120 0.860 3.990 ;
        RECT 1.625 2.685 1.925 3.990 ;
        RECT 3.405 2.925 3.705 3.990 ;
        RECT 5.155 2.925 5.455 3.990 ;
        RECT 0.000 3.390 6.150 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.520 1.030 1.820 ;
        RECT 1.210 1.060 1.380 2.305 ;
        RECT 1.210 2.135 2.375 2.305 ;
        RECT 2.175 0.705 2.345 1.230 ;
        RECT 1.210 1.060 2.345 1.230 ;
        RECT 2.205 2.135 2.375 2.810 ;
        RECT 2.205 2.640 2.665 2.810 ;
        RECT 2.175 0.705 3.025 0.875 ;
        RECT 3.255 1.850 3.555 2.020 ;
        RECT 3.385 1.850 3.555 2.395 ;
        RECT 3.955 1.125 4.425 1.295 ;
        RECT 4.255 1.125 4.425 2.395 ;
        RECT 3.385 2.225 4.425 2.395 ;
        RECT 4.255 1.520 4.550 1.820 ;
        RECT 2.580 1.060 2.780 2.460 ;
        RECT 2.580 2.290 3.055 2.460 ;
        RECT 2.885 2.290 3.055 2.745 ;
        RECT 2.580 1.500 4.075 1.670 ;
        RECT 5.420 1.540 5.590 2.745 ;
        RECT 2.885 2.575 5.590 2.745 ;
  END 
END LATNHDLXHT

MACRO LATNHD2XHT
  CLASS  CORE ;
  FOREIGN LATNHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.970 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 6.110 0.715 6.280 2.960 ;
        RECT 6.110 0.715 6.320 1.610 ;
        RECT 6.110 1.260 6.460 1.610 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.490 0.510 2.950 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.020 0.720 5.240 1.195 ;
        RECT 5.050 0.720 5.240 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.945 1.585 2.445 1.950 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.540 -0.300 0.840 0.745 ;
        RECT 1.780 -0.300 1.950 1.040 ;
        RECT 3.515 -0.300 3.815 0.635 ;
        RECT 4.485 -0.300 4.785 0.715 ;
        RECT 5.525 -0.300 5.825 1.055 ;
        RECT 6.565 -0.300 6.865 1.055 ;
        RECT 0.000 -0.300 6.970 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.280 0.860 3.990 ;
        RECT 1.715 2.635 2.015 3.990 ;
        RECT 3.465 2.895 3.765 3.990 ;
        RECT 4.485 2.975 4.785 3.990 ;
        RECT 5.525 2.975 5.825 3.990 ;
        RECT 6.565 2.295 6.865 3.990 ;
        RECT 0.000 3.390 6.970 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.520 1.000 1.820 ;
        RECT 1.180 1.060 1.350 2.310 ;
        RECT 1.180 1.980 1.380 2.310 ;
        RECT 1.180 2.140 2.440 2.310 ;
        RECT 2.265 0.515 2.435 1.400 ;
        RECT 1.180 1.230 2.435 1.400 ;
        RECT 2.270 2.140 2.440 3.145 ;
        RECT 2.265 0.515 3.185 0.685 ;
        RECT 2.270 2.975 3.185 3.145 ;
        RECT 3.315 1.825 3.615 1.995 ;
        RECT 3.445 1.825 3.615 2.365 ;
        RECT 4.065 1.125 4.830 1.295 ;
        RECT 4.660 1.125 4.830 2.365 ;
        RECT 3.445 2.195 4.830 2.365 ;
        RECT 2.670 0.960 2.840 2.715 ;
        RECT 2.670 1.475 4.135 1.645 ;
        RECT 3.835 1.475 4.135 1.665 ;
        RECT 5.760 1.520 5.930 2.715 ;
        RECT 2.670 2.545 5.930 2.715 ;
  END 
END LATNHD2XHT

MACRO LATNHD1XHT
  CLASS  CORE ;
  FOREIGN LATNHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.150 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.770 0.720 5.940 2.960 ;
        RECT 5.770 2.085 6.050 2.430 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.495 0.510 2.950 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.610 0.835 4.900 1.225 ;
        RECT 4.730 0.720 4.900 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.655 1.585 2.145 1.950 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 1.655 -0.300 1.955 0.920 ;
        RECT 3.500 -0.300 3.800 1.195 ;
        RECT 5.185 -0.300 5.485 1.055 ;
        RECT 0.000 -0.300 6.150 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.280 0.860 3.990 ;
        RECT 1.655 2.545 1.955 3.990 ;
        RECT 3.465 2.925 3.765 3.990 ;
        RECT 5.185 2.975 5.485 3.990 ;
        RECT 0.000 3.390 6.150 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.520 1.030 1.820 ;
        RECT 1.210 1.125 1.380 2.300 ;
        RECT 1.210 2.130 2.375 2.300 ;
        RECT 2.205 2.130 2.375 3.095 ;
        RECT 2.240 0.605 2.410 1.295 ;
        RECT 1.145 1.125 2.410 1.295 ;
        RECT 2.205 2.925 2.665 3.095 ;
        RECT 2.240 0.605 3.060 0.775 ;
        RECT 3.255 1.850 3.555 2.020 ;
        RECT 3.385 1.850 3.555 2.395 ;
        RECT 4.045 1.025 4.385 1.195 ;
        RECT 4.215 1.025 4.385 2.395 ;
        RECT 3.385 2.225 4.385 2.395 ;
        RECT 4.215 1.520 4.550 1.820 ;
        RECT 2.610 0.960 2.780 2.745 ;
        RECT 2.610 0.960 2.810 1.260 ;
        RECT 2.610 1.500 4.035 1.670 ;
        RECT 5.420 1.520 5.590 2.745 ;
        RECT 2.610 2.575 5.590 2.745 ;
  END 
END LATNHD1XHT

MACRO LATHDMXHT
  CLASS  CORE ;
  FOREIGN LATHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.150 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.770 1.060 5.940 2.430 ;
        RECT 5.770 2.085 6.050 2.430 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.610 0.835 4.905 1.360 ;
        RECT 4.735 0.835 4.905 2.280 ;
        RECT 4.650 1.980 4.905 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.645 1.585 2.165 1.950 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.490 0.510 2.930 ;
    END
  END G
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 1.655 -0.300 1.955 0.930 ;
        RECT 3.465 -0.300 3.765 1.295 ;
        RECT 5.150 -0.300 5.450 1.145 ;
        RECT 0.000 -0.300 6.150 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.130 0.860 3.990 ;
        RECT 1.655 2.500 1.955 3.990 ;
        RECT 3.495 2.925 3.795 3.990 ;
        RECT 5.135 2.925 5.435 3.990 ;
        RECT 0.000 3.390 6.150 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.520 1.030 1.820 ;
        RECT 1.210 1.125 1.380 2.315 ;
        RECT 1.210 2.145 2.405 2.315 ;
        RECT 2.235 2.145 2.405 3.095 ;
        RECT 2.290 0.705 2.460 1.295 ;
        RECT 1.145 1.125 2.460 1.295 ;
        RECT 2.290 0.705 2.695 0.875 ;
        RECT 2.235 2.925 3.055 3.095 ;
        RECT 3.285 1.850 3.585 2.020 ;
        RECT 3.415 1.850 3.585 2.395 ;
        RECT 4.050 1.125 4.415 1.295 ;
        RECT 4.245 1.125 4.415 2.395 ;
        RECT 3.415 2.225 4.415 2.395 ;
        RECT 4.245 1.585 4.555 1.755 ;
        RECT 2.640 1.060 2.810 2.745 ;
        RECT 2.640 1.500 4.065 1.670 ;
        RECT 5.420 1.520 5.590 2.745 ;
        RECT 2.640 2.575 5.590 2.745 ;
  END 
END LATHDMXHT

MACRO LATHD1XHT
  CLASS  CORE ;
  FOREIGN LATHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.150 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.770 0.720 5.940 2.960 ;
        RECT 5.770 2.090 6.050 2.425 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.610 0.850 4.900 1.205 ;
        RECT 4.730 0.720 4.900 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.680 1.585 2.135 1.950 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.495 0.510 2.955 ;
    END
  END G
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 1.625 -0.300 1.925 0.780 ;
        RECT 3.435 -0.300 3.735 1.295 ;
        RECT 5.185 -0.300 5.485 1.055 ;
        RECT 0.000 -0.300 6.150 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.280 0.860 3.990 ;
        RECT 1.655 2.545 1.955 3.990 ;
        RECT 3.405 2.995 3.705 3.990 ;
        RECT 5.185 2.975 5.485 3.990 ;
        RECT 0.000 3.390 6.150 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.520 1.030 1.820 ;
        RECT 1.210 1.060 1.380 2.300 ;
        RECT 1.210 2.130 2.375 2.300 ;
        RECT 2.205 2.130 2.375 3.095 ;
        RECT 2.260 0.605 2.430 1.230 ;
        RECT 1.210 1.060 2.430 1.230 ;
        RECT 2.260 0.605 2.665 0.775 ;
        RECT 2.205 2.925 3.025 3.095 ;
        RECT 3.255 1.850 3.555 2.020 ;
        RECT 3.385 1.850 3.555 2.395 ;
        RECT 3.955 1.125 4.430 1.295 ;
        RECT 4.260 1.125 4.430 2.395 ;
        RECT 3.385 2.225 4.430 2.395 ;
        RECT 4.260 1.520 4.550 1.820 ;
        RECT 2.610 1.060 2.780 2.745 ;
        RECT 2.610 1.500 4.075 1.670 ;
        RECT 5.420 1.520 5.590 2.745 ;
        RECT 2.610 2.575 5.590 2.745 ;
  END 
END LATHD1XHT

MACRO INVTSHDUXHT
  CLASS  CORE ;
  FOREIGN INVTSHDUXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.240 1.585 0.810 1.950 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.895 1.495 2.360 2.015 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 0.785 ;
        RECT 2.025 -0.300 2.325 0.845 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 1.040 1.060 1.230 2.770 ;
        RECT 0.855 2.560 1.230 2.770 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.265 0.405 3.990 ;
        RECT 2.025 2.750 2.325 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.425 1.120 1.605 2.380 ;
        RECT 1.425 1.120 1.805 1.300 ;
        RECT 1.425 2.200 1.805 2.380 ;
  END 
END INVTSHDUXHT

MACRO INVTSHDMXHT
  CLASS  CORE ;
  FOREIGN INVTSHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.330 1.500 0.860 1.950 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.910 1.520 2.360 2.015 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.005 ;
        RECT 2.025 -0.300 2.325 1.295 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 0.855 2.560 1.230 2.770 ;
        RECT 1.060 1.060 1.230 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.235 0.405 3.990 ;
        RECT 2.025 2.325 2.325 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.425 1.120 1.605 2.380 ;
        RECT 1.425 1.120 1.805 1.300 ;
        RECT 1.425 2.200 1.805 2.380 ;
  END 
END INVTSHDMXHT

MACRO INVTSHD2XHT
  CLASS  CORE ;
  FOREIGN INVTSHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.740 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.585 0.850 1.950 ;
        RECT 0.440 1.585 2.130 1.755 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.200 1.250 4.435 1.860 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.875 ;
        RECT 1.665 -0.300 1.965 0.875 ;
        RECT 5.295 -0.300 5.595 1.235 ;
        RECT 0.000 -0.300 5.740 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 2.705 0.975 3.005 2.555 ;
        RECT 2.705 1.540 4.000 1.840 ;
        RECT 3.790 0.910 4.000 2.620 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.545 0.925 3.990 ;
        RECT 1.665 2.545 1.965 3.990 ;
        RECT 5.295 2.545 5.595 3.990 ;
        RECT 0.000 3.390 5.740 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 2.140 0.340 3.120 ;
        RECT 1.210 2.140 1.380 3.120 ;
        RECT 0.170 2.140 2.420 2.310 ;
        RECT 2.250 2.140 2.420 3.120 ;
        RECT 3.290 2.135 3.460 3.120 ;
        RECT 4.330 2.140 4.500 3.120 ;
        RECT 2.250 2.950 4.500 3.120 ;
        RECT 0.170 0.920 0.340 1.300 ;
        RECT 1.210 0.910 1.380 1.300 ;
        RECT 2.250 0.560 2.420 1.300 ;
        RECT 0.170 1.130 2.420 1.300 ;
        RECT 3.290 0.560 3.460 0.940 ;
        RECT 2.250 0.560 4.500 0.730 ;
        RECT 4.330 0.560 4.500 0.940 ;
        RECT 4.700 0.720 5.025 2.780 ;
  END 
END INVTSHD2XHT

MACRO INVTSHD1XHT
  CLASS  CORE ;
  FOREIGN INVTSHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.435 1.585 1.100 1.950 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.145 1.265 2.375 1.860 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.875 ;
        RECT 3.215 -0.300 3.515 1.245 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 1.665 0.975 1.965 2.555 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.545 0.925 3.990 ;
        RECT 3.215 2.395 3.515 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 2.140 0.340 3.120 ;
        RECT 0.170 2.140 1.380 2.310 ;
        RECT 1.210 2.140 1.380 3.120 ;
        RECT 2.250 2.140 2.420 3.120 ;
        RECT 1.210 2.950 2.420 3.120 ;
        RECT 0.170 0.920 0.340 1.300 ;
        RECT 1.210 0.580 1.380 1.300 ;
        RECT 0.170 1.130 1.380 1.300 ;
        RECT 1.210 0.580 2.420 0.750 ;
        RECT 2.250 0.580 2.420 0.940 ;
        RECT 2.620 1.060 2.945 2.440 ;
  END 
END INVTSHD1XHT

MACRO INVTSHDLXHT
  CLASS  CORE ;
  FOREIGN INVTSHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.240 1.585 0.810 1.950 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.895 1.495 2.360 2.015 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.195 ;
        RECT 2.025 -0.300 2.325 1.295 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 1.040 1.060 1.230 2.770 ;
        RECT 0.855 2.560 1.230 2.770 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.185 0.405 3.990 ;
        RECT 2.025 2.325 2.325 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.425 1.120 1.605 2.380 ;
        RECT 1.425 1.120 1.805 1.300 ;
        RECT 1.425 2.200 1.805 2.380 ;
  END 
END INVTSHDLXHT

MACRO INVTSHD8XHT
  CLASS  CORE ;
  FOREIGN INVTSHD8XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 9.890 1.575 10.195 2.020 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.610 0.685 2.020 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.745 -0.300 1.045 0.715 ;
        RECT 3.695 -0.300 3.995 1.055 ;
        RECT 4.735 -0.300 5.035 1.055 ;
        RECT 5.775 -0.300 6.075 1.055 ;
        RECT 6.815 -0.300 7.115 1.055 ;
        RECT 8.595 -0.300 8.895 0.715 ;
        RECT 9.635 -0.300 9.935 0.715 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 3.240 0.720 3.410 2.965 ;
        RECT 4.280 0.720 4.450 2.965 ;
        RECT 5.320 0.720 5.490 2.960 ;
        RECT 6.360 0.720 6.530 2.960 ;
        RECT 3.240 1.360 7.570 2.090 ;
        RECT 7.400 0.720 7.570 2.960 ;
        RECT 7.390 1.360 7.570 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.745 2.975 1.045 3.990 ;
        RECT 3.695 2.290 3.995 3.990 ;
        RECT 4.735 2.290 5.035 3.990 ;
        RECT 5.775 2.290 6.075 3.990 ;
        RECT 6.815 2.290 7.115 3.990 ;
        RECT 8.595 2.295 8.895 3.990 ;
        RECT 9.635 2.635 9.935 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.140 0.480 0.460 0.650 ;
        RECT 0.290 0.480 0.460 1.365 ;
        RECT 0.290 1.175 1.110 1.365 ;
        RECT 0.940 1.175 1.110 2.380 ;
        RECT 0.225 2.205 1.110 2.380 ;
        RECT 0.940 2.105 1.845 2.275 ;
        RECT 1.330 1.020 1.500 1.520 ;
        RECT 2.025 1.320 2.195 2.645 ;
        RECT 1.785 2.475 2.195 2.645 ;
        RECT 2.305 1.085 2.605 1.690 ;
        RECT 1.330 1.320 2.605 1.520 ;
        RECT 2.025 1.390 2.680 1.690 ;
        RECT 1.330 2.710 1.500 3.075 ;
        RECT 1.850 0.720 2.020 1.020 ;
        RECT 2.375 2.010 2.545 3.075 ;
        RECT 1.330 2.875 2.545 3.075 ;
        RECT 1.850 0.720 3.040 0.890 ;
        RECT 2.870 0.720 3.040 2.210 ;
        RECT 2.375 2.010 3.040 2.210 ;
        RECT 7.765 1.770 7.945 2.105 ;
        RECT 8.140 1.925 8.310 2.965 ;
        RECT 7.765 1.925 9.355 2.105 ;
        RECT 9.175 1.925 9.355 2.960 ;
        RECT 7.765 1.215 7.945 1.570 ;
        RECT 8.140 0.720 8.310 1.395 ;
        RECT 9.175 0.720 9.355 1.395 ;
        RECT 7.765 1.215 9.355 1.395 ;
        RECT 8.480 1.575 9.710 1.745 ;
        RECT 9.540 1.035 9.710 2.455 ;
        RECT 9.540 2.285 10.390 2.455 ;
        RECT 10.220 0.565 10.390 1.205 ;
        RECT 9.540 1.035 10.390 1.205 ;
        RECT 10.220 2.285 10.390 2.925 ;
  END 
END INVTSHD8XHT

MACRO INVTSHD7XHT
  CLASS  CORE ;
  FOREIGN INVTSHD7XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 9.940 1.540 10.265 2.160 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.890 1.540 1.465 2.020 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.130 -0.300 1.430 0.715 ;
        RECT 3.275 -0.300 3.575 1.120 ;
        RECT 4.315 -0.300 4.615 1.120 ;
        RECT 5.355 -0.300 5.655 1.120 ;
        RECT 6.395 -0.300 6.695 0.780 ;
        RECT 7.435 -0.300 7.735 1.120 ;
        RECT 8.475 -0.300 8.775 1.055 ;
        RECT 10.025 -0.300 10.325 1.200 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 3.795 0.610 4.095 1.470 ;
        RECT 3.795 2.220 4.095 3.210 ;
        RECT 3.795 1.300 6.095 1.470 ;
        RECT 4.835 0.610 5.135 3.110 ;
        RECT 5.875 0.610 6.095 3.110 ;
        RECT 4.335 1.300 6.095 2.455 ;
        RECT 5.875 0.610 6.175 1.215 ;
        RECT 5.875 2.130 6.175 3.110 ;
        RECT 4.335 2.130 6.555 2.455 ;
        RECT 4.335 2.200 7.215 2.455 ;
        RECT 3.795 2.220 7.215 2.455 ;
        RECT 6.915 0.575 7.215 1.215 ;
        RECT 5.875 0.980 7.215 1.215 ;
        RECT 6.915 2.200 7.215 3.180 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.085 2.975 1.385 3.990 ;
        RECT 3.275 2.230 3.575 3.990 ;
        RECT 4.315 2.635 4.615 3.990 ;
        RECT 5.355 2.635 5.655 3.990 ;
        RECT 6.395 2.635 6.695 3.990 ;
        RECT 7.435 2.460 7.735 3.990 ;
        RECT 8.475 2.460 8.775 3.990 ;
        RECT 10.025 2.460 10.325 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.140 1.495 0.640 1.665 ;
        RECT 0.470 1.125 0.640 2.400 ;
        RECT 0.470 2.165 0.780 2.400 ;
        RECT 0.470 1.125 0.785 1.295 ;
        RECT 1.720 2.105 1.890 2.400 ;
        RECT 0.470 2.230 1.890 2.400 ;
        RECT 1.720 2.105 2.245 2.275 ;
        RECT 0.350 0.565 0.770 0.735 ;
        RECT 1.105 0.945 1.885 1.115 ;
        RECT 1.715 0.535 1.885 1.585 ;
        RECT 1.715 1.405 2.595 1.585 ;
        RECT 2.425 1.405 2.595 2.645 ;
        RECT 2.215 2.475 2.595 2.645 ;
        RECT 1.715 0.535 3.050 0.705 ;
        RECT 2.750 0.535 3.050 0.805 ;
        RECT 1.035 0.885 1.045 1.115 ;
        RECT 1.045 0.895 1.055 1.115 ;
        RECT 1.055 0.905 1.065 1.115 ;
        RECT 1.065 0.915 1.075 1.115 ;
        RECT 1.075 0.925 1.085 1.115 ;
        RECT 1.085 0.935 1.095 1.115 ;
        RECT 1.095 0.945 1.105 1.115 ;
        RECT 0.950 0.800 0.960 1.030 ;
        RECT 0.960 0.810 0.970 1.040 ;
        RECT 0.970 0.820 0.980 1.050 ;
        RECT 0.980 0.830 0.990 1.060 ;
        RECT 0.990 0.840 1.000 1.070 ;
        RECT 1.000 0.850 1.010 1.080 ;
        RECT 1.010 0.860 1.020 1.090 ;
        RECT 1.020 0.870 1.030 1.100 ;
        RECT 1.030 0.875 1.036 1.109 ;
        RECT 0.770 0.565 0.780 0.849 ;
        RECT 0.780 0.565 0.790 0.859 ;
        RECT 0.790 0.565 0.800 0.869 ;
        RECT 0.800 0.565 0.810 0.879 ;
        RECT 0.810 0.565 0.820 0.889 ;
        RECT 0.820 0.565 0.830 0.899 ;
        RECT 0.830 0.565 0.840 0.909 ;
        RECT 0.840 0.565 0.850 0.919 ;
        RECT 0.850 0.565 0.860 0.929 ;
        RECT 0.860 0.565 0.870 0.939 ;
        RECT 0.870 0.565 0.880 0.949 ;
        RECT 0.880 0.565 0.890 0.959 ;
        RECT 0.890 0.565 0.900 0.969 ;
        RECT 0.900 0.565 0.910 0.979 ;
        RECT 0.910 0.565 0.920 0.989 ;
        RECT 0.920 0.565 0.930 0.999 ;
        RECT 0.930 0.565 0.940 1.009 ;
        RECT 0.940 0.565 0.950 1.019 ;
        RECT 0.550 2.625 0.720 3.060 ;
        RECT 0.550 2.625 1.965 2.795 ;
        RECT 1.665 2.625 1.965 3.145 ;
        RECT 2.200 0.885 2.500 1.155 ;
        RECT 2.200 0.985 3.000 1.155 ;
        RECT 2.830 0.985 3.000 3.145 ;
        RECT 1.665 2.975 3.000 3.145 ;
        RECT 2.830 1.825 4.135 1.995 ;
        RECT 6.755 1.825 8.125 1.995 ;
        RECT 7.955 1.825 8.125 3.005 ;
        RECT 7.955 2.090 8.255 3.005 ;
        RECT 7.955 2.090 9.295 2.260 ;
        RECT 8.995 2.090 9.295 3.005 ;
        RECT 7.955 0.640 8.125 1.565 ;
        RECT 6.275 1.395 8.125 1.565 ;
        RECT 7.955 0.640 8.255 1.405 ;
        RECT 7.955 1.235 9.295 1.405 ;
        RECT 8.995 0.640 9.295 1.405 ;
        RECT 8.315 1.675 9.685 1.845 ;
        RECT 9.505 0.720 9.685 2.930 ;
        RECT 9.505 0.720 9.805 1.360 ;
        RECT 9.505 2.290 9.805 2.930 ;
  END 
END INVTSHD7XHT

MACRO INVTSHD6XHT
  CLASS  CORE ;
  FOREIGN INVTSHD6XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.610 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.760 1.310 8.100 2.020 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.540 0.870 2.020 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 -0.300 0.990 1.120 ;
        RECT 3.355 -0.300 3.655 1.055 ;
        RECT 4.395 -0.300 4.695 1.055 ;
        RECT 5.435 -0.300 5.735 0.780 ;
        RECT 6.475 -0.300 6.775 1.120 ;
        RECT 7.515 -0.300 7.815 0.780 ;
        RECT 0.000 -0.300 8.610 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 2.835 2.220 6.255 2.435 ;
        RECT 2.835 0.590 3.135 1.625 ;
        RECT 2.835 2.220 3.135 3.210 ;
        RECT 2.835 1.255 5.445 1.625 ;
        RECT 2.835 2.220 4.175 2.455 ;
        RECT 3.875 0.590 4.175 3.140 ;
        RECT 4.915 0.590 5.215 3.140 ;
        RECT 4.915 0.980 5.445 2.455 ;
        RECT 3.875 1.255 5.445 2.435 ;
        RECT 4.915 2.195 6.255 2.455 ;
        RECT 5.955 0.575 6.255 1.215 ;
        RECT 4.915 0.980 6.255 1.215 ;
        RECT 5.955 2.195 6.255 3.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.705 2.570 1.005 3.990 ;
        RECT 3.355 2.635 3.655 3.990 ;
        RECT 4.395 2.635 4.695 3.990 ;
        RECT 5.435 2.635 5.735 3.990 ;
        RECT 6.475 2.570 6.775 3.990 ;
        RECT 7.515 2.230 7.815 3.990 ;
        RECT 0.000 3.390 8.610 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.480 0.330 2.400 ;
        RECT 0.105 2.100 0.340 2.400 ;
        RECT 0.105 0.480 0.405 1.360 ;
        RECT 0.105 2.200 0.405 2.400 ;
        RECT 1.570 2.040 1.740 2.370 ;
        RECT 0.105 2.200 1.740 2.370 ;
        RECT 1.275 0.535 1.445 1.585 ;
        RECT 1.275 1.405 2.155 1.585 ;
        RECT 1.985 1.405 2.155 2.720 ;
        RECT 1.775 2.550 2.155 2.720 ;
        RECT 1.275 0.535 2.610 0.705 ;
        RECT 2.310 0.535 2.610 0.805 ;
        RECT 1.225 2.570 1.525 3.190 ;
        RECT 1.760 0.885 2.060 1.155 ;
        RECT 1.760 0.985 2.560 1.155 ;
        RECT 2.390 0.985 2.560 3.190 ;
        RECT 1.225 3.020 2.560 3.190 ;
        RECT 2.390 1.825 3.695 1.995 ;
        RECT 6.135 1.825 6.605 1.995 ;
        RECT 6.435 1.825 6.605 2.195 ;
        RECT 6.435 2.025 7.230 2.195 ;
        RECT 7.060 2.025 7.230 3.005 ;
        RECT 6.435 1.300 6.605 1.565 ;
        RECT 5.655 1.395 6.605 1.565 ;
        RECT 6.435 1.300 7.230 1.470 ;
        RECT 6.995 0.560 7.230 1.470 ;
        RECT 7.410 0.960 7.580 1.845 ;
        RECT 6.835 1.670 7.580 1.845 ;
        RECT 7.410 0.960 8.450 1.130 ;
        RECT 8.280 0.960 8.450 2.870 ;
        RECT 8.065 2.230 8.450 2.870 ;
  END 
END INVTSHD6XHT

MACRO INVTSHD5XHT
  CLASS  CORE ;
  FOREIGN INVTSHD5XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.790 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.040 1.390 7.280 2.020 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.540 1.020 2.020 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 -0.300 0.990 1.120 ;
        RECT 2.700 -0.300 2.870 1.120 ;
        RECT 3.675 -0.300 3.975 1.120 ;
        RECT 4.715 -0.300 5.015 0.780 ;
        RECT 5.755 -0.300 6.055 1.180 ;
        RECT 6.795 -0.300 7.095 0.860 ;
        RECT 0.000 -0.300 7.790 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 3.155 0.590 3.455 3.210 ;
        RECT 3.155 1.320 4.495 2.450 ;
        RECT 4.195 0.590 4.495 3.210 ;
        RECT 3.155 2.225 5.535 2.450 ;
        RECT 5.235 0.560 5.535 1.175 ;
        RECT 4.195 0.960 5.535 1.175 ;
        RECT 5.235 2.225 5.535 3.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.705 2.570 1.005 3.990 ;
        RECT 2.700 2.570 2.870 3.990 ;
        RECT 3.675 2.635 3.975 3.990 ;
        RECT 4.715 2.635 5.015 3.990 ;
        RECT 5.755 2.570 6.055 3.990 ;
        RECT 6.795 2.230 7.095 3.990 ;
        RECT 0.000 3.390 7.790 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.480 0.305 2.370 ;
        RECT 0.105 0.480 0.405 1.360 ;
        RECT 1.570 2.000 1.740 2.370 ;
        RECT 0.105 2.200 1.740 2.370 ;
        RECT 1.275 0.640 1.445 1.585 ;
        RECT 1.275 1.415 2.170 1.585 ;
        RECT 1.990 1.415 2.170 2.740 ;
        RECT 1.745 2.570 2.170 2.740 ;
        RECT 1.290 2.570 1.460 3.145 ;
        RECT 1.795 0.595 1.965 1.235 ;
        RECT 1.795 1.065 2.520 1.235 ;
        RECT 2.350 1.065 2.520 3.145 ;
        RECT 1.225 2.975 2.520 3.145 ;
        RECT 4.735 1.875 5.905 2.045 ;
        RECT 5.735 1.875 5.905 2.305 ;
        RECT 5.735 2.135 6.510 2.305 ;
        RECT 6.340 2.135 6.510 3.115 ;
        RECT 6.340 0.720 6.510 1.545 ;
        RECT 4.735 1.375 6.510 1.545 ;
        RECT 6.690 1.040 6.860 1.915 ;
        RECT 6.115 1.745 6.860 1.915 ;
        RECT 7.345 0.820 7.645 1.210 ;
        RECT 6.690 1.040 7.645 1.210 ;
        RECT 7.475 0.820 7.645 2.840 ;
        RECT 7.345 2.200 7.645 2.840 ;
  END 
END INVTSHD5XHT

MACRO INVTSHD4XHT
  CLASS  CORE ;
  FOREIGN INVTSHD4XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.380 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.615 1.475 6.870 2.015 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.675 0.705 2.015 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.705 -0.300 1.005 0.895 ;
        RECT 3.185 -0.300 3.485 0.935 ;
        RECT 4.225 -0.300 4.525 0.935 ;
        RECT 5.265 -0.300 5.565 0.895 ;
        RECT 6.375 -0.300 6.675 0.895 ;
        RECT 0.000 -0.300 7.380 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 2.730 0.720 2.900 1.360 ;
        RECT 2.730 2.150 2.900 3.140 ;
        RECT 2.730 1.190 4.105 1.360 ;
        RECT 3.530 1.190 4.105 2.320 ;
        RECT 2.730 2.150 4.105 2.320 ;
        RECT 3.770 0.720 3.940 3.130 ;
        RECT 3.770 1.145 4.105 2.580 ;
        RECT 3.770 1.145 4.980 1.315 ;
        RECT 3.770 2.410 4.980 2.580 ;
        RECT 4.810 0.675 4.980 1.315 ;
        RECT 2.730 1.190 4.980 1.315 ;
        RECT 4.810 2.410 4.980 3.050 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.705 2.635 1.005 3.990 ;
        RECT 3.185 2.565 3.485 3.990 ;
        RECT 4.225 2.895 4.525 3.990 ;
        RECT 5.265 2.555 5.565 3.990 ;
        RECT 6.375 2.215 6.675 3.990 ;
        RECT 0.000 3.390 7.380 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.480 0.340 1.490 ;
        RECT 0.105 0.480 0.405 0.650 ;
        RECT 0.170 1.320 1.100 1.490 ;
        RECT 0.930 1.320 1.100 2.365 ;
        RECT 0.105 2.195 1.100 2.365 ;
        RECT 0.930 2.115 1.805 2.285 ;
        RECT 1.290 1.015 1.460 1.600 ;
        RECT 1.290 1.430 2.155 1.600 ;
        RECT 1.950 1.430 2.155 1.730 ;
        RECT 1.985 1.430 2.155 2.655 ;
        RECT 1.745 2.485 2.155 2.655 ;
        RECT 1.290 2.715 1.460 3.020 ;
        RECT 1.745 1.080 2.530 1.250 ;
        RECT 2.360 1.080 2.530 3.020 ;
        RECT 1.290 2.835 2.530 3.020 ;
        RECT 4.945 1.845 5.245 2.195 ;
        RECT 4.945 2.025 6.020 2.195 ;
        RECT 5.850 2.025 6.020 3.130 ;
        RECT 5.185 1.125 5.355 1.665 ;
        RECT 4.425 1.495 5.355 1.665 ;
        RECT 5.785 0.785 6.085 1.295 ;
        RECT 5.185 1.125 6.085 1.295 ;
        RECT 6.265 1.125 6.435 1.760 ;
        RECT 5.620 1.590 6.435 1.760 ;
        RECT 7.040 2.150 7.210 2.795 ;
        RECT 7.050 1.125 7.220 2.320 ;
        RECT 7.040 2.150 7.220 2.320 ;
        RECT 6.265 1.125 7.275 1.295 ;
  END 
END INVTSHD4XHT

MACRO INVTSHD3XHT
  CLASS  CORE ;
  FOREIGN INVTSHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.560 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.010 1.520 6.460 2.015 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.310 2.015 ;
        RECT 0.100 1.520 0.520 1.820 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.945 ;
        RECT 2.520 -0.300 2.690 1.340 ;
        RECT 3.495 -0.300 3.795 1.275 ;
        RECT 4.565 -0.300 4.865 1.055 ;
        RECT 6.115 -0.300 6.415 1.295 ;
        RECT 0.000 -0.300 6.560 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 2.970 0.720 3.210 2.815 ;
        RECT 2.970 2.260 4.315 2.430 ;
        RECT 4.080 0.720 4.250 1.625 ;
        RECT 2.970 1.455 4.250 1.625 ;
        RECT 4.015 2.260 4.315 2.770 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.705 2.605 1.005 3.990 ;
        RECT 2.520 2.400 2.690 3.990 ;
        RECT 3.495 2.805 3.795 3.990 ;
        RECT 4.565 2.635 4.865 3.990 ;
        RECT 6.145 2.195 6.445 3.990 ;
        RECT 0.000 3.390 6.560 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 0.915 1.295 ;
        RECT 0.745 1.125 0.915 2.365 ;
        RECT 0.105 2.195 0.915 2.365 ;
        RECT 0.745 1.560 1.110 1.860 ;
        RECT 1.320 1.680 1.490 2.695 ;
        RECT 1.800 1.060 1.970 1.850 ;
        RECT 1.320 1.680 1.970 1.850 ;
        RECT 1.320 2.395 2.320 2.695 ;
        RECT 1.280 0.710 1.450 1.220 ;
        RECT 1.280 0.710 2.340 0.880 ;
        RECT 2.170 0.710 2.340 2.215 ;
        RECT 1.805 2.045 2.340 2.215 ;
        RECT 3.545 1.815 4.185 2.080 ;
        RECT 3.545 1.910 4.715 2.080 ;
        RECT 4.545 1.910 4.715 2.345 ;
        RECT 4.545 2.175 5.320 2.345 ;
        RECT 5.150 2.175 5.320 3.155 ;
        RECT 4.430 1.235 4.600 1.730 ;
        RECT 5.150 0.720 5.320 1.405 ;
        RECT 4.430 1.235 5.320 1.405 ;
        RECT 4.970 1.610 5.830 1.910 ;
        RECT 5.660 1.060 5.830 2.280 ;
  END 
END INVTSHD3XHT

MACRO INVTSHD20XHT
  CLASS  CORE ;
  FOREIGN INVTSHD20XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.550 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 21.185 1.325 21.815 1.845 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.270 1.615 0.585 1.950 ;
        RECT 0.270 1.710 0.995 1.950 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.055 ;
        RECT 1.190 -0.300 1.490 0.805 ;
        RECT 2.230 -0.300 2.530 1.145 ;
        RECT 3.270 -0.300 3.570 1.055 ;
        RECT 6.720 -0.300 7.020 1.055 ;
        RECT 7.760 -0.300 8.060 1.055 ;
        RECT 8.800 -0.300 9.100 1.055 ;
        RECT 9.840 -0.300 10.140 1.055 ;
        RECT 10.880 -0.300 11.180 1.055 ;
        RECT 11.920 -0.300 12.220 1.055 ;
        RECT 12.960 -0.300 13.260 1.055 ;
        RECT 14.000 -0.300 14.300 1.055 ;
        RECT 15.040 -0.300 15.340 1.055 ;
        RECT 16.080 -0.300 16.380 1.055 ;
        RECT 17.770 -0.300 18.070 0.715 ;
        RECT 18.810 -0.300 19.110 0.715 ;
        RECT 19.850 -0.300 20.150 0.715 ;
        RECT 20.890 -0.300 21.190 0.715 ;
        RECT 21.930 -0.300 22.230 1.055 ;
        RECT 0.000 -0.300 22.550 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 6.265 0.720 6.435 2.960 ;
        RECT 7.240 0.785 7.540 2.895 ;
        RECT 8.280 0.785 8.580 2.895 ;
        RECT 9.320 0.785 9.620 2.895 ;
        RECT 10.360 0.785 10.660 2.895 ;
        RECT 11.400 0.785 11.700 2.895 ;
        RECT 12.440 0.785 12.740 2.895 ;
        RECT 13.480 0.765 13.780 2.895 ;
        RECT 14.575 0.785 14.755 2.960 ;
        RECT 14.520 0.785 14.820 2.015 ;
        RECT 15.560 0.765 15.860 2.895 ;
        RECT 6.265 1.370 16.835 2.015 ;
        RECT 16.665 0.720 16.835 2.960 ;
        RECT 16.655 1.370 16.835 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.290 0.405 3.990 ;
        RECT 1.190 2.875 1.490 3.990 ;
        RECT 2.230 2.885 2.530 3.990 ;
        RECT 3.300 3.220 3.600 3.990 ;
        RECT 6.720 2.295 7.020 3.990 ;
        RECT 7.760 2.295 8.060 3.990 ;
        RECT 8.800 2.295 9.100 3.990 ;
        RECT 9.840 2.295 10.140 3.990 ;
        RECT 10.880 2.295 11.180 3.990 ;
        RECT 11.920 2.295 12.220 3.990 ;
        RECT 12.960 2.295 13.260 3.990 ;
        RECT 14.000 2.295 14.300 3.990 ;
        RECT 15.040 2.295 15.340 3.990 ;
        RECT 16.080 2.295 16.380 3.990 ;
        RECT 17.770 2.635 18.070 3.990 ;
        RECT 18.810 2.635 19.110 3.990 ;
        RECT 19.850 2.635 20.150 3.990 ;
        RECT 20.890 2.635 21.190 3.990 ;
        RECT 21.930 2.295 22.230 3.990 ;
        RECT 0.000 3.390 22.550 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.685 0.480 0.875 1.290 ;
        RECT 0.685 2.130 0.875 3.110 ;
        RECT 0.685 1.120 1.090 1.290 ;
        RECT 0.885 1.120 1.090 1.515 ;
        RECT 0.885 1.325 1.445 1.515 ;
        RECT 1.255 1.325 1.445 2.315 ;
        RECT 0.685 2.130 1.445 2.315 ;
        RECT 1.255 1.785 4.475 1.985 ;
        RECT 1.760 0.720 1.960 1.525 ;
        RECT 2.810 0.720 2.990 1.525 ;
        RECT 3.835 0.720 4.015 1.525 ;
        RECT 1.760 1.325 5.075 1.525 ;
        RECT 3.780 2.175 5.075 2.355 ;
        RECT 4.875 1.020 5.075 2.420 ;
        RECT 4.875 1.475 5.715 1.675 ;
        RECT 5.535 1.430 5.715 1.730 ;
        RECT 1.775 2.185 1.945 2.825 ;
        RECT 2.815 2.185 2.985 2.840 ;
        RECT 1.775 2.185 3.480 2.385 ;
        RECT 3.280 2.185 3.480 2.945 ;
        RECT 4.300 0.520 4.600 1.075 ;
        RECT 4.300 0.520 5.640 0.720 ;
        RECT 5.390 2.300 5.590 2.945 ;
        RECT 3.280 2.745 5.590 2.945 ;
        RECT 5.340 0.520 5.640 1.140 ;
        RECT 5.340 0.960 6.075 1.140 ;
        RECT 5.895 0.960 6.075 2.500 ;
        RECT 5.390 2.300 6.075 2.500 ;
        RECT 17.030 1.770 17.210 2.160 ;
        RECT 17.305 1.980 17.505 3.120 ;
        RECT 18.335 1.980 18.535 2.965 ;
        RECT 19.380 1.980 19.580 2.970 ;
        RECT 17.030 1.980 20.605 2.160 ;
        RECT 20.425 1.980 20.605 2.960 ;
        RECT 17.030 1.180 17.210 1.570 ;
        RECT 17.300 0.480 17.500 1.360 ;
        RECT 18.340 0.720 18.540 1.360 ;
        RECT 19.380 0.720 19.580 1.360 ;
        RECT 20.425 0.720 20.605 1.360 ;
        RECT 17.030 1.180 20.605 1.360 ;
        RECT 17.685 1.575 20.985 1.745 ;
        RECT 20.795 0.935 20.985 2.390 ;
        RECT 20.795 2.200 21.660 2.390 ;
        RECT 21.475 0.480 21.645 1.125 ;
        RECT 20.795 0.935 21.645 1.125 ;
        RECT 21.470 2.200 21.660 3.190 ;
  END 
END INVTSHD20XHT

MACRO INVTSHD12XHT
  CLASS  CORE ;
  FOREIGN INVTSHD12XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.940 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 13.100 1.265 13.435 1.875 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.675 0.630 2.055 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.120 ;
        RECT 1.695 -0.300 1.995 1.120 ;
        RECT 4.660 -0.300 4.960 1.055 ;
        RECT 5.700 -0.300 6.000 1.055 ;
        RECT 6.740 -0.300 7.040 1.055 ;
        RECT 7.780 -0.300 8.080 1.055 ;
        RECT 8.820 -0.300 9.120 1.055 ;
        RECT 9.860 -0.300 10.160 1.055 ;
        RECT 11.640 -0.300 11.940 0.715 ;
        RECT 12.680 -0.300 12.980 0.715 ;
        RECT 0.000 -0.300 13.940 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 4.205 0.720 4.375 2.960 ;
        RECT 5.245 0.720 5.415 2.960 ;
        RECT 6.285 0.720 6.455 2.960 ;
        RECT 7.325 0.720 7.495 2.960 ;
        RECT 8.365 0.720 8.535 2.960 ;
        RECT 9.405 0.700 9.575 2.960 ;
        RECT 4.205 1.365 10.615 1.980 ;
        RECT 10.445 0.715 10.615 2.960 ;
        RECT 10.435 1.365 10.615 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.885 0.955 3.990 ;
        RECT 1.695 2.885 1.995 3.990 ;
        RECT 4.660 2.295 4.960 3.990 ;
        RECT 5.700 2.295 6.000 3.990 ;
        RECT 6.740 2.295 7.040 3.990 ;
        RECT 7.780 2.295 8.080 3.990 ;
        RECT 8.820 2.295 9.120 3.990 ;
        RECT 9.860 2.295 10.160 3.990 ;
        RECT 11.640 2.635 11.940 3.990 ;
        RECT 12.680 2.635 12.980 3.990 ;
        RECT 0.000 3.390 13.940 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.900 0.340 1.480 ;
        RECT 0.170 2.295 0.340 2.945 ;
        RECT 0.170 1.300 1.060 1.480 ;
        RECT 0.880 1.300 1.060 2.485 ;
        RECT 0.170 2.295 1.060 2.485 ;
        RECT 0.880 1.825 2.505 2.025 ;
        RECT 1.240 0.655 1.410 1.600 ;
        RECT 1.240 1.400 2.980 1.600 ;
        RECT 1.240 1.430 3.620 1.600 ;
        RECT 2.780 1.060 2.980 2.480 ;
        RECT 2.780 1.430 3.620 1.730 ;
        RECT 1.240 2.225 1.410 2.875 ;
        RECT 1.240 2.225 2.455 2.460 ;
        RECT 2.255 2.225 2.455 3.060 ;
        RECT 2.205 0.520 2.505 1.080 ;
        RECT 2.205 0.520 3.545 0.720 ;
        RECT 3.300 2.420 3.500 3.060 ;
        RECT 2.255 2.855 3.500 3.060 ;
        RECT 3.245 0.520 3.545 1.075 ;
        RECT 3.245 0.895 4.010 1.075 ;
        RECT 3.830 0.895 4.010 2.620 ;
        RECT 3.300 2.420 4.010 2.620 ;
        RECT 10.810 1.770 10.990 2.160 ;
        RECT 11.170 1.980 11.370 2.960 ;
        RECT 10.810 1.980 12.400 2.160 ;
        RECT 12.220 1.980 12.400 2.960 ;
        RECT 10.810 1.215 10.990 1.570 ;
        RECT 11.170 0.720 11.370 1.395 ;
        RECT 12.220 0.720 12.400 1.395 ;
        RECT 10.810 1.215 12.400 1.395 ;
        RECT 11.525 1.575 12.920 1.745 ;
        RECT 12.730 0.915 12.920 2.340 ;
        RECT 12.730 2.165 13.435 2.335 ;
        RECT 13.265 2.165 13.435 3.210 ;
        RECT 13.200 0.545 13.500 1.085 ;
        RECT 12.730 0.915 13.500 1.085 ;
  END 
END INVTSHD12XHT

MACRO INVODHD8XHT
  CLASS  CORE ;
  FOREIGN INVODHD8XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.360 0.405 2.015 ;
    END
  END A
  PIN Z0
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 1.720 0.720 1.955 1.360 ;
    END
  END Z0
  PIN Z1
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 2.150 0.720 2.450 1.360 ;
    END
  END Z1
  PIN Z2
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 3.200 0.720 3.590 1.360 ;
    END
  END Z2
  PIN Z3
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 3.085 2.060 3.385 3.180 ;
        RECT 2.905 2.965 3.385 3.180 ;
    END
  END Z3
  PIN Z4
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 4.130 2.060 4.430 2.815 ;
        RECT 4.130 2.480 4.490 2.815 ;
    END
  END Z4
  PIN Z5
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 1.535 2.060 1.835 2.835 ;
        RECT 1.325 2.495 1.835 2.835 ;
    END
  END Z5
  PIN Z6
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 2.560 2.060 2.885 2.635 ;
    END
  END Z6
  PIN Z7
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 3.790 0.720 4.100 1.360 ;
    END
  END Z7
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.135 0.915 1.525 1.120 ;
        RECT 0.105 -0.300 0.405 1.055 ;
        RECT 1.355 -0.300 1.435 1.865 ;
        RECT 1.135 -0.300 1.435 1.120 ;
        RECT 1.355 0.915 1.525 1.865 ;
        RECT 2.065 1.695 2.365 2.460 ;
        RECT 2.685 -0.300 2.985 1.865 ;
        RECT 3.615 1.695 3.915 2.460 ;
        RECT 4.320 -0.300 4.620 1.865 ;
        RECT 1.355 1.695 4.620 1.865 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.685 0.720 0.875 2.960 ;
        RECT 0.685 1.430 1.165 1.730 ;
  END 
END INVODHD8XHT

MACRO INVHDUXHT
  CLASS  CORE ;
  FOREIGN INVHDUXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.230 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.310 2.015 ;
        RECT 0.100 1.520 0.665 1.820 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.180 -0.300 0.480 1.295 ;
        RECT 0.000 -0.300 1.230 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.845 1.060 1.015 2.430 ;
        RECT 0.845 1.060 1.060 1.605 ;
        RECT 0.845 1.265 1.130 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.180 2.195 0.480 3.990 ;
        RECT 0.000 3.390 1.230 3.990 ;
    END
  END VDD
END INVHDUXHT

MACRO INVHDPXHT
  CLASS  CORE ;
  FOREIGN INVHDPXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.230 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.590 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.190 -0.300 0.490 1.145 ;
        RECT 0.000 -0.300 1.230 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.770 0.720 0.960 2.960 ;
        RECT 0.770 1.265 1.130 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.190 2.515 0.490 3.990 ;
        RECT 0.000 3.390 1.230 3.990 ;
    END
  END VDD
END INVHDPXHT

MACRO INVHD3XHT
  CLASS  CORE ;
  FOREIGN INVHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.610 1.545 1.280 1.950 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.300 -0.300 0.600 1.055 ;
        RECT 1.340 -0.300 1.640 0.715 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.820 0.785 1.120 1.360 ;
        RECT 0.820 2.140 1.120 3.060 ;
        RECT 0.820 1.170 2.160 1.360 ;
        RECT 1.480 1.170 2.160 2.410 ;
        RECT 0.820 2.140 2.160 2.410 ;
        RECT 1.860 0.785 2.160 2.895 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.300 2.295 0.600 3.990 ;
        RECT 1.340 2.635 1.640 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
END INVHD3XHT

MACRO INVHD2XHT
  CLASS  CORE ;
  FOREIGN INVHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.505 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.055 ;
        RECT 1.145 -0.300 1.445 1.055 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.685 0.715 0.875 2.960 ;
        RECT 0.685 1.265 1.130 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 1.145 2.295 1.445 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
END INVHD2XHT

MACRO INVHD16XHT
  CLASS  CORE ;
  FOREIGN INVHD16XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.120 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.445 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.055 ;
        RECT 1.145 -0.300 1.445 1.255 ;
        RECT 2.185 -0.300 2.485 0.715 ;
        RECT 3.225 -0.300 3.525 0.715 ;
        RECT 4.265 -0.300 4.565 0.715 ;
        RECT 5.305 -0.300 5.605 0.715 ;
        RECT 6.345 -0.300 6.645 0.715 ;
        RECT 7.385 -0.300 7.685 0.715 ;
        RECT 8.425 -0.300 8.725 0.715 ;
        RECT 9.465 -0.300 9.765 0.715 ;
        RECT 10.505 -0.300 10.805 0.715 ;
        RECT 11.545 -0.300 11.845 0.715 ;
        RECT 12.585 -0.300 12.885 1.055 ;
        RECT 0.000 -0.300 13.120 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.785 0.785 5.085 1.295 ;
        RECT 4.785 2.045 5.090 2.895 ;
        RECT 5.825 0.785 6.125 1.295 ;
        RECT 5.825 2.045 6.125 2.895 ;
        RECT 6.865 0.785 7.165 1.295 ;
        RECT 6.865 2.045 7.170 2.895 ;
        RECT 7.905 0.785 8.205 1.295 ;
        RECT 7.905 2.045 8.205 2.895 ;
        RECT 4.785 0.940 12.365 1.295 ;
        RECT 8.645 0.940 9.250 2.415 ;
        RECT 4.785 2.045 9.250 2.415 ;
        RECT 8.945 0.785 9.245 2.895 ;
        RECT 8.945 0.940 9.250 2.895 ;
        RECT 9.985 0.785 10.285 2.895 ;
        RECT 11.025 0.785 11.325 2.895 ;
        RECT 11.025 0.940 11.330 2.895 ;
        RECT 8.645 0.940 12.365 2.410 ;
        RECT 4.785 2.045 12.365 2.410 ;
        RECT 12.065 0.785 12.365 2.895 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 1.145 2.365 1.445 3.990 ;
        RECT 2.185 2.635 2.485 3.990 ;
        RECT 3.225 2.635 3.525 3.990 ;
        RECT 4.265 2.635 4.565 3.990 ;
        RECT 5.305 2.635 5.605 3.990 ;
        RECT 6.345 2.635 6.645 3.990 ;
        RECT 7.385 2.635 7.685 3.990 ;
        RECT 8.425 2.635 8.725 3.990 ;
        RECT 9.465 2.635 9.765 3.990 ;
        RECT 10.505 2.635 10.805 3.990 ;
        RECT 11.545 2.635 11.845 3.990 ;
        RECT 12.585 2.295 12.885 3.990 ;
        RECT 0.000 3.390 13.120 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.685 0.720 0.875 2.620 ;
        RECT 0.685 1.585 2.820 1.755 ;
        RECT 1.665 0.785 1.965 1.295 ;
        RECT 1.665 2.045 1.970 2.895 ;
        RECT 1.665 2.045 4.045 2.255 ;
        RECT 2.705 0.785 3.005 1.295 ;
        RECT 2.705 2.045 3.005 2.895 ;
        RECT 1.665 0.940 4.045 1.295 ;
        RECT 3.095 0.940 4.045 2.325 ;
        RECT 2.705 2.045 4.045 2.325 ;
        RECT 3.745 0.825 4.045 2.965 ;
        RECT 3.095 1.580 8.070 1.755 ;
  END 
END INVHD16XHT

MACRO INVHDLXHT
  CLASS  CORE ;
  FOREIGN INVHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.230 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.310 2.015 ;
        RECT 0.100 1.520 0.665 1.820 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.260 -0.300 0.560 1.295 ;
        RECT 0.000 -0.300 1.230 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.845 1.060 1.015 2.310 ;
        RECT 0.845 1.265 1.130 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.180 2.195 0.480 3.990 ;
        RECT 0.000 3.390 1.230 3.990 ;
    END
  END VDD
END INVHDLXHT

MACRO INVHD7XHT
  CLASS  CORE ;
  FOREIGN INVHD7XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.510 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.445 1.645 0.825 1.950 ;
        RECT 0.445 1.645 2.445 1.815 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.120 ;
        RECT 1.145 -0.300 1.445 1.100 ;
        RECT 2.185 -0.300 2.485 1.100 ;
        RECT 3.225 -0.300 3.525 1.100 ;
        RECT 0.000 -0.300 4.510 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.625 0.720 0.925 1.465 ;
        RECT 0.625 2.220 0.925 3.210 ;
        RECT 1.665 0.720 1.965 1.465 ;
        RECT 1.665 2.015 1.965 2.960 ;
        RECT 0.625 1.295 4.045 1.465 ;
        RECT 1.070 2.015 4.045 2.455 ;
        RECT 2.705 0.720 3.005 2.960 ;
        RECT 2.705 1.295 3.015 2.960 ;
        RECT 2.705 1.295 4.045 2.455 ;
        RECT 0.625 2.220 4.045 2.455 ;
        RECT 3.745 0.720 4.045 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.230 0.405 3.990 ;
        RECT 1.145 2.635 1.445 3.990 ;
        RECT 2.185 2.635 2.485 3.990 ;
        RECT 3.225 2.635 3.525 3.990 ;
        RECT 0.000 3.390 4.510 3.990 ;
    END
  END VDD
END INVHD7XHT

MACRO INVHD6XHT
  CLASS  CORE ;
  FOREIGN INVHD6XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.445 1.645 1.430 1.950 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.120 ;
        RECT 1.145 -0.300 1.445 1.110 ;
        RECT 2.185 -0.300 2.485 1.110 ;
        RECT 3.225 -0.300 3.525 1.120 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.625 0.720 0.925 1.460 ;
        RECT 0.625 2.220 0.925 3.210 ;
        RECT 0.625 1.290 3.005 1.460 ;
        RECT 0.625 2.220 1.965 2.455 ;
        RECT 1.665 0.720 1.965 2.960 ;
        RECT 1.665 1.290 3.005 2.450 ;
        RECT 0.625 2.220 3.005 2.450 ;
        RECT 2.705 0.720 3.005 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.230 0.405 3.990 ;
        RECT 1.145 2.635 1.445 3.990 ;
        RECT 2.185 2.630 2.485 3.990 ;
        RECT 3.225 2.230 3.525 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
END INVHD6XHT

MACRO INVHD5XHT
  CLASS  CORE ;
  FOREIGN INVHD5XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.445 1.645 1.455 1.950 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.120 ;
        RECT 1.145 -0.300 1.445 1.110 ;
        RECT 2.185 -0.300 2.485 1.120 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.625 0.720 0.925 1.465 ;
        RECT 0.625 2.130 0.925 3.120 ;
        RECT 0.625 1.295 1.965 1.465 ;
        RECT 0.625 1.305 3.005 1.465 ;
        RECT 1.665 0.720 1.965 2.960 ;
        RECT 1.665 1.305 3.005 2.455 ;
        RECT 0.625 2.130 3.005 2.455 ;
        RECT 2.705 0.720 3.005 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.230 0.405 3.990 ;
        RECT 1.145 2.635 1.445 3.990 ;
        RECT 2.185 2.635 2.485 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
END INVHD5XHT

MACRO INVHD4XHT
  CLASS  CORE ;
  FOREIGN INVHD4XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.435 1.545 1.175 1.950 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.215 -0.300 0.515 1.055 ;
        RECT 1.255 -0.300 1.555 0.715 ;
        RECT 2.295 -0.300 2.595 1.055 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.735 0.785 1.035 1.360 ;
        RECT 0.735 2.140 1.035 3.050 ;
        RECT 0.735 0.940 2.075 1.360 ;
        RECT 1.395 0.940 2.075 2.410 ;
        RECT 0.735 2.140 2.075 2.410 ;
        RECT 1.775 0.785 2.075 2.895 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.215 2.295 0.515 3.990 ;
        RECT 1.255 2.635 1.555 3.990 ;
        RECT 2.295 2.295 2.595 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
END INVHD4XHT

MACRO INVHD1XHT
  CLASS  CORE ;
  FOREIGN INVHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.230 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.605 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.205 -0.300 0.505 1.055 ;
        RECT 0.000 -0.300 1.230 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.785 0.720 0.975 2.960 ;
        RECT 0.785 1.265 1.130 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.205 2.295 0.505 3.990 ;
        RECT 0.000 3.390 1.230 3.990 ;
    END
  END VDD
END INVHD1XHT

MACRO INVHD20XHT
  CLASS  CORE ;
  FOREIGN INVHD20XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.400 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.430 0.505 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.055 ;
        RECT 1.145 -0.300 1.445 1.055 ;
        RECT 2.185 -0.300 2.485 0.715 ;
        RECT 3.225 -0.300 3.525 0.715 ;
        RECT 4.265 -0.300 4.565 0.715 ;
        RECT 5.815 -0.300 6.115 0.715 ;
        RECT 6.855 -0.300 7.155 0.715 ;
        RECT 7.895 -0.300 8.195 0.715 ;
        RECT 8.935 -0.300 9.235 0.715 ;
        RECT 9.975 -0.300 10.275 0.715 ;
        RECT 11.015 -0.300 11.315 0.715 ;
        RECT 12.055 -0.300 12.355 0.715 ;
        RECT 13.095 -0.300 13.395 0.715 ;
        RECT 14.135 -0.300 14.435 0.715 ;
        RECT 15.175 -0.300 15.475 0.715 ;
        RECT 0.000 -0.300 16.400 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.295 0.785 5.595 1.295 ;
        RECT 5.295 2.045 5.595 2.895 ;
        RECT 5.295 2.045 15.995 2.380 ;
        RECT 6.335 0.785 6.635 1.295 ;
        RECT 6.335 2.045 6.640 2.895 ;
        RECT 7.375 0.785 7.675 1.295 ;
        RECT 7.375 2.045 7.675 2.895 ;
        RECT 8.415 0.785 8.715 2.895 ;
        RECT 8.380 0.940 9.755 2.410 ;
        RECT 6.335 2.045 9.755 2.410 ;
        RECT 9.455 0.785 9.755 2.895 ;
        RECT 10.495 0.785 10.795 1.295 ;
        RECT 10.495 2.045 10.795 2.960 ;
        RECT 11.535 0.785 11.835 1.295 ;
        RECT 11.535 2.045 11.835 2.895 ;
        RECT 5.295 0.940 15.995 1.295 ;
        RECT 12.575 0.785 12.875 2.895 ;
        RECT 12.575 0.940 13.915 2.410 ;
        RECT 13.615 0.785 13.915 2.895 ;
        RECT 14.655 0.785 14.955 2.895 ;
        RECT 12.535 0.940 15.995 2.385 ;
        RECT 6.335 2.045 15.995 2.385 ;
        RECT 15.695 0.785 15.995 2.895 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 1.145 2.295 1.445 3.990 ;
        RECT 2.185 2.635 2.485 3.990 ;
        RECT 3.225 2.635 3.525 3.990 ;
        RECT 4.265 2.635 4.565 3.990 ;
        RECT 5.815 2.635 6.115 3.990 ;
        RECT 6.855 2.635 7.155 3.990 ;
        RECT 7.895 2.635 8.195 3.990 ;
        RECT 8.935 2.635 9.235 3.990 ;
        RECT 9.975 2.635 10.275 3.990 ;
        RECT 11.015 2.635 11.315 3.990 ;
        RECT 12.055 2.635 12.355 3.990 ;
        RECT 13.095 2.635 13.395 3.990 ;
        RECT 14.135 2.635 14.435 3.990 ;
        RECT 15.175 2.635 15.475 3.990 ;
        RECT 0.000 3.390 16.400 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.685 0.720 0.875 2.960 ;
        RECT 0.685 1.585 3.365 1.755 ;
        RECT 1.665 0.785 1.965 1.295 ;
        RECT 1.665 2.045 1.970 2.895 ;
        RECT 2.705 0.785 3.005 1.295 ;
        RECT 2.705 2.045 3.005 2.895 ;
        RECT 3.745 0.635 4.045 1.295 ;
        RECT 1.665 0.940 5.085 1.295 ;
        RECT 3.775 0.635 4.045 3.105 ;
        RECT 3.745 2.045 4.045 3.105 ;
        RECT 3.775 0.940 5.085 2.410 ;
        RECT 1.665 2.045 5.085 2.410 ;
        RECT 4.785 0.635 5.085 3.105 ;
        RECT 3.775 1.585 7.880 1.755 ;
        RECT 10.285 1.585 12.195 1.755 ;
  END 
END INVHD20XHT

MACRO INVCLKHDUXHT
  CLASS  CORE ;
  FOREIGN INVCLKHDUXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.230 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.590 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.160 -0.300 0.460 1.295 ;
        RECT 0.000 -0.300 1.230 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.775 1.060 0.945 2.410 ;
        RECT 0.775 1.060 0.975 1.615 ;
        RECT 0.775 1.265 1.130 1.615 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.190 2.285 0.490 3.990 ;
        RECT 0.000 3.390 1.230 3.990 ;
    END
  END VDD
END INVCLKHDUXHT

MACRO INVCLKHDMXHT
  CLASS  CORE ;
  FOREIGN INVCLKHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.230 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.610 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.210 -0.300 0.510 1.235 ;
        RECT 0.000 -0.300 1.230 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.795 1.060 0.965 2.620 ;
        RECT 0.795 1.270 1.130 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.210 2.305 0.510 3.990 ;
        RECT 0.000 3.390 1.230 3.990 ;
    END
  END VDD
END INVCLKHDMXHT

MACRO INVCLKHD8XHT
  CLASS  CORE ;
  FOREIGN INVCLKHD8XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.445 1.585 0.820 1.950 ;
        RECT 0.445 1.585 2.145 1.765 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.000 ;
        RECT 1.145 -0.300 1.445 1.000 ;
        RECT 2.185 -0.300 2.485 1.000 ;
        RECT 3.225 -0.300 3.525 1.000 ;
        RECT 4.265 -0.300 4.565 1.000 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.625 0.990 0.925 1.385 ;
        RECT 0.625 2.130 0.925 2.705 ;
        RECT 1.665 0.990 1.965 1.385 ;
        RECT 1.665 1.965 1.965 3.045 ;
        RECT 0.625 1.200 4.045 1.385 ;
        RECT 1.050 1.965 4.045 2.335 ;
        RECT 2.705 0.990 3.005 3.045 ;
        RECT 2.400 1.200 4.045 2.335 ;
        RECT 0.625 2.130 4.045 2.335 ;
        RECT 3.745 0.990 4.045 3.045 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.395 0.405 3.990 ;
        RECT 1.145 2.535 1.445 3.990 ;
        RECT 2.185 2.535 2.485 3.990 ;
        RECT 3.225 2.535 3.525 3.990 ;
        RECT 4.265 2.195 4.565 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
END INVCLKHD8XHT

MACRO INVCLKHD4XHT
  CLASS  CORE ;
  FOREIGN INVCLKHD4XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.425 1.585 0.810 1.950 ;
        RECT 0.425 1.585 1.520 1.755 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.200 -0.300 0.500 1.000 ;
        RECT 1.240 -0.300 1.540 1.000 ;
        RECT 2.280 -0.300 2.580 1.015 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.720 1.050 1.020 1.385 ;
        RECT 0.720 2.190 1.020 3.105 ;
        RECT 0.720 1.205 2.060 1.385 ;
        RECT 0.720 2.190 2.060 2.410 ;
        RECT 1.760 1.050 2.060 1.385 ;
        RECT 0.720 1.330 2.465 1.385 ;
        RECT 1.780 1.050 2.060 2.895 ;
        RECT 1.760 2.190 2.060 2.895 ;
        RECT 1.780 1.330 2.465 1.540 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.200 2.295 0.500 3.990 ;
        RECT 1.240 2.635 1.540 3.990 ;
        RECT 2.280 2.295 2.580 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
END INVCLKHD4XHT

MACRO INVHD12XHT
  CLASS  CORE ;
  FOREIGN INVHD12XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.430 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.610 0.585 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.055 ;
        RECT 1.665 -0.300 1.965 0.715 ;
        RECT 2.705 -0.300 3.005 1.055 ;
        RECT 3.745 -0.300 4.045 0.715 ;
        RECT 4.785 -0.300 5.085 0.715 ;
        RECT 5.825 -0.300 6.125 0.715 ;
        RECT 6.865 -0.300 7.165 0.715 ;
        RECT 7.905 -0.300 8.205 0.715 ;
        RECT 8.945 -0.300 9.245 1.055 ;
        RECT 0.000 -0.300 9.430 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.225 0.785 3.525 1.295 ;
        RECT 3.225 2.045 3.530 2.895 ;
        RECT 4.265 0.785 4.565 1.295 ;
        RECT 4.265 2.045 4.565 2.895 ;
        RECT 5.305 0.785 5.605 1.295 ;
        RECT 5.305 2.045 5.610 2.895 ;
        RECT 3.225 0.940 8.725 1.295 ;
        RECT 6.345 0.785 6.645 2.895 ;
        RECT 7.385 0.785 7.685 2.895 ;
        RECT 6.160 0.940 8.725 2.410 ;
        RECT 3.225 2.045 8.725 2.410 ;
        RECT 8.425 0.785 8.725 2.895 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.635 0.925 3.990 ;
        RECT 1.665 2.635 1.965 3.990 ;
        RECT 2.705 2.295 3.005 3.990 ;
        RECT 3.745 2.635 4.045 3.990 ;
        RECT 4.785 2.635 5.085 3.990 ;
        RECT 5.825 2.635 6.125 3.990 ;
        RECT 6.865 2.635 7.165 3.990 ;
        RECT 7.905 2.635 8.205 3.990 ;
        RECT 8.945 2.295 9.245 3.990 ;
        RECT 0.000 3.390 9.430 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.720 0.340 1.410 ;
        RECT 0.170 2.230 0.340 3.210 ;
        RECT 0.170 1.240 0.965 1.410 ;
        RECT 0.795 1.240 0.965 2.400 ;
        RECT 0.170 2.230 0.965 2.400 ;
        RECT 0.795 1.610 1.945 1.780 ;
        RECT 1.145 0.785 1.445 1.295 ;
        RECT 1.145 2.040 1.450 2.895 ;
        RECT 1.145 2.040 2.485 2.255 ;
        RECT 2.185 0.785 2.485 1.295 ;
        RECT 1.145 0.940 2.485 1.295 ;
        RECT 2.220 0.785 2.485 2.895 ;
        RECT 2.185 2.040 2.485 2.895 ;
        RECT 2.220 1.555 5.920 1.780 ;
  END 
END INVHD12XHT

MACRO INVCLKHD2XHT
  CLASS  CORE ;
  FOREIGN INVCLKHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.375 0.505 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.095 ;
        RECT 1.145 -0.300 1.445 1.095 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.685 1.060 0.875 2.960 ;
        RECT 0.685 1.325 1.195 1.545 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 1.145 2.295 1.445 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
END INVCLKHD2XHT

MACRO INVCLKHD1XHT
  CLASS  CORE ;
  FOREIGN INVCLKHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.230 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.520 0.590 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.190 -0.300 0.490 1.105 ;
        RECT 0.000 -0.300 1.230 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.770 1.060 0.960 2.960 ;
        RECT 0.770 1.265 1.130 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.190 2.295 0.490 3.990 ;
        RECT 0.000 3.390 1.230 3.990 ;
    END
  END VDD
END INVCLKHD1XHT

MACRO INVCLKHD16XHT
  CLASS  CORE ;
  FOREIGN INVCLKHD16XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.020 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.445 1.675 0.850 1.950 ;
        RECT 0.445 1.675 5.875 1.845 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.050 ;
        RECT 1.145 -0.300 1.445 1.050 ;
        RECT 2.185 -0.300 2.485 1.050 ;
        RECT 3.225 -0.300 3.525 1.050 ;
        RECT 4.265 -0.300 4.565 1.050 ;
        RECT 5.305 -0.300 5.605 1.050 ;
        RECT 6.345 -0.300 6.645 1.050 ;
        RECT 7.385 -0.300 7.685 1.050 ;
        RECT 8.425 -0.300 8.725 1.105 ;
        RECT 0.000 -0.300 9.020 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.625 1.060 0.925 1.495 ;
        RECT 0.625 2.130 0.925 3.095 ;
        RECT 1.665 1.060 1.965 1.495 ;
        RECT 1.665 2.130 1.965 3.095 ;
        RECT 2.705 1.060 3.005 1.495 ;
        RECT 2.705 2.130 3.005 3.095 ;
        RECT 3.745 1.060 4.045 1.495 ;
        RECT 3.745 2.130 4.045 3.095 ;
        RECT 4.785 1.060 5.085 1.495 ;
        RECT 4.785 2.130 5.085 3.095 ;
        RECT 0.625 2.130 8.205 2.400 ;
        RECT 5.825 1.060 6.125 1.495 ;
        RECT 5.825 2.130 6.125 3.095 ;
        RECT 0.625 1.230 8.205 1.495 ;
        RECT 6.865 1.060 7.165 2.895 ;
        RECT 6.370 1.230 8.205 2.410 ;
        RECT 5.825 2.130 8.205 2.410 ;
        RECT 7.905 1.060 8.205 2.895 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.245 0.405 3.990 ;
        RECT 1.145 2.585 1.445 3.990 ;
        RECT 2.185 2.585 2.485 3.990 ;
        RECT 3.225 2.585 3.525 3.990 ;
        RECT 4.265 2.585 4.565 3.990 ;
        RECT 5.305 2.585 5.605 3.990 ;
        RECT 6.345 2.605 6.645 3.990 ;
        RECT 7.385 2.605 7.685 3.990 ;
        RECT 8.425 2.245 8.725 3.990 ;
        RECT 0.000 3.390 9.020 3.990 ;
    END
  END VDD
END INVCLKHD16XHT

MACRO INVCLKHD14XHT
  CLASS  CORE ;
  FOREIGN INVCLKHD14XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.380 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.395 1.675 0.855 1.955 ;
        RECT 0.395 1.675 4.540 1.845 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.160 -0.300 0.460 1.030 ;
        RECT 1.200 -0.300 1.500 1.030 ;
        RECT 2.240 -0.300 2.540 1.030 ;
        RECT 3.280 -0.300 3.580 1.030 ;
        RECT 4.320 -0.300 4.620 1.080 ;
        RECT 5.360 -0.300 5.660 1.080 ;
        RECT 6.400 -0.300 6.700 1.080 ;
        RECT 0.000 -0.300 7.380 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.680 1.060 0.980 1.495 ;
        RECT 0.680 2.145 0.980 2.995 ;
        RECT 1.720 1.060 2.020 1.495 ;
        RECT 1.720 2.145 2.020 2.995 ;
        RECT 2.760 1.060 3.060 1.495 ;
        RECT 2.760 2.145 3.060 2.995 ;
        RECT 3.800 1.060 4.100 1.495 ;
        RECT 0.680 1.210 4.100 1.495 ;
        RECT 3.800 2.145 4.100 2.995 ;
        RECT 0.680 1.305 7.220 1.495 ;
        RECT 4.840 1.060 5.140 2.895 ;
        RECT 4.840 1.305 6.180 2.395 ;
        RECT 0.680 2.145 6.180 2.395 ;
        RECT 5.880 1.060 6.180 2.895 ;
        RECT 4.840 1.305 7.220 2.375 ;
        RECT 0.680 2.145 7.220 2.375 ;
        RECT 6.920 1.060 7.220 2.895 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.160 2.235 0.460 3.990 ;
        RECT 1.200 2.575 1.500 3.990 ;
        RECT 2.240 2.575 2.540 3.990 ;
        RECT 3.280 2.575 3.580 3.990 ;
        RECT 4.320 2.575 4.620 3.990 ;
        RECT 5.360 2.575 5.660 3.990 ;
        RECT 6.400 2.555 6.700 3.990 ;
        RECT 0.000 3.390 7.380 3.990 ;
    END
  END VDD
END INVCLKHD14XHT

MACRO INVCLKHDLXHT
  CLASS  CORE ;
  FOREIGN INVCLKHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.230 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.590 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.190 -0.300 0.490 1.295 ;
        RECT 0.000 -0.300 1.230 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.775 1.055 0.945 2.660 ;
        RECT 0.775 1.265 1.130 1.615 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.190 2.195 0.490 3.990 ;
        RECT 0.000 3.390 1.230 3.990 ;
    END
  END VDD
END INVCLKHDLXHT

MACRO INVCLKHD80XHT
  CLASS  CORE ;
  FOREIGN INVCLKHD80XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 49.200 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.445 1.585 0.785 1.950 ;
        RECT 0.445 1.585 1.765 1.755 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.145 -0.300 1.445 0.990 ;
        RECT 2.185 -0.300 2.485 0.990 ;
        RECT 3.225 -0.300 3.525 0.990 ;
        RECT 4.265 -0.300 4.565 0.990 ;
        RECT 5.305 -0.300 5.605 0.990 ;
        RECT 6.345 -0.300 6.645 0.990 ;
        RECT 7.385 -0.300 7.685 0.990 ;
        RECT 8.425 -0.300 8.725 0.990 ;
        RECT 9.465 -0.300 9.765 0.990 ;
        RECT 10.505 -0.300 10.805 0.990 ;
        RECT 11.545 -0.300 11.845 0.990 ;
        RECT 12.585 -0.300 12.885 0.990 ;
        RECT 13.625 -0.300 13.925 0.990 ;
        RECT 14.665 -0.300 14.965 0.715 ;
        RECT 15.705 -0.300 16.005 0.715 ;
        RECT 16.745 -0.300 17.045 0.715 ;
        RECT 17.785 -0.300 18.085 0.715 ;
        RECT 18.825 -0.300 19.125 0.715 ;
        RECT 19.865 -0.300 20.165 0.715 ;
        RECT 20.905 -0.300 21.205 0.715 ;
        RECT 21.945 -0.300 22.245 0.715 ;
        RECT 22.985 -0.300 23.285 0.715 ;
        RECT 24.025 -0.300 24.325 0.715 ;
        RECT 25.065 -0.300 25.365 0.715 ;
        RECT 26.105 -0.300 26.405 0.715 ;
        RECT 27.145 -0.300 27.445 0.715 ;
        RECT 28.185 -0.300 28.485 0.715 ;
        RECT 29.225 -0.300 29.525 0.715 ;
        RECT 30.265 -0.300 30.565 0.715 ;
        RECT 31.305 -0.300 31.605 0.715 ;
        RECT 32.345 -0.300 32.645 0.715 ;
        RECT 33.385 -0.300 33.685 1.055 ;
        RECT 34.425 -0.300 34.725 1.055 ;
        RECT 35.465 -0.300 35.765 1.055 ;
        RECT 36.505 -0.300 36.805 1.055 ;
        RECT 37.545 -0.300 37.845 1.055 ;
        RECT 38.585 -0.300 38.885 1.055 ;
        RECT 39.655 -0.300 39.955 0.715 ;
        RECT 0.000 -0.300 49.200 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.145 1.235 41.515 1.435 ;
        RECT 14.145 0.780 14.445 1.435 ;
        RECT 14.145 2.045 14.445 2.895 ;
        RECT 15.185 0.780 15.485 1.435 ;
        RECT 15.185 2.045 15.485 2.895 ;
        RECT 16.225 0.780 16.525 1.435 ;
        RECT 16.225 2.045 16.525 2.895 ;
        RECT 17.265 0.785 17.565 1.435 ;
        RECT 17.265 2.045 17.565 2.895 ;
        RECT 18.305 0.785 18.605 1.435 ;
        RECT 18.305 2.045 18.605 2.895 ;
        RECT 19.345 0.785 19.645 1.435 ;
        RECT 19.345 2.045 19.645 2.895 ;
        RECT 20.385 0.785 20.685 1.435 ;
        RECT 20.385 2.045 20.685 2.895 ;
        RECT 21.425 0.785 21.725 1.435 ;
        RECT 21.425 2.045 21.725 2.895 ;
        RECT 22.465 0.785 22.765 1.435 ;
        RECT 22.465 2.045 22.765 2.895 ;
        RECT 23.505 0.785 23.805 1.435 ;
        RECT 23.505 2.045 23.805 2.895 ;
        RECT 24.545 0.780 24.845 1.435 ;
        RECT 24.545 2.045 24.845 2.895 ;
        RECT 25.585 0.785 25.885 1.435 ;
        RECT 25.585 2.045 25.885 2.895 ;
        RECT 26.625 0.785 26.925 1.435 ;
        RECT 26.625 2.045 26.925 2.895 ;
        RECT 27.665 0.775 27.965 1.435 ;
        RECT 27.665 2.045 27.965 2.895 ;
        RECT 28.705 0.785 29.005 1.435 ;
        RECT 28.705 2.045 29.005 2.895 ;
        RECT 29.745 0.785 30.045 1.435 ;
        RECT 29.745 2.045 30.045 2.895 ;
        RECT 30.785 0.785 31.085 1.435 ;
        RECT 30.785 2.045 31.085 2.895 ;
        RECT 31.825 0.785 32.125 2.895 ;
        RECT 31.365 0.895 33.165 2.410 ;
        RECT 14.145 0.895 33.165 1.435 ;
        RECT 32.865 0.785 33.165 2.895 ;
        RECT 33.905 0.785 34.205 2.895 ;
        RECT 34.945 0.785 35.245 2.895 ;
        RECT 35.985 0.785 36.285 2.895 ;
        RECT 37.025 0.785 37.325 2.895 ;
        RECT 38.065 0.775 38.365 2.895 ;
        RECT 39.105 0.785 39.405 2.895 ;
        RECT 31.365 1.235 41.515 2.410 ;
        RECT 40.440 0.560 40.445 2.895 ;
        RECT 40.145 1.235 40.445 2.895 ;
        RECT 40.440 0.560 41.515 2.410 ;
        RECT 14.145 2.045 41.515 2.410 ;
        RECT 41.215 0.560 41.515 3.125 ;
        RECT 42.255 0.560 42.555 3.125 ;
        RECT 43.295 0.560 43.595 3.125 ;
        RECT 44.335 0.560 44.635 3.125 ;
        RECT 45.375 0.560 45.675 3.125 ;
        RECT 46.415 0.560 46.715 3.125 ;
        RECT 47.455 0.560 47.755 3.125 ;
        RECT 40.440 0.560 48.825 1.365 ;
        RECT 14.145 1.235 48.825 1.365 ;
        RECT 48.525 0.560 48.825 3.005 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.425 0.405 3.990 ;
        RECT 1.145 2.765 1.445 3.990 ;
        RECT 2.185 2.765 2.485 3.990 ;
        RECT 3.225 2.115 3.525 3.990 ;
        RECT 4.265 2.635 4.565 3.990 ;
        RECT 5.305 2.635 5.605 3.990 ;
        RECT 6.345 2.635 6.645 3.990 ;
        RECT 7.385 2.635 7.685 3.990 ;
        RECT 8.425 2.635 8.725 3.990 ;
        RECT 9.465 2.635 9.765 3.990 ;
        RECT 10.505 2.635 10.805 3.990 ;
        RECT 11.545 2.635 11.845 3.990 ;
        RECT 12.585 2.635 12.885 3.990 ;
        RECT 13.625 2.295 13.925 3.990 ;
        RECT 14.665 2.635 14.965 3.990 ;
        RECT 15.705 2.635 16.005 3.990 ;
        RECT 16.745 2.635 17.045 3.990 ;
        RECT 17.785 2.635 18.085 3.990 ;
        RECT 18.825 2.635 19.125 3.990 ;
        RECT 19.865 2.635 20.165 3.990 ;
        RECT 20.905 2.635 21.205 3.990 ;
        RECT 21.945 2.635 22.245 3.990 ;
        RECT 22.985 2.635 23.285 3.990 ;
        RECT 24.025 2.635 24.325 3.990 ;
        RECT 25.065 2.635 25.365 3.990 ;
        RECT 26.105 2.635 26.405 3.990 ;
        RECT 27.145 2.635 27.445 3.990 ;
        RECT 28.185 2.635 28.485 3.990 ;
        RECT 29.225 2.635 29.525 3.990 ;
        RECT 30.265 2.635 30.565 3.990 ;
        RECT 31.305 2.635 31.605 3.990 ;
        RECT 32.345 2.635 32.645 3.990 ;
        RECT 33.385 2.635 33.685 3.990 ;
        RECT 34.425 2.635 34.725 3.990 ;
        RECT 35.465 2.635 35.765 3.990 ;
        RECT 36.505 2.635 36.805 3.990 ;
        RECT 37.545 2.635 37.845 3.990 ;
        RECT 38.585 2.635 38.885 3.990 ;
        RECT 39.625 2.635 39.925 3.990 ;
        RECT 40.665 2.635 40.965 3.990 ;
        RECT 41.735 1.615 42.035 3.990 ;
        RECT 42.775 1.615 43.075 3.990 ;
        RECT 43.815 1.615 44.115 3.990 ;
        RECT 44.855 1.615 45.155 3.990 ;
        RECT 45.895 1.615 46.195 3.990 ;
        RECT 46.935 1.615 47.235 3.990 ;
        RECT 47.975 1.615 48.275 3.990 ;
        RECT 0.000 3.390 49.200 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.625 1.000 0.925 1.385 ;
        RECT 0.625 2.140 0.925 2.725 ;
        RECT 1.665 1.000 1.965 1.385 ;
        RECT 1.665 2.140 1.965 2.725 ;
        RECT 0.625 1.215 3.005 1.385 ;
        RECT 2.130 1.215 3.005 2.320 ;
        RECT 0.625 2.140 3.005 2.320 ;
        RECT 2.705 1.000 3.005 2.895 ;
        RECT 2.130 1.675 8.020 1.845 ;
        RECT 3.745 1.070 4.045 1.455 ;
        RECT 3.745 2.170 4.045 3.105 ;
        RECT 4.785 1.070 5.085 1.455 ;
        RECT 4.785 2.170 5.085 3.105 ;
        RECT 5.825 1.070 6.125 1.455 ;
        RECT 5.825 2.170 6.125 3.105 ;
        RECT 6.865 1.070 7.165 1.455 ;
        RECT 6.865 2.170 7.165 3.105 ;
        RECT 7.905 1.070 8.205 1.455 ;
        RECT 7.905 2.170 8.205 3.105 ;
        RECT 3.745 1.215 13.405 1.455 ;
        RECT 8.945 1.070 9.245 2.895 ;
        RECT 9.985 1.070 10.285 2.895 ;
        RECT 11.025 1.070 11.325 2.895 ;
        RECT 12.065 1.070 12.365 2.895 ;
        RECT 8.260 1.215 13.405 2.410 ;
        RECT 3.745 2.170 13.405 2.410 ;
        RECT 13.105 0.930 13.405 2.895 ;
        RECT 8.260 1.655 30.925 1.825 ;
  END 
END INVCLKHD80XHT

MACRO INVCLKHD7XHT
  CLASS  CORE ;
  FOREIGN INVCLKHD7XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.365 1.255 0.865 1.950 ;
        RECT 0.365 1.255 1.765 1.490 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 0.790 ;
        RECT 1.145 -0.300 1.445 0.725 ;
        RECT 2.245 -0.300 2.545 0.725 ;
        RECT 3.285 -0.300 3.585 0.825 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.625 0.740 0.925 1.075 ;
        RECT 0.625 2.220 0.925 3.210 ;
        RECT 1.265 1.810 1.995 2.455 ;
        RECT 0.625 2.220 1.995 2.455 ;
        RECT 1.665 0.740 1.965 1.075 ;
        RECT 1.695 1.810 1.995 3.065 ;
        RECT 0.625 0.905 3.065 1.075 ;
        RECT 1.265 1.810 3.065 2.450 ;
        RECT 2.025 0.905 3.065 2.450 ;
        RECT 0.625 2.220 3.065 2.450 ;
        RECT 2.765 0.655 3.065 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.230 0.405 3.990 ;
        RECT 1.145 2.635 1.445 3.990 ;
        RECT 2.245 2.635 2.545 3.990 ;
        RECT 3.285 2.200 3.585 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
END INVCLKHD7XHT

MACRO INVCLKHD6XHT
  CLASS  CORE ;
  FOREIGN INVCLKHD6XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.445 1.585 0.840 1.950 ;
        RECT 0.445 1.585 2.105 1.755 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 0.980 ;
        RECT 1.145 -0.300 1.445 0.980 ;
        RECT 2.185 -0.300 2.485 0.980 ;
        RECT 3.225 -0.300 3.525 0.980 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.625 0.970 0.925 1.385 ;
        RECT 0.625 2.130 0.925 2.980 ;
        RECT 1.665 0.970 1.965 1.385 ;
        RECT 1.665 2.130 1.965 2.980 ;
        RECT 0.625 1.160 3.005 1.385 ;
        RECT 2.345 1.160 3.005 2.345 ;
        RECT 0.625 2.130 3.005 2.345 ;
        RECT 2.705 0.970 3.005 2.895 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.185 0.405 3.990 ;
        RECT 1.145 2.525 1.445 3.990 ;
        RECT 2.185 2.525 2.485 3.990 ;
        RECT 3.225 2.185 3.525 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
END INVCLKHD6XHT

MACRO INVCLKHD40XHT
  CLASS  CORE ;
  FOREIGN INVCLKHD40XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.420 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.360 1.585 0.910 1.950 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.980 ;
        RECT 1.665 -0.300 1.965 0.980 ;
        RECT 2.705 -0.300 3.005 0.980 ;
        RECT 3.745 -0.300 4.045 0.980 ;
        RECT 4.785 -0.300 5.085 0.980 ;
        RECT 5.825 -0.300 6.125 0.980 ;
        RECT 6.865 -0.300 7.165 1.055 ;
        RECT 7.905 -0.300 8.205 0.715 ;
        RECT 8.945 -0.300 9.245 0.715 ;
        RECT 9.985 -0.300 10.285 0.715 ;
        RECT 11.025 -0.300 11.325 0.715 ;
        RECT 12.065 -0.300 12.365 0.715 ;
        RECT 13.105 -0.300 13.405 0.715 ;
        RECT 14.145 -0.300 14.445 0.715 ;
        RECT 15.185 -0.300 15.485 0.715 ;
        RECT 16.225 -0.300 16.525 0.715 ;
        RECT 17.265 -0.300 17.565 0.715 ;
        RECT 18.305 -0.300 18.605 0.715 ;
        RECT 19.345 -0.300 19.645 0.715 ;
        RECT 20.385 -0.300 20.685 0.715 ;
        RECT 0.000 -0.300 25.420 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.385 1.125 24.325 1.455 ;
        RECT 7.385 0.785 7.685 1.455 ;
        RECT 7.385 2.090 7.685 2.940 ;
        RECT 8.425 0.785 8.725 1.455 ;
        RECT 8.425 2.090 8.725 2.940 ;
        RECT 9.465 0.785 9.765 1.455 ;
        RECT 9.465 2.090 9.765 2.940 ;
        RECT 10.505 0.785 10.805 1.455 ;
        RECT 7.385 0.895 10.805 1.455 ;
        RECT 10.505 2.090 10.805 2.940 ;
        RECT 11.545 0.785 11.845 1.455 ;
        RECT 11.545 2.090 11.845 2.985 ;
        RECT 12.585 0.785 12.885 1.455 ;
        RECT 12.585 2.090 12.885 2.940 ;
        RECT 13.625 0.785 13.925 1.455 ;
        RECT 13.625 2.090 13.925 2.940 ;
        RECT 14.665 0.785 14.965 1.455 ;
        RECT 14.665 2.090 14.965 2.940 ;
        RECT 15.705 0.785 16.005 1.455 ;
        RECT 15.705 2.090 16.005 2.940 ;
        RECT 16.745 0.785 17.045 1.455 ;
        RECT 17.000 0.785 17.045 2.940 ;
        RECT 16.745 2.090 17.045 2.940 ;
        RECT 17.785 0.785 18.085 2.895 ;
        RECT 18.825 0.785 19.125 2.895 ;
        RECT 17.000 0.900 20.165 2.410 ;
        RECT 7.385 0.900 20.165 1.455 ;
        RECT 19.865 0.645 20.165 2.895 ;
        RECT 20.905 1.125 21.205 2.895 ;
        RECT 21.945 0.810 22.245 3.085 ;
        RECT 22.985 0.810 23.285 3.085 ;
        RECT 17.000 1.125 24.325 2.410 ;
        RECT 7.385 2.090 24.325 2.410 ;
        RECT 24.025 0.810 24.325 3.085 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.635 0.925 3.990 ;
        RECT 1.665 2.385 1.965 3.990 ;
        RECT 2.705 2.635 3.005 3.990 ;
        RECT 3.745 2.635 4.045 3.990 ;
        RECT 4.785 2.635 5.085 3.990 ;
        RECT 5.825 2.635 6.125 3.990 ;
        RECT 6.865 2.635 7.165 3.990 ;
        RECT 7.905 2.635 8.205 3.990 ;
        RECT 8.945 2.635 9.245 3.990 ;
        RECT 9.985 2.635 10.285 3.990 ;
        RECT 11.025 2.635 11.325 3.990 ;
        RECT 12.065 2.635 12.365 3.990 ;
        RECT 13.105 2.635 13.405 3.990 ;
        RECT 14.145 2.635 14.445 3.990 ;
        RECT 15.185 2.635 15.485 3.990 ;
        RECT 16.225 2.635 16.525 3.990 ;
        RECT 17.265 2.635 17.565 3.990 ;
        RECT 18.305 2.635 18.605 3.990 ;
        RECT 19.345 2.635 19.645 3.990 ;
        RECT 20.385 2.635 20.685 3.990 ;
        RECT 21.425 2.635 21.725 3.990 ;
        RECT 22.465 2.635 22.765 3.990 ;
        RECT 23.505 2.635 23.805 3.990 ;
        RECT 24.545 2.295 24.845 3.990 ;
        RECT 0.000 3.390 25.420 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.920 0.405 1.385 ;
        RECT 0.105 2.170 0.405 3.105 ;
        RECT 0.105 1.205 1.445 1.385 ;
        RECT 1.145 0.920 1.445 2.410 ;
        RECT 0.105 2.170 1.445 2.410 ;
        RECT 1.145 1.675 4.130 1.845 ;
        RECT 2.185 1.060 2.485 1.475 ;
        RECT 2.185 2.170 2.485 3.105 ;
        RECT 3.225 1.060 3.525 1.475 ;
        RECT 3.225 2.170 3.525 3.105 ;
        RECT 4.265 1.060 4.565 1.475 ;
        RECT 4.265 2.170 4.565 3.105 ;
        RECT 2.185 1.205 6.645 1.475 ;
        RECT 5.305 1.060 5.605 3.105 ;
        RECT 4.720 1.205 6.645 2.410 ;
        RECT 2.185 2.170 6.645 2.410 ;
        RECT 6.345 1.010 6.645 3.105 ;
        RECT 4.720 1.675 16.685 1.845 ;
  END 
END INVCLKHD40XHT

MACRO INVCLKHD30XHT
  CLASS  CORE ;
  FOREIGN INVCLKHD30XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.320 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.495 0.445 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 0.975 ;
        RECT 1.145 -0.300 1.445 0.975 ;
        RECT 2.185 -0.300 2.485 0.975 ;
        RECT 3.225 -0.300 3.525 0.975 ;
        RECT 4.265 -0.300 4.565 0.975 ;
        RECT 5.305 -0.300 5.605 0.975 ;
        RECT 6.345 -0.300 6.645 0.975 ;
        RECT 7.385 -0.300 7.685 0.975 ;
        RECT 8.425 -0.300 8.725 0.975 ;
        RECT 9.465 -0.300 9.765 0.975 ;
        RECT 10.505 -0.300 10.805 0.975 ;
        RECT 11.545 -0.300 11.845 0.975 ;
        RECT 12.585 -0.300 12.885 0.975 ;
        RECT 13.625 -0.300 13.925 0.975 ;
        RECT 14.665 -0.300 14.965 0.975 ;
        RECT 15.705 -0.300 16.005 0.975 ;
        RECT 16.745 -0.300 17.045 0.975 ;
        RECT 17.785 -0.300 18.085 0.975 ;
        RECT 18.825 -0.300 19.125 0.975 ;
        RECT 19.865 -0.300 20.165 0.975 ;
        RECT 20.905 -0.300 21.205 0.975 ;
        RECT 0.000 -0.300 21.320 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.825 1.055 6.125 1.495 ;
        RECT 5.825 2.065 6.125 3.105 ;
        RECT 6.865 1.055 7.165 1.495 ;
        RECT 6.865 2.065 7.165 3.105 ;
        RECT 7.905 1.055 8.205 1.495 ;
        RECT 7.905 2.065 8.205 3.105 ;
        RECT 8.945 1.055 9.245 1.495 ;
        RECT 8.945 2.065 9.245 3.105 ;
        RECT 9.985 1.055 10.285 1.495 ;
        RECT 9.985 2.065 10.285 3.105 ;
        RECT 11.025 1.055 11.325 1.495 ;
        RECT 11.025 2.065 11.325 3.105 ;
        RECT 12.065 1.055 12.365 1.495 ;
        RECT 12.065 2.065 12.365 3.105 ;
        RECT 13.105 1.055 13.405 1.495 ;
        RECT 13.105 2.065 13.405 3.105 ;
        RECT 5.825 1.205 20.685 1.495 ;
        RECT 14.145 1.055 14.445 2.895 ;
        RECT 15.185 1.055 15.485 2.895 ;
        RECT 16.225 1.055 16.525 2.895 ;
        RECT 17.265 1.055 17.565 2.895 ;
        RECT 18.305 1.055 18.605 2.895 ;
        RECT 19.345 1.055 19.645 2.895 ;
        RECT 13.455 1.205 20.685 2.410 ;
        RECT 5.825 2.065 20.685 2.410 ;
        RECT 20.385 0.905 20.685 2.895 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 1.145 2.295 1.445 3.990 ;
        RECT 2.185 2.635 2.485 3.990 ;
        RECT 3.225 2.635 3.525 3.990 ;
        RECT 4.265 2.635 4.565 3.990 ;
        RECT 5.305 2.295 5.605 3.990 ;
        RECT 6.345 2.635 6.645 3.990 ;
        RECT 7.385 2.635 7.685 3.990 ;
        RECT 8.425 2.635 8.725 3.990 ;
        RECT 9.465 2.635 9.765 3.990 ;
        RECT 10.505 2.635 10.805 3.990 ;
        RECT 11.545 2.635 11.845 3.990 ;
        RECT 12.585 2.635 12.885 3.990 ;
        RECT 13.625 2.635 13.925 3.990 ;
        RECT 14.665 2.635 14.965 3.990 ;
        RECT 15.705 2.635 16.005 3.990 ;
        RECT 16.745 2.635 17.045 3.990 ;
        RECT 17.785 2.635 18.085 3.990 ;
        RECT 18.825 2.635 19.125 3.990 ;
        RECT 19.865 2.635 20.165 3.990 ;
        RECT 20.905 2.295 21.205 3.990 ;
        RECT 0.000 3.390 21.320 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 0.960 0.870 2.960 ;
        RECT 0.690 1.630 3.220 1.800 ;
        RECT 1.665 1.055 1.965 1.450 ;
        RECT 1.665 1.985 1.965 2.895 ;
        RECT 2.705 1.055 3.005 1.450 ;
        RECT 2.705 1.985 3.005 2.895 ;
        RECT 3.745 1.055 4.045 1.450 ;
        RECT 1.665 1.205 5.085 1.450 ;
        RECT 3.855 1.055 4.045 2.895 ;
        RECT 3.745 1.985 4.045 2.895 ;
        RECT 3.855 1.205 5.085 2.250 ;
        RECT 4.780 1.055 5.085 2.250 ;
        RECT 1.665 1.985 5.085 2.250 ;
        RECT 4.785 1.055 5.085 3.105 ;
        RECT 3.855 1.675 12.470 1.845 ;
  END 
END INVCLKHD30XHT

MACRO INVCLKHD20XHT
  CLASS  CORE ;
  FOREIGN INVCLKHD20XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.070 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.445 1.675 0.825 1.955 ;
        RECT 0.445 1.675 6.625 1.845 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 0.980 ;
        RECT 1.145 -0.300 1.445 0.980 ;
        RECT 2.185 -0.300 2.485 0.980 ;
        RECT 3.225 -0.300 3.525 0.980 ;
        RECT 4.265 -0.300 4.565 0.980 ;
        RECT 5.305 -0.300 5.605 1.030 ;
        RECT 6.345 -0.300 6.645 1.030 ;
        RECT 7.385 -0.300 7.685 1.030 ;
        RECT 8.425 -0.300 8.725 1.030 ;
        RECT 9.465 -0.300 9.765 1.120 ;
        RECT 10.505 -0.300 10.805 1.120 ;
        RECT 0.000 -0.300 11.070 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.625 1.300 10.285 1.495 ;
        RECT 0.625 1.060 0.925 1.495 ;
        RECT 0.625 2.140 0.925 3.105 ;
        RECT 1.665 1.060 1.965 1.495 ;
        RECT 1.665 2.140 1.965 3.105 ;
        RECT 2.705 1.060 3.005 1.495 ;
        RECT 2.705 2.140 3.005 3.105 ;
        RECT 3.745 1.060 4.045 1.495 ;
        RECT 3.745 2.140 4.045 3.105 ;
        RECT 4.785 1.060 5.085 1.495 ;
        RECT 0.625 1.205 5.085 1.495 ;
        RECT 4.785 2.140 5.085 3.105 ;
        RECT 5.825 1.060 6.125 1.495 ;
        RECT 5.825 2.140 6.125 3.105 ;
        RECT 6.865 1.060 7.165 1.495 ;
        RECT 6.865 2.140 7.165 3.105 ;
        RECT 7.905 1.060 8.205 2.895 ;
        RECT 7.245 1.215 9.245 2.410 ;
        RECT 0.625 1.215 9.245 1.495 ;
        RECT 8.945 1.060 9.245 2.895 ;
        RECT 7.245 1.300 10.285 2.410 ;
        RECT 0.625 2.140 10.285 2.410 ;
        RECT 9.985 1.060 10.285 2.895 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 1.145 2.635 1.445 3.990 ;
        RECT 2.185 2.635 2.485 3.990 ;
        RECT 3.225 2.635 3.525 3.990 ;
        RECT 4.265 2.635 4.565 3.990 ;
        RECT 5.305 2.635 5.605 3.990 ;
        RECT 6.345 2.635 6.645 3.990 ;
        RECT 7.385 2.635 7.685 3.990 ;
        RECT 8.425 2.635 8.725 3.990 ;
        RECT 9.465 2.635 9.765 3.990 ;
        RECT 10.505 2.295 10.805 3.990 ;
        RECT 0.000 3.390 11.070 3.990 ;
    END
  END VDD
END INVCLKHD20XHT

MACRO INVCLKHD10XHT
  CLASS  CORE ;
  FOREIGN INVCLKHD10XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.315 1.585 0.890 1.950 ;
        RECT 0.315 1.585 3.535 1.755 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.175 -0.300 0.475 1.000 ;
        RECT 1.215 -0.300 1.515 1.000 ;
        RECT 2.255 -0.300 2.555 1.000 ;
        RECT 3.295 -0.300 3.595 0.960 ;
        RECT 4.335 -0.300 4.635 0.960 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.695 0.990 0.995 1.385 ;
        RECT 0.695 2.130 0.995 3.065 ;
        RECT 1.735 0.990 2.035 1.385 ;
        RECT 1.735 2.130 2.035 3.065 ;
        RECT 2.775 0.990 3.075 1.385 ;
        RECT 2.775 2.130 3.075 3.065 ;
        RECT 0.695 1.180 5.155 1.385 ;
        RECT 3.750 1.180 5.155 2.375 ;
        RECT 3.815 0.990 4.115 3.065 ;
        RECT 3.815 1.140 5.155 2.375 ;
        RECT 0.695 2.130 5.155 2.375 ;
        RECT 4.855 0.990 5.155 3.065 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.175 2.215 0.475 3.990 ;
        RECT 1.215 2.555 1.515 3.990 ;
        RECT 2.255 2.555 2.555 3.990 ;
        RECT 3.295 2.555 3.595 3.990 ;
        RECT 4.335 2.555 4.635 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
END INVCLKHD10XHT

MACRO HOLDHDHT
  CLASS  CORE ;
  FOREIGN HOLDHDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.750 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION INOUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 2.535 1.540 2.705 ;
        RECT 0.655 1.125 1.540 1.295 ;
        RECT 1.330 2.465 1.540 2.835 ;
        RECT 1.370 1.125 1.540 2.835 ;
        RECT 1.300 2.535 1.540 2.835 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.885 0.955 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.515 0.340 2.280 ;
        RECT 0.170 1.585 1.190 1.755 ;
  END 
END HOLDHDHT

MACRO HAHDMXHT
  CLASS  CORE ;
  FOREIGN HAHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.150 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.495 0.520 2.915 ;
        RECT 2.605 2.525 2.775 2.915 ;
        RECT 0.100 2.745 2.775 2.915 ;
        RECT 2.605 2.525 4.115 2.695 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.190 1.265 3.590 1.820 ;
    END
  END B
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.770 1.060 5.230 1.360 ;
        RECT 5.020 1.060 5.230 2.215 ;
        RECT 4.705 2.045 5.230 2.215 ;
    END
  END S
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.185 ;
        RECT 3.160 -0.300 3.460 0.595 ;
        RECT 5.195 -0.300 5.495 0.595 ;
        RECT 0.000 -0.300 6.150 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 3.095 0.955 3.990 ;
        RECT 3.160 2.880 3.460 3.990 ;
        RECT 4.185 2.870 4.485 3.990 ;
        RECT 5.195 2.925 5.495 3.990 ;
        RECT 0.000 3.390 6.150 3.990 ;
    END
  END VDD
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.810 1.060 6.055 2.435 ;
    END
  END CO
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.375 1.755 ;
        RECT 1.205 1.585 1.375 2.565 ;
        RECT 2.165 0.950 2.335 2.565 ;
        RECT 1.205 2.395 2.335 2.565 ;
        RECT 2.515 1.125 2.685 2.215 ;
        RECT 2.515 1.125 2.910 1.295 ;
        RECT 2.515 2.045 2.910 2.215 ;
        RECT 1.640 0.600 1.810 2.215 ;
        RECT 1.575 2.045 1.875 2.215 ;
        RECT 1.640 0.600 2.695 0.770 ;
        RECT 2.525 0.600 2.695 0.945 ;
        RECT 3.665 0.705 3.885 0.945 ;
        RECT 2.525 0.775 3.885 0.945 ;
        RECT 3.665 0.705 4.590 0.875 ;
        RECT 4.420 0.705 4.590 1.840 ;
        RECT 4.420 1.540 4.835 1.840 ;
        RECT 4.070 1.060 4.240 2.215 ;
        RECT 3.635 2.045 4.520 2.215 ;
        RECT 4.350 2.045 4.520 2.620 ;
        RECT 5.460 1.520 5.630 2.620 ;
        RECT 4.350 2.450 5.630 2.620 ;
  END 
END HAHDMXHT

MACRO FILLERC6HDHT
  CLASS  CORE ;
  FOREIGN FILLERC6HDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.160 -0.300 2.300 0.595 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.160 0.865 2.300 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
END FILLERC6HDHT

MACRO FILLERC3HDHT
  CLASS  CORE ;
  FOREIGN FILLERC3HDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.230 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 -0.300 1.100 1.665 ;
        RECT 0.000 -0.300 1.230 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 1.980 1.100 3.990 ;
        RECT 0.000 3.390 1.230 3.990 ;
    END
  END VDD
END FILLERC3HDHT

MACRO HAHDLXHT
  CLASS  CORE ;
  FOREIGN HAHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.150 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.495 0.475 2.915 ;
        RECT 2.605 2.525 2.775 2.915 ;
        RECT 0.100 2.745 2.775 2.915 ;
        RECT 2.605 2.525 4.115 2.695 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.190 1.265 3.590 1.820 ;
    END
  END B
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.770 1.060 5.230 1.360 ;
        RECT 5.020 1.060 5.230 2.215 ;
        RECT 4.705 2.045 5.230 2.215 ;
    END
  END S
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.185 ;
        RECT 3.160 -0.300 3.460 0.595 ;
        RECT 5.195 -0.300 5.495 0.745 ;
        RECT 0.000 -0.300 6.150 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 3.095 0.955 3.990 ;
        RECT 3.160 2.880 3.460 3.990 ;
        RECT 4.185 2.870 4.485 3.990 ;
        RECT 5.195 2.800 5.495 3.990 ;
        RECT 0.000 3.390 6.150 3.990 ;
    END
  END VDD
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.810 1.060 6.055 2.435 ;
    END
  END CO
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.375 1.755 ;
        RECT 1.205 1.585 1.375 2.565 ;
        RECT 2.165 0.950 2.335 2.565 ;
        RECT 1.205 2.395 2.335 2.565 ;
        RECT 2.515 1.125 2.685 2.215 ;
        RECT 2.515 1.125 2.910 1.295 ;
        RECT 2.515 2.045 2.910 2.215 ;
        RECT 1.640 0.600 1.810 2.215 ;
        RECT 1.575 2.045 1.875 2.215 ;
        RECT 1.640 0.600 2.695 0.770 ;
        RECT 2.525 0.600 2.695 0.945 ;
        RECT 3.665 0.705 3.885 0.945 ;
        RECT 2.525 0.775 3.885 0.945 ;
        RECT 3.665 0.705 4.590 0.875 ;
        RECT 4.420 0.705 4.590 1.840 ;
        RECT 4.420 1.540 4.835 1.840 ;
        RECT 4.070 1.060 4.240 2.215 ;
        RECT 3.635 2.045 4.520 2.215 ;
        RECT 4.350 2.045 4.520 2.620 ;
        RECT 5.460 1.520 5.630 2.620 ;
        RECT 4.350 2.450 5.630 2.620 ;
  END 
END HAHDLXHT

MACRO FILLERC8HDHT
  CLASS  CORE ;
  FOREIGN FILLERC8HDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.365 -0.300 2.925 0.595 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.365 0.865 2.925 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
END FILLERC8HDHT

MACRO FILLERC64HDHT
  CLASS  CORE ;
  FOREIGN FILLERC64HDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.240 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.435 -0.300 25.805 0.645 ;
        RECT 0.000 -0.300 26.240 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.435 0.865 25.805 3.990 ;
        RECT 0.000 3.390 26.240 3.990 ;
    END
  END VDD
END FILLERC64HDHT

MACRO FILLERC4HDHT
  CLASS  CORE ;
  FOREIGN FILLERC4HDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 -0.300 1.510 1.595 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 1.980 1.510 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
END FILLERC4HDHT

MACRO FILLERC32HDHT
  CLASS  CORE ;
  FOREIGN FILLERC32HDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.120 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.470 -0.300 12.650 0.620 ;
        RECT 0.000 -0.300 13.120 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.470 0.865 12.650 3.990 ;
        RECT 0.000 3.390 13.120 3.990 ;
    END
  END VDD
END FILLERC32HDHT

MACRO FILLERC1HDHT
  CLASS  CORE ;
  FOREIGN FILLERC1HDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.410 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 -0.300 0.410 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 3.390 0.410 3.990 ;
    END
  END VDD
END FILLERC1HDHT

MACRO FILLER1HDHT
  CLASS  CORE ;
  FOREIGN FILLER1HDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.410 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 -0.300 0.410 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 3.390 0.410 3.990 ;
    END
  END VDD
END FILLER1HDHT

MACRO FILLERC16HDHT
  CLASS  CORE ;
  FOREIGN FILLERC16HDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.560 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.355 -0.300 6.205 0.595 ;
        RECT 0.000 -0.300 6.560 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.355 0.865 6.205 3.990 ;
        RECT 0.000 3.390 6.560 3.990 ;
    END
  END VDD
END FILLERC16HDHT

MACRO HAHD1XHT
  CLASS  CORE ;
  FOREIGN HAHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.150 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.495 0.475 2.915 ;
        RECT 3.880 2.450 4.050 2.915 ;
        RECT 0.100 2.745 4.050 2.915 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.195 1.260 3.590 1.820 ;
    END
  END B
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.770 0.720 4.940 1.360 ;
        RECT 4.770 1.190 5.230 1.360 ;
        RECT 5.020 1.190 5.230 2.215 ;
        RECT 4.705 2.045 5.230 2.215 ;
    END
  END S
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.155 ;
        RECT 3.160 -0.300 3.460 0.595 ;
        RECT 5.225 -0.300 5.525 0.715 ;
        RECT 0.000 -0.300 6.150 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 3.095 0.955 3.990 ;
        RECT 3.160 3.095 3.460 3.990 ;
        RECT 4.250 2.835 4.425 3.990 ;
        RECT 5.225 2.975 5.525 3.990 ;
        RECT 0.000 3.390 6.150 3.990 ;
    END
  END VDD
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.810 0.720 6.050 2.960 ;
    END
  END CO
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.180 1.755 ;
        RECT 1.010 1.585 1.180 2.565 ;
        RECT 2.165 0.950 2.335 2.565 ;
        RECT 1.010 2.395 2.335 2.565 ;
        RECT 2.515 1.125 2.685 2.215 ;
        RECT 2.515 1.125 2.910 1.295 ;
        RECT 2.515 2.045 2.910 2.215 ;
        RECT 1.640 0.600 1.810 2.215 ;
        RECT 1.575 2.045 1.875 2.215 ;
        RECT 1.640 0.600 2.695 0.770 ;
        RECT 2.525 0.600 2.695 0.945 ;
        RECT 3.675 0.680 3.885 0.945 ;
        RECT 2.525 0.775 3.885 0.945 ;
        RECT 3.675 0.680 4.590 0.850 ;
        RECT 4.420 0.680 4.590 1.840 ;
        RECT 4.420 1.540 4.835 1.840 ;
        RECT 4.070 1.060 4.240 2.215 ;
        RECT 3.635 2.045 4.525 2.215 ;
        RECT 4.355 2.045 4.525 2.620 ;
        RECT 5.460 1.520 5.630 2.620 ;
        RECT 4.355 2.450 5.630 2.620 ;
  END 
END HAHD1XHT

MACRO FILLER8HDHT
  CLASS  CORE ;
  FOREIGN FILLER8HDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
END FILLER8HDHT

MACRO FILLER6HDHT
  CLASS  CORE ;
  FOREIGN FILLER6HDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
END FILLER6HDHT

MACRO FILLER4HDHT
  CLASS  CORE ;
  FOREIGN FILLER4HDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
END FILLER4HDHT

MACRO FILLER3HDHT
  CLASS  CORE ;
  FOREIGN FILLER3HDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.230 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 -0.300 1.230 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 3.390 1.230 3.990 ;
    END
  END VDD
END FILLER3HDHT

MACRO FILLER2HDHT
  CLASS  CORE ;
  FOREIGN FILLER2HDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.820 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 -0.300 0.820 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 3.390 0.820 3.990 ;
    END
  END VDD
END FILLER2HDHT

MACRO FILLER16HDHT
  CLASS  CORE ;
  FOREIGN FILLER16HDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.560 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 -0.300 6.560 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 3.390 6.560 3.990 ;
    END
  END VDD
END FILLER16HDHT

MACRO FFSEDQHDMXHT
  CLASS  CORE ;
  FOREIGN FFSEDQHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.760 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.420 1.060 14.660 1.360 ;
        RECT 14.450 1.060 14.660 2.280 ;
        RECT 14.420 1.980 14.660 2.280 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 1.325 1.220 1.925 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.625 0.620 2.010 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.835 1.470 3.205 2.020 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.765 -0.300 1.065 0.795 ;
        RECT 2.580 -0.300 2.880 0.570 ;
        RECT 3.640 -0.300 3.940 0.570 ;
        RECT 5.410 -0.300 5.710 0.570 ;
        RECT 6.860 -0.300 7.160 0.520 ;
        RECT 8.165 -0.300 8.335 0.730 ;
        RECT 9.970 -0.300 10.270 0.525 ;
        RECT 10.950 -0.300 11.250 0.565 ;
        RECT 12.760 -0.300 13.060 0.470 ;
        RECT 13.835 -0.300 14.135 1.145 ;
        RECT 0.000 -0.300 14.760 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 6.345 1.525 6.870 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.665 1.465 6.050 2.010 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.755 2.575 1.055 3.990 ;
        RECT 2.655 2.910 2.955 3.990 ;
        RECT 3.520 2.910 3.820 3.990 ;
        RECT 5.410 2.890 5.710 3.990 ;
        RECT 6.810 3.160 7.110 3.990 ;
        RECT 8.045 2.810 8.215 3.990 ;
        RECT 10.090 3.160 10.390 3.990 ;
        RECT 10.950 3.160 11.250 3.990 ;
        RECT 12.850 2.745 13.150 3.990 ;
        RECT 13.805 2.745 14.105 3.990 ;
        RECT 0.000 3.390 14.760 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.270 0.975 0.440 1.345 ;
        RECT 0.205 2.205 0.505 2.430 ;
        RECT 0.270 0.975 1.600 1.145 ;
        RECT 1.430 0.975 1.600 2.375 ;
        RECT 0.205 2.205 1.600 2.375 ;
        RECT 1.430 1.705 1.700 2.005 ;
        RECT 1.780 1.045 2.050 1.345 ;
        RECT 1.880 1.045 2.050 2.730 ;
        RECT 1.780 2.215 2.050 2.730 ;
        RECT 3.805 1.775 3.975 2.730 ;
        RECT 1.780 2.550 3.975 2.730 ;
        RECT 3.430 1.110 3.600 2.370 ;
        RECT 3.130 2.200 3.600 2.370 ;
        RECT 3.130 1.110 4.280 1.280 ;
        RECT 4.110 1.110 4.280 1.650 ;
        RECT 4.165 1.480 4.335 3.060 ;
        RECT 4.110 1.480 4.520 1.650 ;
        RECT 4.165 2.890 5.020 3.060 ;
        RECT 5.215 1.110 5.385 2.360 ;
        RECT 5.215 1.110 6.140 1.280 ;
        RECT 5.215 2.190 6.140 2.360 ;
        RECT 4.515 1.890 4.685 2.710 ;
        RECT 4.460 1.110 4.870 1.280 ;
        RECT 4.700 1.110 4.870 2.070 ;
        RECT 4.515 1.890 4.870 2.070 ;
        RECT 4.515 2.540 6.345 2.710 ;
        RECT 6.175 2.540 6.345 2.980 ;
        RECT 6.175 2.810 7.845 2.980 ;
        RECT 7.675 2.810 7.845 3.110 ;
        RECT 9.205 0.955 9.375 2.280 ;
        RECT 9.140 0.955 9.440 1.125 ;
        RECT 9.205 1.675 10.640 1.845 ;
        RECT 10.550 1.125 10.850 1.495 ;
        RECT 9.860 1.325 11.360 1.495 ;
        RECT 11.190 1.325 11.360 2.215 ;
        RECT 10.520 2.045 11.360 2.215 ;
        RECT 6.350 1.125 7.220 1.295 ;
        RECT 6.350 2.190 7.220 2.360 ;
        RECT 7.050 1.125 7.220 2.630 ;
        RECT 7.050 1.525 7.275 1.825 ;
        RECT 7.050 2.460 8.655 2.630 ;
        RECT 8.485 2.460 8.655 2.980 ;
        RECT 8.485 2.810 11.830 2.980 ;
        RECT 7.455 1.060 7.625 2.280 ;
        RECT 7.455 1.325 8.190 1.495 ;
        RECT 7.455 2.110 9.005 2.280 ;
        RECT 8.835 1.655 9.005 2.630 ;
        RECT 11.540 1.310 11.710 2.630 ;
        RECT 11.540 1.310 11.940 1.480 ;
        RECT 8.835 2.460 12.345 2.630 ;
        RECT 12.175 2.460 12.345 2.945 ;
        RECT 2.470 0.750 2.640 1.820 ;
        RECT 6.845 0.700 7.015 0.930 ;
        RECT 2.470 0.750 7.015 0.930 ;
        RECT 6.845 0.700 7.985 0.880 ;
        RECT 7.805 0.700 7.985 1.090 ;
        RECT 7.805 0.910 8.485 1.090 ;
        RECT 8.880 0.595 9.655 0.775 ;
        RECT 9.950 0.765 11.550 0.945 ;
        RECT 11.810 0.575 12.370 0.760 ;
        RECT 12.430 0.575 12.445 0.820 ;
        RECT 12.520 0.650 12.750 0.820 ;
        RECT 12.580 0.650 12.750 1.480 ;
        RECT 12.580 1.310 13.705 1.480 ;
        RECT 13.375 0.875 13.545 1.480 ;
        RECT 13.535 1.310 13.705 2.215 ;
        RECT 13.280 2.045 13.705 2.215 ;
        RECT 12.445 0.585 12.455 0.819 ;
        RECT 12.455 0.595 12.465 0.819 ;
        RECT 12.465 0.605 12.475 0.819 ;
        RECT 12.475 0.615 12.485 0.819 ;
        RECT 12.485 0.625 12.495 0.819 ;
        RECT 12.495 0.635 12.505 0.819 ;
        RECT 12.505 0.645 12.515 0.819 ;
        RECT 12.515 0.650 12.521 0.820 ;
        RECT 12.370 0.575 12.380 0.759 ;
        RECT 12.380 0.575 12.390 0.769 ;
        RECT 12.390 0.575 12.400 0.779 ;
        RECT 12.400 0.575 12.410 0.789 ;
        RECT 12.410 0.575 12.420 0.799 ;
        RECT 12.420 0.575 12.430 0.809 ;
        RECT 11.740 0.575 11.750 0.819 ;
        RECT 11.750 0.575 11.760 0.809 ;
        RECT 11.760 0.575 11.770 0.799 ;
        RECT 11.770 0.575 11.780 0.789 ;
        RECT 11.780 0.575 11.790 0.779 ;
        RECT 11.790 0.575 11.800 0.769 ;
        RECT 11.800 0.575 11.810 0.759 ;
        RECT 11.625 0.690 11.635 0.934 ;
        RECT 11.635 0.680 11.645 0.924 ;
        RECT 11.645 0.670 11.655 0.914 ;
        RECT 11.655 0.660 11.665 0.904 ;
        RECT 11.665 0.650 11.675 0.894 ;
        RECT 11.675 0.640 11.685 0.884 ;
        RECT 11.685 0.630 11.695 0.874 ;
        RECT 11.695 0.620 11.705 0.864 ;
        RECT 11.705 0.610 11.715 0.854 ;
        RECT 11.715 0.600 11.725 0.844 ;
        RECT 11.725 0.590 11.735 0.834 ;
        RECT 11.735 0.580 11.741 0.830 ;
        RECT 11.550 0.765 11.560 0.945 ;
        RECT 11.560 0.755 11.570 0.945 ;
        RECT 11.570 0.745 11.580 0.945 ;
        RECT 11.580 0.735 11.590 0.945 ;
        RECT 11.590 0.725 11.600 0.945 ;
        RECT 11.600 0.715 11.610 0.945 ;
        RECT 11.610 0.705 11.620 0.945 ;
        RECT 11.620 0.695 11.626 0.945 ;
        RECT 9.825 0.650 9.835 0.944 ;
        RECT 9.835 0.660 9.845 0.944 ;
        RECT 9.845 0.670 9.855 0.944 ;
        RECT 9.855 0.680 9.865 0.944 ;
        RECT 9.865 0.690 9.875 0.944 ;
        RECT 9.875 0.700 9.885 0.944 ;
        RECT 9.885 0.710 9.895 0.944 ;
        RECT 9.895 0.720 9.905 0.944 ;
        RECT 9.905 0.730 9.915 0.944 ;
        RECT 9.915 0.740 9.925 0.944 ;
        RECT 9.925 0.750 9.935 0.944 ;
        RECT 9.935 0.760 9.945 0.944 ;
        RECT 9.945 0.765 9.951 0.945 ;
        RECT 9.780 0.605 9.790 0.899 ;
        RECT 9.790 0.615 9.800 0.909 ;
        RECT 9.800 0.625 9.810 0.919 ;
        RECT 9.810 0.635 9.820 0.929 ;
        RECT 9.820 0.640 9.826 0.940 ;
        RECT 9.655 0.595 9.665 0.775 ;
        RECT 9.665 0.595 9.675 0.785 ;
        RECT 9.675 0.595 9.685 0.795 ;
        RECT 9.685 0.595 9.695 0.805 ;
        RECT 9.695 0.595 9.705 0.815 ;
        RECT 9.705 0.595 9.715 0.825 ;
        RECT 9.715 0.595 9.725 0.835 ;
        RECT 9.725 0.595 9.735 0.845 ;
        RECT 9.735 0.595 9.745 0.855 ;
        RECT 9.745 0.595 9.755 0.865 ;
        RECT 9.755 0.595 9.765 0.875 ;
        RECT 9.765 0.595 9.775 0.885 ;
        RECT 9.775 0.595 9.781 0.895 ;
        RECT 8.800 0.595 8.810 0.845 ;
        RECT 8.810 0.595 8.820 0.835 ;
        RECT 8.820 0.595 8.830 0.825 ;
        RECT 8.830 0.595 8.840 0.815 ;
        RECT 8.840 0.595 8.850 0.805 ;
        RECT 8.850 0.595 8.860 0.795 ;
        RECT 8.860 0.595 8.870 0.785 ;
        RECT 8.870 0.595 8.880 0.775 ;
        RECT 8.565 0.830 8.575 1.080 ;
        RECT 8.575 0.820 8.585 1.070 ;
        RECT 8.585 0.810 8.595 1.060 ;
        RECT 8.595 0.800 8.605 1.050 ;
        RECT 8.605 0.790 8.615 1.040 ;
        RECT 8.615 0.780 8.625 1.030 ;
        RECT 8.625 0.770 8.635 1.020 ;
        RECT 8.635 0.760 8.645 1.010 ;
        RECT 8.645 0.750 8.655 1.000 ;
        RECT 8.655 0.740 8.665 0.990 ;
        RECT 8.665 0.730 8.675 0.980 ;
        RECT 8.675 0.720 8.685 0.970 ;
        RECT 8.685 0.710 8.695 0.960 ;
        RECT 8.695 0.700 8.705 0.950 ;
        RECT 8.705 0.690 8.715 0.940 ;
        RECT 8.715 0.680 8.725 0.930 ;
        RECT 8.725 0.670 8.735 0.920 ;
        RECT 8.735 0.660 8.745 0.910 ;
        RECT 8.745 0.650 8.755 0.900 ;
        RECT 8.755 0.640 8.765 0.890 ;
        RECT 8.765 0.630 8.775 0.880 ;
        RECT 8.775 0.620 8.785 0.870 ;
        RECT 8.785 0.610 8.795 0.860 ;
        RECT 8.795 0.600 8.801 0.854 ;
        RECT 8.485 0.910 8.495 1.090 ;
        RECT 8.495 0.900 8.505 1.090 ;
        RECT 8.505 0.890 8.515 1.090 ;
        RECT 8.515 0.880 8.525 1.090 ;
        RECT 8.525 0.870 8.535 1.090 ;
        RECT 8.535 0.860 8.545 1.090 ;
        RECT 8.545 0.850 8.555 1.090 ;
        RECT 8.555 0.840 8.565 1.090 ;
        RECT 11.890 0.940 12.190 1.110 ;
        RECT 12.090 1.040 12.290 1.120 ;
        RECT 12.100 1.040 12.290 1.130 ;
        RECT 12.110 1.040 12.290 1.140 ;
        RECT 11.890 2.045 12.190 2.215 ;
        RECT 11.890 0.950 12.200 1.110 ;
        RECT 11.890 0.960 12.210 1.110 ;
        RECT 11.890 0.970 12.220 1.110 ;
        RECT 11.890 0.980 12.230 1.110 ;
        RECT 11.890 0.990 12.240 1.110 ;
        RECT 11.890 1.000 12.250 1.110 ;
        RECT 11.890 1.010 12.260 1.110 ;
        RECT 11.890 1.020 12.270 1.110 ;
        RECT 11.890 1.030 12.280 1.110 ;
        RECT 12.120 1.040 12.290 2.214 ;
        RECT 12.930 1.675 13.100 2.565 ;
        RECT 12.120 1.675 13.355 1.845 ;
        RECT 14.070 1.520 14.240 2.565 ;
        RECT 12.930 2.395 14.240 2.565 ;
        RECT 14.070 1.520 14.260 1.820 ;
  END 
END FFSEDQHDMXHT

MACRO FFSEDQHDLXHT
  CLASS  CORE ;
  FOREIGN FFSEDQHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.760 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.420 1.060 14.660 1.360 ;
        RECT 14.450 1.060 14.660 2.280 ;
        RECT 14.420 1.980 14.660 2.280 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 1.325 1.220 1.945 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.605 0.620 2.010 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.845 1.495 3.205 2.020 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.765 -0.300 1.065 0.795 ;
        RECT 2.570 -0.300 2.870 0.570 ;
        RECT 3.640 -0.300 3.940 0.570 ;
        RECT 5.410 -0.300 5.710 0.570 ;
        RECT 6.810 -0.300 7.110 0.520 ;
        RECT 8.165 -0.300 8.335 0.730 ;
        RECT 9.970 -0.300 10.270 0.525 ;
        RECT 10.940 -0.300 11.240 0.565 ;
        RECT 12.730 -0.300 13.030 0.470 ;
        RECT 13.900 -0.300 14.070 1.360 ;
        RECT 0.000 -0.300 14.760 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 6.345 1.525 6.870 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.665 1.465 6.050 2.010 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.765 2.575 1.065 3.990 ;
        RECT 2.655 2.910 2.955 3.990 ;
        RECT 3.520 2.910 3.820 3.990 ;
        RECT 5.410 2.890 5.710 3.990 ;
        RECT 6.810 3.160 7.110 3.990 ;
        RECT 8.045 2.810 8.215 3.990 ;
        RECT 10.090 3.160 10.390 3.990 ;
        RECT 10.940 3.160 11.240 3.990 ;
        RECT 12.850 2.745 13.150 3.990 ;
        RECT 13.805 2.745 14.105 3.990 ;
        RECT 0.000 3.390 14.760 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.270 0.975 0.440 1.345 ;
        RECT 0.270 0.975 1.600 1.145 ;
        RECT 1.430 0.975 1.600 2.375 ;
        RECT 0.205 2.205 1.600 2.375 ;
        RECT 1.430 1.705 1.700 2.005 ;
        RECT 1.790 0.575 2.050 0.875 ;
        RECT 1.880 0.575 2.050 2.730 ;
        RECT 1.780 2.215 2.050 2.730 ;
        RECT 3.805 1.775 3.975 2.730 ;
        RECT 1.780 2.550 3.975 2.730 ;
        RECT 3.430 1.110 3.600 2.370 ;
        RECT 3.130 2.200 3.600 2.370 ;
        RECT 3.120 1.110 4.280 1.280 ;
        RECT 4.110 1.110 4.280 1.650 ;
        RECT 4.165 1.480 4.335 3.060 ;
        RECT 4.110 1.480 4.520 1.650 ;
        RECT 4.165 2.890 4.970 3.060 ;
        RECT 5.215 1.110 5.385 2.360 ;
        RECT 5.215 1.110 6.140 1.280 ;
        RECT 5.215 2.190 6.140 2.360 ;
        RECT 4.515 1.890 4.685 2.710 ;
        RECT 4.460 1.110 4.870 1.280 ;
        RECT 4.700 1.110 4.870 2.070 ;
        RECT 4.515 1.890 4.870 2.070 ;
        RECT 4.515 2.540 6.425 2.710 ;
        RECT 6.255 2.540 6.425 2.980 ;
        RECT 6.255 2.810 7.845 2.980 ;
        RECT 7.675 2.810 7.845 3.110 ;
        RECT 9.205 0.955 9.375 2.280 ;
        RECT 9.140 0.955 9.440 1.125 ;
        RECT 9.205 1.675 10.640 1.845 ;
        RECT 10.550 1.125 10.850 1.495 ;
        RECT 9.860 1.325 11.360 1.495 ;
        RECT 11.190 1.325 11.360 2.215 ;
        RECT 10.520 2.045 11.360 2.215 ;
        RECT 6.350 1.125 7.220 1.295 ;
        RECT 6.350 2.190 7.220 2.360 ;
        RECT 7.050 1.125 7.220 2.630 ;
        RECT 7.050 1.525 7.275 1.825 ;
        RECT 7.050 2.460 8.655 2.630 ;
        RECT 8.485 2.460 8.655 2.980 ;
        RECT 8.485 2.810 11.855 2.980 ;
        RECT 7.455 1.060 7.625 2.280 ;
        RECT 7.455 1.325 8.190 1.495 ;
        RECT 7.455 2.110 9.005 2.280 ;
        RECT 8.835 1.655 9.005 2.630 ;
        RECT 11.540 1.310 11.710 2.630 ;
        RECT 11.540 1.310 11.940 1.480 ;
        RECT 8.835 2.460 12.395 2.630 ;
        RECT 12.225 2.460 12.395 2.835 ;
        RECT 2.460 0.750 2.630 1.825 ;
        RECT 6.845 0.700 7.040 0.930 ;
        RECT 2.460 0.750 7.040 0.930 ;
        RECT 6.845 0.700 7.985 0.880 ;
        RECT 7.805 0.700 7.985 1.090 ;
        RECT 8.625 0.595 8.795 1.090 ;
        RECT 7.805 0.910 8.795 1.090 ;
        RECT 8.625 0.595 9.655 0.775 ;
        RECT 9.950 0.765 11.550 0.945 ;
        RECT 11.810 0.575 12.370 0.760 ;
        RECT 12.430 0.575 12.445 0.820 ;
        RECT 12.520 0.650 12.750 0.820 ;
        RECT 12.580 0.650 12.750 1.480 ;
        RECT 12.580 1.310 13.705 1.480 ;
        RECT 13.375 0.875 13.545 1.480 ;
        RECT 13.535 1.310 13.705 2.215 ;
        RECT 13.280 2.045 13.705 2.215 ;
        RECT 12.445 0.585 12.455 0.819 ;
        RECT 12.455 0.595 12.465 0.819 ;
        RECT 12.465 0.605 12.475 0.819 ;
        RECT 12.475 0.615 12.485 0.819 ;
        RECT 12.485 0.625 12.495 0.819 ;
        RECT 12.495 0.635 12.505 0.819 ;
        RECT 12.505 0.645 12.515 0.819 ;
        RECT 12.515 0.650 12.521 0.820 ;
        RECT 12.370 0.575 12.380 0.759 ;
        RECT 12.380 0.575 12.390 0.769 ;
        RECT 12.390 0.575 12.400 0.779 ;
        RECT 12.400 0.575 12.410 0.789 ;
        RECT 12.410 0.575 12.420 0.799 ;
        RECT 12.420 0.575 12.430 0.809 ;
        RECT 11.740 0.575 11.750 0.819 ;
        RECT 11.750 0.575 11.760 0.809 ;
        RECT 11.760 0.575 11.770 0.799 ;
        RECT 11.770 0.575 11.780 0.789 ;
        RECT 11.780 0.575 11.790 0.779 ;
        RECT 11.790 0.575 11.800 0.769 ;
        RECT 11.800 0.575 11.810 0.759 ;
        RECT 11.625 0.690 11.635 0.934 ;
        RECT 11.635 0.680 11.645 0.924 ;
        RECT 11.645 0.670 11.655 0.914 ;
        RECT 11.655 0.660 11.665 0.904 ;
        RECT 11.665 0.650 11.675 0.894 ;
        RECT 11.675 0.640 11.685 0.884 ;
        RECT 11.685 0.630 11.695 0.874 ;
        RECT 11.695 0.620 11.705 0.864 ;
        RECT 11.705 0.610 11.715 0.854 ;
        RECT 11.715 0.600 11.725 0.844 ;
        RECT 11.725 0.590 11.735 0.834 ;
        RECT 11.735 0.580 11.741 0.830 ;
        RECT 11.550 0.765 11.560 0.945 ;
        RECT 11.560 0.755 11.570 0.945 ;
        RECT 11.570 0.745 11.580 0.945 ;
        RECT 11.580 0.735 11.590 0.945 ;
        RECT 11.590 0.725 11.600 0.945 ;
        RECT 11.600 0.715 11.610 0.945 ;
        RECT 11.610 0.705 11.620 0.945 ;
        RECT 11.620 0.695 11.626 0.945 ;
        RECT 9.825 0.650 9.835 0.944 ;
        RECT 9.835 0.660 9.845 0.944 ;
        RECT 9.845 0.670 9.855 0.944 ;
        RECT 9.855 0.680 9.865 0.944 ;
        RECT 9.865 0.690 9.875 0.944 ;
        RECT 9.875 0.700 9.885 0.944 ;
        RECT 9.885 0.710 9.895 0.944 ;
        RECT 9.895 0.720 9.905 0.944 ;
        RECT 9.905 0.730 9.915 0.944 ;
        RECT 9.915 0.740 9.925 0.944 ;
        RECT 9.925 0.750 9.935 0.944 ;
        RECT 9.935 0.760 9.945 0.944 ;
        RECT 9.945 0.765 9.951 0.945 ;
        RECT 9.780 0.605 9.790 0.899 ;
        RECT 9.790 0.615 9.800 0.909 ;
        RECT 9.800 0.625 9.810 0.919 ;
        RECT 9.810 0.635 9.820 0.929 ;
        RECT 9.820 0.640 9.826 0.940 ;
        RECT 9.655 0.595 9.665 0.775 ;
        RECT 9.665 0.595 9.675 0.785 ;
        RECT 9.675 0.595 9.685 0.795 ;
        RECT 9.685 0.595 9.695 0.805 ;
        RECT 9.695 0.595 9.705 0.815 ;
        RECT 9.705 0.595 9.715 0.825 ;
        RECT 9.715 0.595 9.725 0.835 ;
        RECT 9.725 0.595 9.735 0.845 ;
        RECT 9.735 0.595 9.745 0.855 ;
        RECT 9.745 0.595 9.755 0.865 ;
        RECT 9.755 0.595 9.765 0.875 ;
        RECT 9.765 0.595 9.775 0.885 ;
        RECT 9.775 0.595 9.781 0.895 ;
        RECT 11.890 0.940 12.190 1.110 ;
        RECT 12.090 1.040 12.290 1.120 ;
        RECT 12.100 1.040 12.290 1.130 ;
        RECT 12.110 1.040 12.290 1.140 ;
        RECT 11.890 2.045 12.190 2.215 ;
        RECT 11.890 0.950 12.200 1.110 ;
        RECT 11.890 0.960 12.210 1.110 ;
        RECT 11.890 0.970 12.220 1.110 ;
        RECT 11.890 0.980 12.230 1.110 ;
        RECT 11.890 0.990 12.240 1.110 ;
        RECT 11.890 1.000 12.250 1.110 ;
        RECT 11.890 1.010 12.260 1.110 ;
        RECT 11.890 1.020 12.270 1.110 ;
        RECT 11.890 1.030 12.280 1.110 ;
        RECT 12.120 1.040 12.290 2.214 ;
        RECT 12.930 1.675 13.100 2.565 ;
        RECT 12.120 1.675 13.355 1.845 ;
        RECT 14.070 1.540 14.240 2.565 ;
        RECT 12.930 2.395 14.240 2.565 ;
        RECT 14.070 1.540 14.260 1.840 ;
  END 
END FFSEDQHDLXHT

MACRO FFSEDQHD2XHT
  CLASS  CORE ;
  FOREIGN FFSEDQHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.990 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 15.130 0.720 15.300 2.960 ;
        RECT 15.130 2.030 15.485 2.425 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.835 1.475 1.130 2.020 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.625 0.580 2.010 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.805 1.545 3.180 2.020 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.675 -0.300 0.975 0.930 ;
        RECT 2.555 -0.300 2.855 0.570 ;
        RECT 3.540 -0.300 3.840 0.570 ;
        RECT 5.310 -0.300 5.610 0.570 ;
        RECT 6.940 -0.300 7.240 0.520 ;
        RECT 8.235 -0.300 8.405 0.730 ;
        RECT 10.270 -0.300 10.570 0.525 ;
        RECT 11.360 -0.300 11.660 0.565 ;
        RECT 13.550 -0.300 13.850 0.445 ;
        RECT 14.610 -0.300 14.780 1.120 ;
        RECT 15.650 -0.300 15.820 1.120 ;
        RECT 0.000 -0.300 15.990 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 6.385 1.525 6.870 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.705 1.465 6.050 2.010 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.685 2.640 0.985 3.990 ;
        RECT 2.555 2.910 2.855 3.990 ;
        RECT 3.420 2.910 3.720 3.990 ;
        RECT 5.310 2.890 5.610 3.990 ;
        RECT 6.940 3.160 7.240 3.990 ;
        RECT 8.205 2.810 8.375 3.990 ;
        RECT 10.280 3.160 10.580 3.990 ;
        RECT 11.265 3.160 11.565 3.990 ;
        RECT 13.480 2.765 13.780 3.990 ;
        RECT 14.545 2.975 14.845 3.990 ;
        RECT 15.650 2.570 15.820 3.990 ;
        RECT 0.000 3.390 15.990 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.110 1.500 1.280 ;
        RECT 1.330 1.110 1.500 2.375 ;
        RECT 0.105 2.205 1.500 2.375 ;
        RECT 1.330 1.705 1.600 2.005 ;
        RECT 1.680 0.945 1.950 1.245 ;
        RECT 1.780 0.945 1.950 2.875 ;
        RECT 1.680 2.235 1.950 2.875 ;
        RECT 3.710 1.775 3.880 2.730 ;
        RECT 1.680 2.550 3.880 2.730 ;
        RECT 3.360 1.110 3.530 2.370 ;
        RECT 3.030 2.200 3.530 2.370 ;
        RECT 3.030 1.110 4.190 1.280 ;
        RECT 4.020 1.110 4.190 1.650 ;
        RECT 4.065 1.480 4.235 3.060 ;
        RECT 4.020 1.480 4.420 1.650 ;
        RECT 4.065 2.890 4.920 3.060 ;
        RECT 5.165 1.110 5.335 2.360 ;
        RECT 5.165 1.110 6.180 1.280 ;
        RECT 5.165 2.190 6.180 2.360 ;
        RECT 4.415 1.890 4.585 2.710 ;
        RECT 4.370 1.110 4.770 1.280 ;
        RECT 4.600 1.110 4.770 2.070 ;
        RECT 4.415 1.890 4.770 2.070 ;
        RECT 4.415 2.540 6.440 2.710 ;
        RECT 6.270 2.540 6.440 2.980 ;
        RECT 6.270 2.810 8.005 2.980 ;
        RECT 7.835 2.810 8.005 3.110 ;
        RECT 9.275 0.955 9.445 2.280 ;
        RECT 9.210 0.955 9.510 1.125 ;
        RECT 9.275 1.675 10.880 1.845 ;
        RECT 10.850 1.125 11.150 1.495 ;
        RECT 10.040 1.325 11.755 1.495 ;
        RECT 11.585 1.325 11.755 2.215 ;
        RECT 10.830 2.045 11.755 2.215 ;
        RECT 7.495 1.060 7.665 2.215 ;
        RECT 7.495 1.325 8.260 1.495 ;
        RECT 7.495 2.045 9.075 2.215 ;
        RECT 8.905 1.655 9.075 2.630 ;
        RECT 8.905 2.460 12.815 2.630 ;
        RECT 12.645 2.460 12.815 2.795 ;
        RECT 6.390 1.125 7.250 1.295 ;
        RECT 6.390 2.190 7.250 2.360 ;
        RECT 7.080 1.125 7.250 2.630 ;
        RECT 7.080 1.525 7.315 1.825 ;
        RECT 7.080 2.460 8.725 2.630 ;
        RECT 8.555 2.460 8.725 2.980 ;
        RECT 8.555 2.810 12.360 2.980 ;
        RECT 12.190 2.810 12.360 3.210 ;
        RECT 12.730 1.350 13.175 1.520 ;
        RECT 12.995 1.350 13.175 3.210 ;
        RECT 12.190 3.040 13.175 3.210 ;
        RECT 2.360 0.750 2.530 1.825 ;
        RECT 6.885 0.700 7.285 0.930 ;
        RECT 2.360 0.750 7.285 0.930 ;
        RECT 6.885 0.700 8.055 0.880 ;
        RECT 7.875 0.700 8.055 1.090 ;
        RECT 8.730 0.595 8.900 1.090 ;
        RECT 7.875 0.910 8.900 1.090 ;
        RECT 9.780 0.595 9.950 0.945 ;
        RECT 8.730 0.595 9.950 0.775 ;
        RECT 9.780 0.765 11.790 0.945 ;
        RECT 12.050 0.575 12.800 0.760 ;
        RECT 13.050 0.480 13.350 0.820 ;
        RECT 12.860 0.575 13.350 0.820 ;
        RECT 12.860 0.650 14.430 0.820 ;
        RECT 14.035 1.125 14.430 1.295 ;
        RECT 14.260 0.650 14.430 2.225 ;
        RECT 14.035 2.055 14.430 2.225 ;
        RECT 12.800 0.575 12.810 0.759 ;
        RECT 12.810 0.575 12.820 0.769 ;
        RECT 12.820 0.575 12.830 0.779 ;
        RECT 12.830 0.575 12.840 0.789 ;
        RECT 12.840 0.575 12.850 0.799 ;
        RECT 12.850 0.575 12.860 0.809 ;
        RECT 11.980 0.575 11.990 0.819 ;
        RECT 11.990 0.575 12.000 0.809 ;
        RECT 12.000 0.575 12.010 0.799 ;
        RECT 12.010 0.575 12.020 0.789 ;
        RECT 12.020 0.575 12.030 0.779 ;
        RECT 12.030 0.575 12.040 0.769 ;
        RECT 12.040 0.575 12.050 0.759 ;
        RECT 11.865 0.690 11.875 0.934 ;
        RECT 11.875 0.680 11.885 0.924 ;
        RECT 11.885 0.670 11.895 0.914 ;
        RECT 11.895 0.660 11.905 0.904 ;
        RECT 11.905 0.650 11.915 0.894 ;
        RECT 11.915 0.640 11.925 0.884 ;
        RECT 11.925 0.630 11.935 0.874 ;
        RECT 11.935 0.620 11.945 0.864 ;
        RECT 11.945 0.610 11.955 0.854 ;
        RECT 11.955 0.600 11.965 0.844 ;
        RECT 11.965 0.590 11.975 0.834 ;
        RECT 11.975 0.580 11.981 0.830 ;
        RECT 11.790 0.765 11.800 0.945 ;
        RECT 11.800 0.755 11.810 0.945 ;
        RECT 11.810 0.745 11.820 0.945 ;
        RECT 11.820 0.735 11.830 0.945 ;
        RECT 11.830 0.725 11.840 0.945 ;
        RECT 11.840 0.715 11.850 0.945 ;
        RECT 11.850 0.705 11.860 0.945 ;
        RECT 11.860 0.695 11.866 0.945 ;
        RECT 12.065 1.000 12.245 2.240 ;
        RECT 12.065 2.070 12.590 2.240 ;
        RECT 12.065 1.000 13.820 1.170 ;
        RECT 13.650 1.000 13.820 2.585 ;
        RECT 13.650 1.595 13.995 1.765 ;
        RECT 14.780 1.540 14.950 2.585 ;
        RECT 13.650 2.415 14.950 2.585 ;
  END 
END FFSEDQHD2XHT

MACRO FFSEDQHD1XHT
  CLASS  CORE ;
  FOREIGN FFSEDQHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.760 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.420 0.720 14.660 1.360 ;
        RECT 14.450 0.720 14.660 2.960 ;
        RECT 14.420 1.980 14.660 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 1.325 1.220 1.880 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.540 0.620 2.010 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.840 1.465 3.245 1.950 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.775 -0.300 1.075 0.795 ;
        RECT 2.560 -0.300 2.880 0.570 ;
        RECT 3.640 -0.300 3.960 0.570 ;
        RECT 5.410 -0.300 5.710 0.570 ;
        RECT 6.810 -0.300 7.110 0.520 ;
        RECT 8.165 -0.300 8.335 0.730 ;
        RECT 9.970 -0.300 10.270 0.525 ;
        RECT 10.950 -0.300 11.250 0.565 ;
        RECT 12.840 -0.300 13.140 0.550 ;
        RECT 13.900 -0.300 14.070 1.120 ;
        RECT 0.000 -0.300 14.760 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 6.345 1.525 6.870 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.665 1.465 6.050 2.010 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.785 2.640 1.085 3.990 ;
        RECT 2.655 2.910 2.955 3.990 ;
        RECT 3.520 2.910 3.820 3.990 ;
        RECT 5.410 2.890 5.710 3.990 ;
        RECT 6.810 3.160 7.110 3.990 ;
        RECT 8.115 2.810 8.285 3.990 ;
        RECT 10.090 3.160 10.390 3.990 ;
        RECT 10.950 3.160 11.250 3.990 ;
        RECT 12.850 2.830 13.150 3.990 ;
        RECT 13.835 2.975 14.135 3.990 ;
        RECT 0.000 3.390 14.760 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.270 0.975 0.440 1.345 ;
        RECT 0.270 0.975 1.600 1.145 ;
        RECT 1.430 0.975 1.600 2.430 ;
        RECT 0.205 2.260 1.600 2.430 ;
        RECT 1.430 1.705 1.700 2.005 ;
        RECT 1.780 1.045 2.050 1.345 ;
        RECT 1.880 1.045 2.050 2.875 ;
        RECT 1.780 2.235 2.050 2.875 ;
        RECT 3.805 1.775 3.975 2.730 ;
        RECT 1.780 2.550 3.975 2.730 ;
        RECT 3.430 1.110 3.600 2.310 ;
        RECT 3.130 2.140 3.600 2.310 ;
        RECT 3.130 1.110 4.290 1.280 ;
        RECT 4.120 1.110 4.290 1.650 ;
        RECT 4.165 1.480 4.335 3.060 ;
        RECT 4.120 1.480 4.520 1.650 ;
        RECT 4.165 2.890 5.020 3.060 ;
        RECT 5.215 1.110 5.385 2.360 ;
        RECT 5.215 1.110 6.140 1.280 ;
        RECT 5.215 2.190 6.140 2.360 ;
        RECT 4.515 1.890 4.685 2.710 ;
        RECT 4.470 1.110 4.870 1.280 ;
        RECT 4.700 1.110 4.870 2.070 ;
        RECT 4.515 1.890 4.870 2.070 ;
        RECT 4.515 2.540 6.860 2.710 ;
        RECT 6.690 2.540 6.860 2.980 ;
        RECT 6.690 2.810 7.915 2.980 ;
        RECT 7.745 2.810 7.915 3.110 ;
        RECT 9.205 0.955 9.375 2.280 ;
        RECT 9.140 0.955 9.440 1.125 ;
        RECT 9.205 1.675 10.640 1.845 ;
        RECT 10.550 1.125 10.850 1.495 ;
        RECT 9.860 1.325 11.360 1.495 ;
        RECT 11.190 1.325 11.360 2.215 ;
        RECT 10.520 2.045 11.360 2.215 ;
        RECT 6.350 1.125 7.220 1.295 ;
        RECT 6.350 2.190 7.220 2.360 ;
        RECT 7.050 1.125 7.220 2.630 ;
        RECT 7.050 1.525 7.275 1.825 ;
        RECT 7.050 2.460 8.655 2.630 ;
        RECT 8.485 2.460 8.655 2.980 ;
        RECT 8.485 2.810 11.940 2.980 ;
        RECT 7.455 1.060 7.625 2.280 ;
        RECT 7.455 1.325 8.190 1.495 ;
        RECT 7.455 2.110 9.005 2.280 ;
        RECT 8.835 1.655 9.005 2.630 ;
        RECT 11.540 1.310 11.710 2.630 ;
        RECT 11.540 1.310 11.940 1.480 ;
        RECT 8.835 2.460 12.395 2.630 ;
        RECT 12.225 2.460 12.395 2.945 ;
        RECT 2.460 0.750 2.630 1.825 ;
        RECT 6.175 0.700 6.400 0.930 ;
        RECT 2.460 0.750 6.400 0.930 ;
        RECT 6.175 0.700 7.985 0.880 ;
        RECT 7.805 0.700 7.985 1.090 ;
        RECT 8.685 0.595 8.855 1.090 ;
        RECT 7.805 0.910 8.855 1.090 ;
        RECT 8.685 0.595 9.655 0.775 ;
        RECT 11.500 0.575 11.670 0.945 ;
        RECT 9.950 0.765 11.670 0.945 ;
        RECT 11.500 0.575 12.530 0.760 ;
        RECT 12.580 0.575 12.605 1.480 ;
        RECT 12.760 0.940 12.880 1.480 ;
        RECT 12.760 0.940 13.705 1.110 ;
        RECT 13.535 0.940 13.705 2.215 ;
        RECT 13.280 2.045 13.705 2.215 ;
        RECT 12.605 0.585 12.615 1.479 ;
        RECT 12.615 0.595 12.625 1.479 ;
        RECT 12.625 0.605 12.635 1.479 ;
        RECT 12.635 0.615 12.645 1.479 ;
        RECT 12.645 0.625 12.655 1.479 ;
        RECT 12.655 0.635 12.665 1.479 ;
        RECT 12.665 0.645 12.675 1.479 ;
        RECT 12.675 0.655 12.685 1.479 ;
        RECT 12.685 0.665 12.695 1.479 ;
        RECT 12.695 0.675 12.705 1.479 ;
        RECT 12.705 0.685 12.715 1.479 ;
        RECT 12.715 0.695 12.725 1.479 ;
        RECT 12.725 0.705 12.735 1.479 ;
        RECT 12.735 0.715 12.745 1.479 ;
        RECT 12.745 0.725 12.755 1.479 ;
        RECT 12.755 0.730 12.761 1.480 ;
        RECT 12.530 0.575 12.540 0.759 ;
        RECT 12.540 0.575 12.550 0.769 ;
        RECT 12.550 0.575 12.560 0.779 ;
        RECT 12.560 0.575 12.570 0.789 ;
        RECT 12.570 0.575 12.580 0.799 ;
        RECT 9.825 0.650 9.835 0.944 ;
        RECT 9.835 0.660 9.845 0.944 ;
        RECT 9.845 0.670 9.855 0.944 ;
        RECT 9.855 0.680 9.865 0.944 ;
        RECT 9.865 0.690 9.875 0.944 ;
        RECT 9.875 0.700 9.885 0.944 ;
        RECT 9.885 0.710 9.895 0.944 ;
        RECT 9.895 0.720 9.905 0.944 ;
        RECT 9.905 0.730 9.915 0.944 ;
        RECT 9.915 0.740 9.925 0.944 ;
        RECT 9.925 0.750 9.935 0.944 ;
        RECT 9.935 0.760 9.945 0.944 ;
        RECT 9.945 0.765 9.951 0.945 ;
        RECT 9.780 0.605 9.790 0.899 ;
        RECT 9.790 0.615 9.800 0.909 ;
        RECT 9.800 0.625 9.810 0.919 ;
        RECT 9.810 0.635 9.820 0.929 ;
        RECT 9.820 0.640 9.826 0.940 ;
        RECT 9.655 0.595 9.665 0.775 ;
        RECT 9.665 0.595 9.675 0.785 ;
        RECT 9.675 0.595 9.685 0.795 ;
        RECT 9.685 0.595 9.695 0.805 ;
        RECT 9.695 0.595 9.705 0.815 ;
        RECT 9.705 0.595 9.715 0.825 ;
        RECT 9.715 0.595 9.725 0.835 ;
        RECT 9.725 0.595 9.735 0.845 ;
        RECT 9.735 0.595 9.745 0.855 ;
        RECT 9.745 0.595 9.755 0.865 ;
        RECT 9.755 0.595 9.765 0.875 ;
        RECT 9.765 0.595 9.775 0.885 ;
        RECT 9.775 0.595 9.781 0.895 ;
        RECT 11.890 0.940 12.290 1.110 ;
        RECT 12.120 0.940 12.290 2.215 ;
        RECT 11.890 2.045 12.290 2.215 ;
        RECT 12.930 1.675 13.100 2.650 ;
        RECT 12.120 1.675 13.355 1.845 ;
        RECT 14.070 1.520 14.240 2.650 ;
        RECT 12.930 2.480 14.240 2.650 ;
        RECT 14.070 1.520 14.260 1.820 ;
  END 
END FFSEDQHD1XHT

MACRO FFSEDHQHD3XHT
  CLASS  CORE ;
  FOREIGN FFSEDHQHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.270 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 17.890 0.720 18.060 1.405 ;
        RECT 17.890 1.980 18.060 2.960 ;
        RECT 17.890 1.235 19.175 1.405 ;
        RECT 17.890 1.980 19.175 2.350 ;
        RECT 18.930 0.720 19.175 3.045 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.795 1.325 1.190 1.920 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.090 1.625 0.560 2.010 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.845 1.545 3.190 2.020 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.715 -0.300 1.015 0.775 ;
        RECT 2.500 -0.300 2.820 0.570 ;
        RECT 3.580 -0.300 3.900 0.570 ;
        RECT 5.350 -0.300 5.650 0.570 ;
        RECT 6.980 -0.300 7.280 0.520 ;
        RECT 7.970 -0.300 8.270 0.520 ;
        RECT 9.225 -0.300 9.525 0.580 ;
        RECT 11.435 -0.300 11.735 0.505 ;
        RECT 12.425 -0.300 12.725 0.585 ;
        RECT 14.280 -0.300 14.580 0.495 ;
        RECT 16.270 -0.300 16.445 0.660 ;
        RECT 17.365 -0.300 17.540 1.120 ;
        RECT 18.345 -0.300 18.645 1.055 ;
        RECT 0.000 -0.300 19.270 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 6.425 1.525 6.875 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.745 1.465 6.070 2.010 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.715 2.640 1.015 3.990 ;
        RECT 2.595 2.910 2.895 3.990 ;
        RECT 3.460 2.910 3.760 3.990 ;
        RECT 5.400 2.890 5.700 3.990 ;
        RECT 6.960 3.005 7.260 3.990 ;
        RECT 7.655 3.005 7.955 3.990 ;
        RECT 9.510 2.780 9.680 3.990 ;
        RECT 11.560 3.220 12.540 3.990 ;
        RECT 13.475 3.255 13.775 3.990 ;
        RECT 16.215 2.765 16.515 3.990 ;
        RECT 17.305 2.975 17.605 3.990 ;
        RECT 18.410 2.570 18.580 3.990 ;
        RECT 0.000 3.390 19.270 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.210 0.975 0.380 1.345 ;
        RECT 0.210 0.975 1.540 1.145 ;
        RECT 1.370 0.975 1.540 2.375 ;
        RECT 0.145 2.205 1.540 2.375 ;
        RECT 1.370 1.705 1.640 2.005 ;
        RECT 1.720 1.045 1.990 1.345 ;
        RECT 1.820 1.045 1.990 2.730 ;
        RECT 1.720 2.375 1.990 2.730 ;
        RECT 3.745 1.775 3.915 2.730 ;
        RECT 1.720 2.550 3.915 2.730 ;
        RECT 3.375 1.110 3.545 2.370 ;
        RECT 3.070 2.200 3.545 2.370 ;
        RECT 3.070 1.110 4.235 1.280 ;
        RECT 4.065 1.110 4.235 1.650 ;
        RECT 4.105 1.480 4.275 3.190 ;
        RECT 4.065 1.480 4.460 1.650 ;
        RECT 4.105 3.020 4.960 3.190 ;
        RECT 5.185 1.110 5.355 2.360 ;
        RECT 5.185 2.190 6.205 2.360 ;
        RECT 5.185 1.110 6.220 1.280 ;
        RECT 6.430 1.125 7.225 1.295 ;
        RECT 7.055 1.125 7.225 2.360 ;
        RECT 6.410 2.190 7.225 2.360 ;
        RECT 7.055 1.525 7.355 1.825 ;
        RECT 4.455 1.890 4.625 2.710 ;
        RECT 4.420 1.110 4.810 1.280 ;
        RECT 4.640 1.110 4.810 2.070 ;
        RECT 4.455 1.890 4.810 2.070 ;
        RECT 4.455 2.540 8.305 2.710 ;
        RECT 8.135 2.540 8.305 3.090 ;
        RECT 8.135 2.920 9.320 3.090 ;
        RECT 9.020 2.920 9.320 3.210 ;
        RECT 7.535 1.125 7.705 2.215 ;
        RECT 7.470 1.125 7.770 1.295 ;
        RECT 7.465 2.045 8.655 2.215 ;
        RECT 8.485 2.045 8.655 2.600 ;
        RECT 8.485 2.430 9.505 2.600 ;
        RECT 10.580 0.890 10.750 2.280 ;
        RECT 11.620 1.620 11.790 2.280 ;
        RECT 10.580 2.110 11.790 2.280 ;
        RECT 11.620 1.620 11.985 1.790 ;
        RECT 8.520 1.125 8.820 1.460 ;
        RECT 8.520 1.290 10.380 1.460 ;
        RECT 8.835 1.290 9.005 2.215 ;
        RECT 8.835 2.045 10.030 2.215 ;
        RECT 9.860 2.045 10.030 3.040 ;
        RECT 10.210 1.175 10.380 1.475 ;
        RECT 8.835 1.290 10.380 1.475 ;
        RECT 9.860 2.870 14.245 3.040 ;
        RECT 13.945 2.870 14.245 3.175 ;
        RECT 11.270 1.235 11.440 1.895 ;
        RECT 11.970 1.980 12.140 2.280 ;
        RECT 11.865 1.125 12.165 1.405 ;
        RECT 11.270 1.235 12.390 1.405 ;
        RECT 12.220 1.235 12.390 2.215 ;
        RECT 11.970 1.980 12.390 2.215 ;
        RECT 12.220 1.450 12.935 1.735 ;
        RECT 12.220 1.450 14.430 1.620 ;
        RECT 12.925 2.520 14.980 2.690 ;
        RECT 14.810 2.520 14.980 3.165 ;
        RECT 9.210 1.675 10.380 1.845 ;
        RECT 10.210 1.655 10.380 2.630 ;
        RECT 12.570 1.940 12.740 2.630 ;
        RECT 10.210 2.460 12.740 2.630 ;
        RECT 12.570 1.940 14.040 2.110 ;
        RECT 13.870 1.815 14.040 2.200 ;
        RECT 13.870 1.815 15.360 1.985 ;
        RECT 15.190 1.375 15.360 1.985 ;
        RECT 2.400 0.760 2.570 1.825 ;
        RECT 2.400 0.760 9.875 0.930 ;
        RECT 10.215 0.500 10.845 0.680 ;
        RECT 11.235 0.765 12.970 0.945 ;
        RECT 13.145 0.675 14.850 0.845 ;
        RECT 15.135 0.520 16.090 0.690 ;
        RECT 15.920 0.520 16.090 1.480 ;
        RECT 15.920 1.310 16.265 1.480 ;
        RECT 15.920 0.935 17.065 1.110 ;
        RECT 16.895 0.935 17.065 2.215 ;
        RECT 16.765 2.045 17.065 2.215 ;
        RECT 15.005 0.520 15.015 0.810 ;
        RECT 15.015 0.520 15.025 0.800 ;
        RECT 15.025 0.520 15.035 0.790 ;
        RECT 15.035 0.520 15.045 0.780 ;
        RECT 15.045 0.520 15.055 0.770 ;
        RECT 15.055 0.520 15.065 0.760 ;
        RECT 15.065 0.520 15.075 0.750 ;
        RECT 15.075 0.520 15.085 0.740 ;
        RECT 15.085 0.520 15.095 0.730 ;
        RECT 15.095 0.520 15.105 0.720 ;
        RECT 15.105 0.520 15.115 0.710 ;
        RECT 15.115 0.520 15.125 0.700 ;
        RECT 15.125 0.520 15.135 0.690 ;
        RECT 14.980 0.545 14.990 0.835 ;
        RECT 14.990 0.535 15.000 0.825 ;
        RECT 15.000 0.525 15.006 0.819 ;
        RECT 14.850 0.675 14.860 0.845 ;
        RECT 14.860 0.665 14.870 0.845 ;
        RECT 14.870 0.655 14.880 0.845 ;
        RECT 14.880 0.645 14.890 0.845 ;
        RECT 14.890 0.635 14.900 0.845 ;
        RECT 14.900 0.625 14.910 0.845 ;
        RECT 14.910 0.615 14.920 0.845 ;
        RECT 14.920 0.605 14.930 0.845 ;
        RECT 14.930 0.595 14.940 0.845 ;
        RECT 14.940 0.585 14.950 0.845 ;
        RECT 14.950 0.575 14.960 0.845 ;
        RECT 14.960 0.565 14.970 0.845 ;
        RECT 14.970 0.555 14.980 0.845 ;
        RECT 13.060 0.675 13.070 0.919 ;
        RECT 13.070 0.675 13.080 0.909 ;
        RECT 13.080 0.675 13.090 0.899 ;
        RECT 13.090 0.675 13.100 0.889 ;
        RECT 13.100 0.675 13.110 0.879 ;
        RECT 13.110 0.675 13.120 0.869 ;
        RECT 13.120 0.675 13.130 0.859 ;
        RECT 13.130 0.675 13.140 0.849 ;
        RECT 13.140 0.675 13.146 0.845 ;
        RECT 13.045 0.690 13.055 0.934 ;
        RECT 13.055 0.680 13.061 0.930 ;
        RECT 12.970 0.765 12.980 0.945 ;
        RECT 12.980 0.755 12.990 0.945 ;
        RECT 12.990 0.745 13.000 0.945 ;
        RECT 13.000 0.735 13.010 0.945 ;
        RECT 13.010 0.725 13.020 0.945 ;
        RECT 13.020 0.715 13.030 0.945 ;
        RECT 13.030 0.705 13.040 0.945 ;
        RECT 13.040 0.695 13.046 0.945 ;
        RECT 11.110 0.650 11.120 0.944 ;
        RECT 11.120 0.660 11.130 0.944 ;
        RECT 11.130 0.670 11.140 0.944 ;
        RECT 11.140 0.680 11.150 0.944 ;
        RECT 11.150 0.690 11.160 0.944 ;
        RECT 11.160 0.700 11.170 0.944 ;
        RECT 11.170 0.710 11.180 0.944 ;
        RECT 11.180 0.720 11.190 0.944 ;
        RECT 11.190 0.730 11.200 0.944 ;
        RECT 11.200 0.740 11.210 0.944 ;
        RECT 11.210 0.750 11.220 0.944 ;
        RECT 11.220 0.760 11.230 0.944 ;
        RECT 11.230 0.765 11.236 0.945 ;
        RECT 10.970 0.510 10.980 0.804 ;
        RECT 10.980 0.520 10.990 0.814 ;
        RECT 10.990 0.530 11.000 0.824 ;
        RECT 11.000 0.540 11.010 0.834 ;
        RECT 11.010 0.550 11.020 0.844 ;
        RECT 11.020 0.560 11.030 0.854 ;
        RECT 11.030 0.570 11.040 0.864 ;
        RECT 11.040 0.580 11.050 0.874 ;
        RECT 11.050 0.590 11.060 0.884 ;
        RECT 11.060 0.600 11.070 0.894 ;
        RECT 11.070 0.610 11.080 0.904 ;
        RECT 11.080 0.620 11.090 0.914 ;
        RECT 11.090 0.630 11.100 0.924 ;
        RECT 11.100 0.640 11.110 0.934 ;
        RECT 10.845 0.500 10.855 0.680 ;
        RECT 10.855 0.500 10.865 0.690 ;
        RECT 10.865 0.500 10.875 0.700 ;
        RECT 10.875 0.500 10.885 0.710 ;
        RECT 10.885 0.500 10.895 0.720 ;
        RECT 10.895 0.500 10.905 0.730 ;
        RECT 10.905 0.500 10.915 0.740 ;
        RECT 10.915 0.500 10.925 0.750 ;
        RECT 10.925 0.500 10.935 0.760 ;
        RECT 10.935 0.500 10.945 0.770 ;
        RECT 10.945 0.500 10.955 0.780 ;
        RECT 10.955 0.500 10.965 0.790 ;
        RECT 10.965 0.500 10.971 0.800 ;
        RECT 10.135 0.500 10.145 0.750 ;
        RECT 10.145 0.500 10.155 0.740 ;
        RECT 10.155 0.500 10.165 0.730 ;
        RECT 10.165 0.500 10.175 0.720 ;
        RECT 10.175 0.500 10.185 0.710 ;
        RECT 10.185 0.500 10.195 0.700 ;
        RECT 10.195 0.500 10.205 0.690 ;
        RECT 10.205 0.500 10.215 0.680 ;
        RECT 9.965 0.670 9.975 0.920 ;
        RECT 9.975 0.660 9.985 0.910 ;
        RECT 9.985 0.650 9.995 0.900 ;
        RECT 9.995 0.640 10.005 0.890 ;
        RECT 10.005 0.630 10.015 0.880 ;
        RECT 10.015 0.620 10.025 0.870 ;
        RECT 10.025 0.610 10.035 0.860 ;
        RECT 10.035 0.600 10.045 0.850 ;
        RECT 10.045 0.590 10.055 0.840 ;
        RECT 10.055 0.580 10.065 0.830 ;
        RECT 10.065 0.570 10.075 0.820 ;
        RECT 10.075 0.560 10.085 0.810 ;
        RECT 10.085 0.550 10.095 0.800 ;
        RECT 10.095 0.540 10.105 0.790 ;
        RECT 10.105 0.530 10.115 0.780 ;
        RECT 10.115 0.520 10.125 0.770 ;
        RECT 10.125 0.510 10.135 0.760 ;
        RECT 9.875 0.760 9.885 0.930 ;
        RECT 9.885 0.750 9.895 0.930 ;
        RECT 9.895 0.740 9.905 0.930 ;
        RECT 9.905 0.730 9.915 0.930 ;
        RECT 9.915 0.720 9.925 0.930 ;
        RECT 9.925 0.710 9.935 0.930 ;
        RECT 9.935 0.700 9.945 0.930 ;
        RECT 9.945 0.690 9.955 0.930 ;
        RECT 9.955 0.680 9.965 0.930 ;
        RECT 15.330 2.165 15.500 3.145 ;
        RECT 15.350 0.875 15.520 1.195 ;
        RECT 13.340 1.025 15.740 1.195 ;
        RECT 15.570 1.025 15.740 2.335 ;
        RECT 14.225 2.165 16.585 2.335 ;
        RECT 16.415 1.675 16.585 2.570 ;
        RECT 16.475 1.540 16.680 1.845 ;
        RECT 16.415 1.675 16.680 1.845 ;
        RECT 17.255 1.585 17.425 2.570 ;
        RECT 16.415 2.400 17.425 2.570 ;
        RECT 17.255 1.585 18.715 1.755 ;
  END 
END FFSEDHQHD3XHT

MACRO FFSEDHQHD2XHT
  CLASS  CORE ;
  FOREIGN FFSEDHQHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.040 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 17.180 0.720 17.440 2.960 ;
        RECT 17.180 1.610 17.530 2.045 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.795 1.325 1.190 1.920 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.090 1.625 0.560 2.010 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.845 1.545 3.190 2.020 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.715 -0.300 1.015 0.775 ;
        RECT 2.500 -0.300 2.820 0.570 ;
        RECT 3.580 -0.300 3.900 0.570 ;
        RECT 5.350 -0.300 5.670 0.570 ;
        RECT 6.980 -0.300 7.300 0.520 ;
        RECT 7.880 -0.300 8.200 0.520 ;
        RECT 9.310 -0.300 9.480 0.800 ;
        RECT 11.070 -0.300 11.370 0.550 ;
        RECT 12.145 -0.300 12.445 0.525 ;
        RECT 14.025 -0.300 14.325 0.480 ;
        RECT 15.720 -0.300 15.890 0.625 ;
        RECT 16.550 -0.300 16.850 0.620 ;
        RECT 17.700 -0.300 17.870 1.245 ;
        RECT 0.000 -0.300 18.040 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 6.425 1.525 6.875 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.745 1.465 6.070 2.010 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.715 2.640 1.015 3.990 ;
        RECT 2.595 2.910 2.895 3.990 ;
        RECT 3.460 2.910 3.760 3.990 ;
        RECT 5.400 2.890 5.700 3.990 ;
        RECT 7.080 2.890 7.720 3.990 ;
        RECT 9.280 2.525 9.450 3.990 ;
        RECT 11.330 3.180 12.310 3.990 ;
        RECT 13.195 3.185 13.495 3.990 ;
        RECT 15.635 2.760 15.935 3.990 ;
        RECT 16.595 2.975 16.895 3.990 ;
        RECT 17.700 2.230 17.870 3.990 ;
        RECT 0.000 3.390 18.040 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.210 0.975 0.380 1.345 ;
        RECT 0.210 0.975 1.540 1.145 ;
        RECT 1.370 0.975 1.540 2.375 ;
        RECT 0.145 2.205 1.540 2.375 ;
        RECT 1.370 1.705 1.640 2.005 ;
        RECT 1.720 1.045 1.990 1.345 ;
        RECT 1.820 1.045 1.990 2.730 ;
        RECT 1.720 2.370 1.990 2.730 ;
        RECT 3.745 1.775 3.915 2.730 ;
        RECT 1.720 2.550 3.915 2.730 ;
        RECT 3.370 1.110 3.540 2.370 ;
        RECT 3.070 2.200 3.540 2.370 ;
        RECT 3.070 1.110 4.230 1.280 ;
        RECT 4.060 1.110 4.230 1.650 ;
        RECT 4.105 1.480 4.275 3.190 ;
        RECT 4.060 1.480 4.460 1.650 ;
        RECT 4.105 3.020 4.960 3.190 ;
        RECT 5.185 1.110 5.355 2.360 ;
        RECT 5.185 1.110 6.220 1.280 ;
        RECT 5.185 2.190 6.220 2.360 ;
        RECT 6.430 1.125 7.225 1.295 ;
        RECT 7.055 1.125 7.225 2.360 ;
        RECT 6.430 2.190 7.225 2.360 ;
        RECT 7.055 1.525 7.355 1.825 ;
        RECT 7.535 1.125 7.705 2.215 ;
        RECT 7.470 1.125 7.770 1.295 ;
        RECT 7.470 2.045 8.455 2.215 ;
        RECT 8.285 2.045 8.455 2.630 ;
        RECT 8.285 2.460 8.940 2.630 ;
        RECT 4.455 1.890 4.625 2.710 ;
        RECT 4.410 1.110 4.810 1.280 ;
        RECT 4.640 1.110 4.810 2.070 ;
        RECT 4.455 1.890 4.810 2.070 ;
        RECT 4.455 2.540 8.085 2.710 ;
        RECT 7.915 2.540 8.085 3.080 ;
        RECT 7.915 2.910 9.080 3.080 ;
        RECT 8.910 2.910 9.080 3.210 ;
        RECT 10.350 0.955 10.520 2.280 ;
        RECT 10.285 0.955 10.585 1.125 ;
        RECT 10.350 1.675 11.785 1.845 ;
        RECT 11.005 1.315 12.145 1.485 ;
        RECT 11.695 1.105 11.995 1.485 ;
        RECT 11.975 1.305 12.145 2.215 ;
        RECT 11.665 2.045 12.145 2.215 ;
        RECT 11.975 1.440 12.690 1.610 ;
        RECT 12.710 2.350 12.880 2.650 ;
        RECT 12.710 2.480 14.455 2.650 ;
        RECT 8.505 1.125 8.805 1.295 ;
        RECT 8.635 1.125 8.805 2.260 ;
        RECT 8.635 2.090 9.800 2.260 ;
        RECT 9.630 2.090 9.800 3.000 ;
        RECT 13.975 2.830 14.190 3.160 ;
        RECT 9.630 2.830 14.190 3.000 ;
        RECT 13.975 2.990 14.615 3.160 ;
        RECT 9.030 1.565 10.150 1.735 ;
        RECT 9.980 1.565 10.150 2.630 ;
        RECT 12.335 1.790 12.505 2.630 ;
        RECT 9.980 2.460 12.505 2.630 ;
        RECT 13.370 1.410 13.540 1.960 ;
        RECT 12.335 1.790 13.540 1.960 ;
        RECT 13.370 1.470 14.830 1.640 ;
        RECT 14.660 1.375 14.830 1.675 ;
        RECT 2.400 0.750 2.570 1.825 ;
        RECT 2.400 0.750 8.920 0.920 ;
        RECT 9.720 0.605 9.890 1.190 ;
        RECT 9.270 1.020 9.890 1.190 ;
        RECT 9.720 0.605 10.730 0.775 ;
        RECT 10.995 0.735 12.650 0.915 ;
        RECT 12.795 0.660 14.450 0.845 ;
        RECT 14.670 0.525 15.540 0.695 ;
        RECT 15.370 0.525 15.540 1.110 ;
        RECT 15.490 0.935 15.660 1.545 ;
        RECT 15.370 0.935 16.555 1.110 ;
        RECT 16.385 0.935 16.555 2.215 ;
        RECT 16.175 2.045 16.555 2.215 ;
        RECT 14.585 0.525 14.595 0.769 ;
        RECT 14.595 0.525 14.605 0.759 ;
        RECT 14.605 0.525 14.615 0.749 ;
        RECT 14.615 0.525 14.625 0.739 ;
        RECT 14.625 0.525 14.635 0.729 ;
        RECT 14.635 0.525 14.645 0.719 ;
        RECT 14.645 0.525 14.655 0.709 ;
        RECT 14.655 0.525 14.665 0.699 ;
        RECT 14.665 0.525 14.671 0.695 ;
        RECT 14.520 0.590 14.530 0.834 ;
        RECT 14.530 0.580 14.540 0.824 ;
        RECT 14.540 0.570 14.550 0.814 ;
        RECT 14.550 0.560 14.560 0.804 ;
        RECT 14.560 0.550 14.570 0.794 ;
        RECT 14.570 0.540 14.580 0.784 ;
        RECT 14.580 0.530 14.586 0.780 ;
        RECT 14.450 0.660 14.460 0.844 ;
        RECT 14.460 0.650 14.470 0.844 ;
        RECT 14.470 0.640 14.480 0.844 ;
        RECT 14.480 0.630 14.490 0.844 ;
        RECT 14.490 0.620 14.500 0.844 ;
        RECT 14.500 0.610 14.510 0.844 ;
        RECT 14.510 0.600 14.520 0.844 ;
        RECT 12.725 0.660 12.735 0.904 ;
        RECT 12.735 0.660 12.745 0.894 ;
        RECT 12.745 0.660 12.755 0.884 ;
        RECT 12.755 0.660 12.765 0.874 ;
        RECT 12.765 0.660 12.775 0.864 ;
        RECT 12.775 0.660 12.785 0.854 ;
        RECT 12.785 0.660 12.795 0.844 ;
        RECT 12.650 0.735 12.660 0.915 ;
        RECT 12.660 0.725 12.670 0.915 ;
        RECT 12.670 0.715 12.680 0.915 ;
        RECT 12.680 0.705 12.690 0.915 ;
        RECT 12.690 0.695 12.700 0.915 ;
        RECT 12.700 0.685 12.710 0.915 ;
        RECT 12.710 0.675 12.720 0.915 ;
        RECT 12.720 0.665 12.726 0.915 ;
        RECT 10.870 0.620 10.880 0.914 ;
        RECT 10.880 0.630 10.890 0.914 ;
        RECT 10.890 0.640 10.900 0.914 ;
        RECT 10.900 0.650 10.910 0.914 ;
        RECT 10.910 0.660 10.920 0.914 ;
        RECT 10.920 0.670 10.930 0.914 ;
        RECT 10.930 0.680 10.940 0.914 ;
        RECT 10.940 0.690 10.950 0.914 ;
        RECT 10.950 0.700 10.960 0.914 ;
        RECT 10.960 0.710 10.970 0.914 ;
        RECT 10.970 0.720 10.980 0.914 ;
        RECT 10.980 0.730 10.990 0.914 ;
        RECT 10.990 0.735 10.996 0.915 ;
        RECT 10.865 0.610 10.871 0.910 ;
        RECT 10.730 0.605 10.740 0.775 ;
        RECT 10.740 0.605 10.750 0.785 ;
        RECT 10.750 0.605 10.760 0.795 ;
        RECT 10.760 0.605 10.770 0.805 ;
        RECT 10.770 0.605 10.780 0.815 ;
        RECT 10.780 0.605 10.790 0.825 ;
        RECT 10.790 0.605 10.800 0.835 ;
        RECT 10.800 0.605 10.810 0.845 ;
        RECT 10.810 0.605 10.820 0.855 ;
        RECT 10.820 0.605 10.830 0.865 ;
        RECT 10.830 0.605 10.840 0.875 ;
        RECT 10.840 0.605 10.850 0.885 ;
        RECT 10.850 0.605 10.860 0.895 ;
        RECT 10.860 0.605 10.866 0.905 ;
        RECT 9.190 0.950 9.200 1.190 ;
        RECT 9.200 0.960 9.210 1.190 ;
        RECT 9.210 0.970 9.220 1.190 ;
        RECT 9.220 0.980 9.230 1.190 ;
        RECT 9.230 0.990 9.240 1.190 ;
        RECT 9.240 1.000 9.250 1.190 ;
        RECT 9.250 1.010 9.260 1.190 ;
        RECT 9.260 1.020 9.270 1.190 ;
        RECT 9.000 0.760 9.010 1.000 ;
        RECT 9.010 0.770 9.020 1.010 ;
        RECT 9.020 0.780 9.030 1.020 ;
        RECT 9.030 0.790 9.040 1.030 ;
        RECT 9.040 0.800 9.050 1.040 ;
        RECT 9.050 0.810 9.060 1.050 ;
        RECT 9.060 0.820 9.070 1.060 ;
        RECT 9.070 0.830 9.080 1.070 ;
        RECT 9.080 0.840 9.090 1.080 ;
        RECT 9.090 0.850 9.100 1.090 ;
        RECT 9.100 0.860 9.110 1.100 ;
        RECT 9.110 0.870 9.120 1.110 ;
        RECT 9.120 0.880 9.130 1.120 ;
        RECT 9.130 0.890 9.140 1.130 ;
        RECT 9.140 0.900 9.150 1.140 ;
        RECT 9.150 0.910 9.160 1.150 ;
        RECT 9.160 0.920 9.170 1.160 ;
        RECT 9.170 0.930 9.180 1.170 ;
        RECT 9.180 0.940 9.190 1.180 ;
        RECT 8.920 0.750 8.930 0.920 ;
        RECT 8.930 0.750 8.940 0.930 ;
        RECT 8.940 0.750 8.950 0.940 ;
        RECT 8.950 0.750 8.960 0.950 ;
        RECT 8.960 0.750 8.970 0.960 ;
        RECT 8.970 0.750 8.980 0.970 ;
        RECT 8.980 0.750 8.990 0.980 ;
        RECT 8.990 0.750 9.000 0.990 ;
        RECT 14.800 0.875 14.970 1.195 ;
        RECT 13.100 1.025 15.190 1.195 ;
        RECT 15.020 1.025 15.190 2.300 ;
        RECT 13.635 2.130 15.995 2.300 ;
        RECT 15.825 1.675 15.995 2.570 ;
        RECT 15.980 1.540 16.185 1.845 ;
        RECT 15.825 1.675 16.185 1.845 ;
        RECT 16.830 1.520 17.000 2.570 ;
        RECT 15.825 2.400 17.000 2.570 ;
  END 
END FFSEDHQHD2XHT

MACRO FFSEDHQHD1XHT
  CLASS  CORE ;
  FOREIGN FFSEDHQHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.990 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 15.650 0.720 15.895 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 1.325 1.220 1.920 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.625 0.620 2.010 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.905 1.495 3.205 2.020 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.775 -0.300 1.075 0.775 ;
        RECT 2.560 -0.300 2.880 0.570 ;
        RECT 3.640 -0.300 3.960 0.570 ;
        RECT 5.410 -0.300 5.710 0.570 ;
        RECT 7.040 -0.300 7.360 0.520 ;
        RECT 7.960 -0.300 8.280 0.520 ;
        RECT 9.370 -0.300 9.540 0.850 ;
        RECT 11.175 -0.300 11.475 0.525 ;
        RECT 12.205 -0.300 12.505 0.565 ;
        RECT 14.095 -0.300 14.395 0.695 ;
        RECT 15.020 -0.300 15.320 0.620 ;
        RECT 0.000 -0.300 15.990 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 6.485 1.525 6.935 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.805 1.465 6.130 2.010 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.775 2.640 1.085 3.990 ;
        RECT 2.655 2.910 2.955 3.990 ;
        RECT 3.520 2.910 3.820 3.990 ;
        RECT 5.460 2.890 5.760 3.990 ;
        RECT 7.070 2.890 7.370 3.990 ;
        RECT 7.705 2.890 8.005 3.990 ;
        RECT 9.340 2.535 9.510 3.990 ;
        RECT 11.390 3.160 12.370 3.990 ;
        RECT 14.105 2.830 14.405 3.990 ;
        RECT 15.065 2.975 15.365 3.990 ;
        RECT 0.000 3.390 15.990 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.270 0.975 0.440 1.345 ;
        RECT 0.270 0.975 1.600 1.145 ;
        RECT 1.430 0.975 1.600 2.375 ;
        RECT 0.205 2.205 1.600 2.375 ;
        RECT 1.430 1.705 1.700 2.005 ;
        RECT 1.780 1.045 2.050 1.345 ;
        RECT 1.880 1.045 2.050 2.730 ;
        RECT 1.780 2.370 2.050 2.730 ;
        RECT 3.805 1.775 3.975 2.730 ;
        RECT 1.780 2.550 3.975 2.730 ;
        RECT 3.430 1.110 3.600 2.370 ;
        RECT 3.130 2.200 3.600 2.370 ;
        RECT 3.130 1.110 4.290 1.280 ;
        RECT 4.120 1.110 4.290 1.650 ;
        RECT 4.165 1.480 4.335 3.190 ;
        RECT 4.120 1.480 4.520 1.650 ;
        RECT 4.165 3.020 5.020 3.190 ;
        RECT 5.245 1.110 5.415 2.360 ;
        RECT 5.245 1.110 6.280 1.280 ;
        RECT 5.245 2.190 6.280 2.360 ;
        RECT 6.490 1.125 7.285 1.295 ;
        RECT 7.115 1.125 7.285 2.360 ;
        RECT 6.490 2.190 7.285 2.360 ;
        RECT 7.115 1.525 7.415 1.825 ;
        RECT 7.635 1.125 7.805 2.280 ;
        RECT 7.530 1.125 7.830 1.295 ;
        RECT 7.635 2.095 8.705 2.280 ;
        RECT 8.535 2.095 8.705 2.630 ;
        RECT 8.535 2.460 9.000 2.630 ;
        RECT 4.515 1.890 4.685 2.710 ;
        RECT 4.470 1.110 4.870 1.280 ;
        RECT 4.700 1.110 4.870 2.070 ;
        RECT 4.515 1.890 4.870 2.070 ;
        RECT 4.515 2.540 8.355 2.710 ;
        RECT 8.185 2.540 8.355 3.075 ;
        RECT 8.185 2.905 9.140 3.075 ;
        RECT 8.970 2.905 9.140 3.205 ;
        RECT 10.410 0.955 10.580 2.280 ;
        RECT 10.345 0.955 10.645 1.125 ;
        RECT 10.410 1.675 11.845 1.845 ;
        RECT 11.755 1.125 12.055 1.495 ;
        RECT 11.065 1.325 12.615 1.495 ;
        RECT 12.445 1.325 12.615 2.215 ;
        RECT 11.725 2.045 12.615 2.215 ;
        RECT 8.565 1.125 8.865 1.295 ;
        RECT 8.695 1.125 8.865 1.560 ;
        RECT 8.695 1.390 9.055 1.560 ;
        RECT 8.885 1.390 9.055 2.260 ;
        RECT 8.885 2.090 9.860 2.260 ;
        RECT 9.690 2.090 9.860 2.980 ;
        RECT 9.690 2.810 13.195 2.980 ;
        RECT 12.895 2.810 13.195 3.195 ;
        RECT 9.240 1.390 9.410 1.690 ;
        RECT 9.240 1.520 10.210 1.690 ;
        RECT 10.040 1.520 10.210 2.630 ;
        RECT 12.795 1.310 12.965 2.630 ;
        RECT 12.795 1.310 13.195 1.480 ;
        RECT 10.040 2.460 13.650 2.630 ;
        RECT 13.480 2.460 13.650 2.945 ;
        RECT 2.460 0.750 2.630 1.825 ;
        RECT 2.460 0.750 8.925 0.920 ;
        RECT 9.295 1.040 9.750 1.210 ;
        RECT 10.040 0.605 10.860 0.775 ;
        RECT 11.155 0.765 12.805 0.945 ;
        RECT 13.065 0.575 13.630 0.760 ;
        RECT 14.005 0.935 14.135 1.480 ;
        RECT 14.005 0.935 15.025 1.110 ;
        RECT 14.855 0.935 15.025 2.215 ;
        RECT 14.645 2.045 15.025 2.215 ;
        RECT 13.835 0.715 13.845 1.479 ;
        RECT 13.845 0.725 13.855 1.479 ;
        RECT 13.855 0.735 13.865 1.479 ;
        RECT 13.865 0.745 13.875 1.479 ;
        RECT 13.875 0.755 13.885 1.479 ;
        RECT 13.885 0.765 13.895 1.479 ;
        RECT 13.895 0.775 13.905 1.479 ;
        RECT 13.905 0.785 13.915 1.479 ;
        RECT 13.915 0.795 13.925 1.479 ;
        RECT 13.925 0.805 13.935 1.479 ;
        RECT 13.935 0.815 13.945 1.479 ;
        RECT 13.945 0.825 13.955 1.479 ;
        RECT 13.955 0.835 13.965 1.479 ;
        RECT 13.965 0.845 13.975 1.479 ;
        RECT 13.975 0.855 13.985 1.479 ;
        RECT 13.985 0.865 13.995 1.479 ;
        RECT 13.995 0.875 14.005 1.479 ;
        RECT 13.705 0.585 13.715 0.835 ;
        RECT 13.715 0.595 13.725 0.845 ;
        RECT 13.725 0.605 13.735 0.855 ;
        RECT 13.735 0.615 13.745 0.865 ;
        RECT 13.745 0.625 13.755 0.875 ;
        RECT 13.755 0.635 13.765 0.885 ;
        RECT 13.765 0.645 13.775 0.895 ;
        RECT 13.775 0.655 13.785 0.905 ;
        RECT 13.785 0.665 13.795 0.915 ;
        RECT 13.795 0.675 13.805 0.925 ;
        RECT 13.805 0.685 13.815 0.935 ;
        RECT 13.815 0.695 13.825 0.945 ;
        RECT 13.825 0.705 13.835 0.955 ;
        RECT 13.630 0.575 13.640 0.759 ;
        RECT 13.640 0.575 13.650 0.769 ;
        RECT 13.650 0.575 13.660 0.779 ;
        RECT 13.660 0.575 13.670 0.789 ;
        RECT 13.670 0.575 13.680 0.799 ;
        RECT 13.680 0.575 13.690 0.809 ;
        RECT 13.690 0.575 13.700 0.819 ;
        RECT 13.700 0.575 13.706 0.829 ;
        RECT 12.995 0.575 13.005 0.819 ;
        RECT 13.005 0.575 13.015 0.809 ;
        RECT 13.015 0.575 13.025 0.799 ;
        RECT 13.025 0.575 13.035 0.789 ;
        RECT 13.035 0.575 13.045 0.779 ;
        RECT 13.045 0.575 13.055 0.769 ;
        RECT 13.055 0.575 13.065 0.759 ;
        RECT 12.880 0.690 12.890 0.934 ;
        RECT 12.890 0.680 12.900 0.924 ;
        RECT 12.900 0.670 12.910 0.914 ;
        RECT 12.910 0.660 12.920 0.904 ;
        RECT 12.920 0.650 12.930 0.894 ;
        RECT 12.930 0.640 12.940 0.884 ;
        RECT 12.940 0.630 12.950 0.874 ;
        RECT 12.950 0.620 12.960 0.864 ;
        RECT 12.960 0.610 12.970 0.854 ;
        RECT 12.970 0.600 12.980 0.844 ;
        RECT 12.980 0.590 12.990 0.834 ;
        RECT 12.990 0.580 12.996 0.830 ;
        RECT 12.805 0.765 12.815 0.945 ;
        RECT 12.815 0.755 12.825 0.945 ;
        RECT 12.825 0.745 12.835 0.945 ;
        RECT 12.835 0.735 12.845 0.945 ;
        RECT 12.845 0.725 12.855 0.945 ;
        RECT 12.855 0.715 12.865 0.945 ;
        RECT 12.865 0.705 12.875 0.945 ;
        RECT 12.875 0.695 12.881 0.945 ;
        RECT 11.030 0.650 11.040 0.944 ;
        RECT 11.040 0.660 11.050 0.944 ;
        RECT 11.050 0.670 11.060 0.944 ;
        RECT 11.060 0.680 11.070 0.944 ;
        RECT 11.070 0.690 11.080 0.944 ;
        RECT 11.080 0.700 11.090 0.944 ;
        RECT 11.090 0.710 11.100 0.944 ;
        RECT 11.100 0.720 11.110 0.944 ;
        RECT 11.110 0.730 11.120 0.944 ;
        RECT 11.120 0.740 11.130 0.944 ;
        RECT 11.130 0.750 11.140 0.944 ;
        RECT 11.140 0.760 11.150 0.944 ;
        RECT 11.150 0.765 11.156 0.945 ;
        RECT 10.995 0.615 11.005 0.909 ;
        RECT 11.005 0.625 11.015 0.919 ;
        RECT 11.015 0.635 11.025 0.929 ;
        RECT 11.025 0.640 11.031 0.940 ;
        RECT 10.860 0.605 10.870 0.775 ;
        RECT 10.870 0.605 10.880 0.785 ;
        RECT 10.880 0.605 10.890 0.795 ;
        RECT 10.890 0.605 10.900 0.805 ;
        RECT 10.900 0.605 10.910 0.815 ;
        RECT 10.910 0.605 10.920 0.825 ;
        RECT 10.920 0.605 10.930 0.835 ;
        RECT 10.930 0.605 10.940 0.845 ;
        RECT 10.940 0.605 10.950 0.855 ;
        RECT 10.950 0.605 10.960 0.865 ;
        RECT 10.960 0.605 10.970 0.875 ;
        RECT 10.970 0.605 10.980 0.885 ;
        RECT 10.980 0.605 10.990 0.895 ;
        RECT 10.990 0.605 10.996 0.905 ;
        RECT 9.870 0.605 9.880 1.169 ;
        RECT 9.880 0.605 9.890 1.159 ;
        RECT 9.890 0.605 9.900 1.149 ;
        RECT 9.900 0.605 9.910 1.139 ;
        RECT 9.910 0.605 9.920 1.129 ;
        RECT 9.920 0.605 9.930 1.119 ;
        RECT 9.930 0.605 9.940 1.109 ;
        RECT 9.940 0.605 9.950 1.099 ;
        RECT 9.950 0.605 9.960 1.089 ;
        RECT 9.960 0.605 9.970 1.079 ;
        RECT 9.970 0.605 9.980 1.069 ;
        RECT 9.980 0.605 9.990 1.059 ;
        RECT 9.990 0.605 10.000 1.049 ;
        RECT 10.000 0.605 10.010 1.039 ;
        RECT 10.010 0.605 10.020 1.029 ;
        RECT 10.020 0.605 10.030 1.019 ;
        RECT 10.030 0.605 10.040 1.009 ;
        RECT 9.840 0.950 9.850 1.200 ;
        RECT 9.850 0.940 9.860 1.190 ;
        RECT 9.860 0.930 9.870 1.180 ;
        RECT 9.750 1.040 9.760 1.210 ;
        RECT 9.760 1.030 9.770 1.210 ;
        RECT 9.770 1.020 9.780 1.210 ;
        RECT 9.780 1.010 9.790 1.210 ;
        RECT 9.790 1.000 9.800 1.210 ;
        RECT 9.800 0.990 9.810 1.210 ;
        RECT 9.810 0.980 9.820 1.210 ;
        RECT 9.820 0.970 9.830 1.210 ;
        RECT 9.830 0.960 9.840 1.210 ;
        RECT 9.215 0.970 9.225 1.210 ;
        RECT 9.225 0.980 9.235 1.210 ;
        RECT 9.235 0.990 9.245 1.210 ;
        RECT 9.245 1.000 9.255 1.210 ;
        RECT 9.255 1.010 9.265 1.210 ;
        RECT 9.265 1.020 9.275 1.210 ;
        RECT 9.275 1.030 9.285 1.210 ;
        RECT 9.285 1.040 9.295 1.210 ;
        RECT 9.005 0.760 9.015 1.000 ;
        RECT 9.015 0.770 9.025 1.010 ;
        RECT 9.025 0.780 9.035 1.020 ;
        RECT 9.035 0.790 9.045 1.030 ;
        RECT 9.045 0.800 9.055 1.040 ;
        RECT 9.055 0.810 9.065 1.050 ;
        RECT 9.065 0.820 9.075 1.060 ;
        RECT 9.075 0.830 9.085 1.070 ;
        RECT 9.085 0.840 9.095 1.080 ;
        RECT 9.095 0.850 9.105 1.090 ;
        RECT 9.105 0.860 9.115 1.100 ;
        RECT 9.115 0.870 9.125 1.110 ;
        RECT 9.125 0.880 9.135 1.120 ;
        RECT 9.135 0.890 9.145 1.130 ;
        RECT 9.145 0.900 9.155 1.140 ;
        RECT 9.155 0.910 9.165 1.150 ;
        RECT 9.165 0.920 9.175 1.160 ;
        RECT 9.175 0.930 9.185 1.170 ;
        RECT 9.185 0.940 9.195 1.180 ;
        RECT 9.195 0.950 9.205 1.190 ;
        RECT 9.205 0.960 9.215 1.200 ;
        RECT 8.925 0.750 8.935 0.920 ;
        RECT 8.935 0.750 8.945 0.930 ;
        RECT 8.945 0.750 8.955 0.940 ;
        RECT 8.955 0.750 8.965 0.950 ;
        RECT 8.965 0.750 8.975 0.960 ;
        RECT 8.975 0.750 8.985 0.970 ;
        RECT 8.985 0.750 8.995 0.980 ;
        RECT 8.995 0.750 9.005 0.990 ;
        RECT 13.145 0.940 13.545 1.110 ;
        RECT 13.375 0.940 13.545 2.215 ;
        RECT 13.145 2.045 13.545 2.215 ;
        RECT 14.295 1.675 14.465 2.650 ;
        RECT 14.485 1.540 14.655 1.845 ;
        RECT 13.375 1.675 14.655 1.845 ;
        RECT 15.300 1.520 15.470 2.650 ;
        RECT 14.295 2.480 15.470 2.650 ;
  END 
END FFSEDHQHD1XHT

MACRO FFSEDHDMXHT
  CLASS  CORE ;
  FOREIGN FFSEDHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.170 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.825 1.060 15.070 1.360 ;
        RECT 14.860 1.060 15.070 2.280 ;
        RECT 14.825 1.980 15.070 2.280 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.845 1.060 14.250 1.360 ;
        RECT 14.040 1.060 14.250 2.300 ;
        RECT 13.845 2.000 14.250 2.300 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.325 1.120 1.540 ;
        RECT 0.950 1.325 1.120 1.960 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.680 0.315 2.010 ;
        RECT 0.100 1.720 0.585 2.010 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.650 1.830 2.850 2.360 ;
        RECT 2.455 2.150 2.850 2.360 ;
        RECT 2.870 1.575 3.040 2.020 ;
        RECT 2.650 1.830 3.040 2.020 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.775 ;
        RECT 2.435 -0.300 2.735 0.570 ;
        RECT 3.495 -0.300 3.795 0.570 ;
        RECT 5.250 -0.300 5.550 0.570 ;
        RECT 6.770 -0.300 7.070 0.520 ;
        RECT 8.125 -0.300 8.295 0.730 ;
        RECT 10.050 -0.300 10.350 0.525 ;
        RECT 10.900 -0.300 11.200 0.565 ;
        RECT 12.800 -0.300 13.100 0.560 ;
        RECT 14.210 -0.300 14.510 0.595 ;
        RECT 0.000 -0.300 15.170 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 6.250 1.525 6.755 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.530 1.465 6.050 2.010 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 2.575 0.890 3.990 ;
        RECT 2.555 2.910 2.855 3.990 ;
        RECT 3.420 2.910 3.720 3.990 ;
        RECT 5.310 2.890 5.610 3.990 ;
        RECT 6.890 3.095 7.190 3.990 ;
        RECT 8.095 2.745 8.265 3.990 ;
        RECT 10.050 3.160 10.350 3.990 ;
        RECT 10.910 3.160 11.210 3.990 ;
        RECT 12.810 2.830 13.110 3.990 ;
        RECT 14.210 2.925 14.510 3.990 ;
        RECT 0.000 3.390 15.170 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.490 1.145 ;
        RECT 1.320 0.975 1.490 2.375 ;
        RECT 1.320 1.770 1.500 2.375 ;
        RECT 0.105 2.205 1.500 2.375 ;
        RECT 1.320 1.770 1.665 1.940 ;
        RECT 1.670 1.045 2.015 1.345 ;
        RECT 1.845 1.045 2.015 2.730 ;
        RECT 1.680 2.120 2.015 2.730 ;
        RECT 3.705 1.775 3.875 2.730 ;
        RECT 1.680 2.550 3.875 2.730 ;
        RECT 3.330 1.110 3.500 2.370 ;
        RECT 3.030 2.200 3.500 2.370 ;
        RECT 2.985 1.110 4.190 1.280 ;
        RECT 4.020 1.110 4.190 1.650 ;
        RECT 4.065 1.480 4.235 3.115 ;
        RECT 4.020 1.480 4.420 1.650 ;
        RECT 4.065 2.945 4.870 3.115 ;
        RECT 5.145 1.110 5.315 2.360 ;
        RECT 5.145 1.110 6.100 1.280 ;
        RECT 5.145 2.190 6.100 2.360 ;
        RECT 4.370 1.110 4.770 1.280 ;
        RECT 4.600 1.110 4.770 2.710 ;
        RECT 4.415 2.390 4.770 2.710 ;
        RECT 4.415 2.540 6.820 2.710 ;
        RECT 6.650 2.540 6.820 2.915 ;
        RECT 6.650 2.745 7.895 2.915 ;
        RECT 7.725 2.745 7.895 3.045 ;
        RECT 9.165 0.955 9.335 2.280 ;
        RECT 9.100 0.955 9.400 1.125 ;
        RECT 9.165 1.675 10.600 1.845 ;
        RECT 10.510 1.125 10.810 1.495 ;
        RECT 9.820 1.325 11.320 1.495 ;
        RECT 11.150 1.325 11.320 2.215 ;
        RECT 10.480 2.045 11.320 2.215 ;
        RECT 6.310 1.125 7.170 1.295 ;
        RECT 6.310 2.190 7.170 2.360 ;
        RECT 7.000 1.125 7.170 2.565 ;
        RECT 7.000 1.525 7.235 1.825 ;
        RECT 7.000 2.395 8.615 2.565 ;
        RECT 8.445 2.395 8.615 2.980 ;
        RECT 8.445 2.810 11.900 2.980 ;
        RECT 7.415 1.060 7.585 2.215 ;
        RECT 7.415 1.325 8.150 1.495 ;
        RECT 7.415 2.045 8.965 2.215 ;
        RECT 8.795 1.655 8.965 2.630 ;
        RECT 11.500 1.310 11.670 2.630 ;
        RECT 11.500 1.310 11.900 1.480 ;
        RECT 8.795 2.460 12.355 2.630 ;
        RECT 12.185 2.460 12.355 2.945 ;
        RECT 2.425 0.750 2.595 1.650 ;
        RECT 2.295 1.480 2.595 1.650 ;
        RECT 6.220 0.700 6.405 0.930 ;
        RECT 2.425 0.750 6.405 0.930 ;
        RECT 6.220 0.700 7.945 0.880 ;
        RECT 7.765 0.700 7.945 1.090 ;
        RECT 8.630 0.595 8.800 1.090 ;
        RECT 7.765 0.910 8.800 1.090 ;
        RECT 9.660 0.595 9.830 0.945 ;
        RECT 8.630 0.595 9.830 0.775 ;
        RECT 11.445 0.575 11.615 0.945 ;
        RECT 9.660 0.765 11.615 0.945 ;
        RECT 11.445 0.575 12.430 0.760 ;
        RECT 12.720 0.940 12.840 1.480 ;
        RECT 12.720 0.940 13.665 1.110 ;
        RECT 13.495 0.940 13.665 2.215 ;
        RECT 13.240 2.045 13.665 2.215 ;
        RECT 13.495 1.650 13.860 1.820 ;
        RECT 12.540 0.620 12.550 1.480 ;
        RECT 12.550 0.630 12.560 1.480 ;
        RECT 12.560 0.640 12.570 1.480 ;
        RECT 12.570 0.650 12.580 1.480 ;
        RECT 12.580 0.660 12.590 1.480 ;
        RECT 12.590 0.670 12.600 1.480 ;
        RECT 12.600 0.680 12.610 1.480 ;
        RECT 12.610 0.690 12.620 1.480 ;
        RECT 12.620 0.700 12.630 1.480 ;
        RECT 12.630 0.710 12.640 1.480 ;
        RECT 12.640 0.720 12.650 1.480 ;
        RECT 12.650 0.730 12.660 1.480 ;
        RECT 12.660 0.740 12.670 1.480 ;
        RECT 12.670 0.750 12.680 1.480 ;
        RECT 12.680 0.760 12.690 1.480 ;
        RECT 12.690 0.770 12.700 1.480 ;
        RECT 12.700 0.780 12.710 1.480 ;
        RECT 12.710 0.790 12.720 1.480 ;
        RECT 12.505 0.585 12.515 0.835 ;
        RECT 12.515 0.595 12.525 0.845 ;
        RECT 12.525 0.605 12.535 0.855 ;
        RECT 12.535 0.610 12.541 0.864 ;
        RECT 12.430 0.575 12.440 0.759 ;
        RECT 12.440 0.575 12.450 0.769 ;
        RECT 12.450 0.575 12.460 0.779 ;
        RECT 12.460 0.575 12.470 0.789 ;
        RECT 12.470 0.575 12.480 0.799 ;
        RECT 12.480 0.575 12.490 0.809 ;
        RECT 12.490 0.575 12.500 0.819 ;
        RECT 12.500 0.575 12.506 0.829 ;
        RECT 11.850 0.940 12.250 1.110 ;
        RECT 12.080 0.940 12.250 2.215 ;
        RECT 11.850 2.045 12.250 2.215 ;
        RECT 12.890 1.675 13.060 2.650 ;
        RECT 12.080 1.675 13.315 1.845 ;
        RECT 14.475 1.520 14.645 2.650 ;
        RECT 12.890 2.480 14.645 2.650 ;
        RECT 14.475 1.520 14.675 1.820 ;
  END 
END FFSEDHDMXHT

MACRO FFSEDHDLXHT
  CLASS  CORE ;
  FOREIGN FFSEDHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.170 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.825 1.060 15.070 1.360 ;
        RECT 14.860 1.060 15.070 2.470 ;
        RECT 14.825 1.980 15.070 2.470 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.785 1.060 14.250 1.360 ;
        RECT 14.040 1.060 14.250 2.300 ;
        RECT 13.785 2.000 14.250 2.300 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.325 1.000 1.540 ;
        RECT 0.830 1.325 1.000 2.005 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.680 0.315 2.010 ;
        RECT 0.100 1.720 0.585 2.010 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.530 1.830 2.730 2.360 ;
        RECT 2.070 2.150 2.730 2.360 ;
        RECT 2.750 1.575 2.920 2.020 ;
        RECT 2.530 1.830 2.920 2.020 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.775 ;
        RECT 2.360 -0.300 2.660 0.570 ;
        RECT 3.420 -0.300 3.720 0.570 ;
        RECT 5.170 -0.300 5.470 0.570 ;
        RECT 6.710 -0.300 7.010 0.520 ;
        RECT 8.065 -0.300 8.235 0.730 ;
        RECT 9.870 -0.300 10.170 0.525 ;
        RECT 10.840 -0.300 11.140 0.565 ;
        RECT 12.740 -0.300 13.040 0.560 ;
        RECT 14.210 -0.300 14.510 0.745 ;
        RECT 0.000 -0.300 15.170 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 6.250 1.525 6.695 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.430 1.465 5.800 2.010 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.830 0.955 3.990 ;
        RECT 2.435 2.910 2.735 3.990 ;
        RECT 3.300 2.910 3.600 3.990 ;
        RECT 5.190 2.890 5.490 3.990 ;
        RECT 6.830 3.095 7.130 3.990 ;
        RECT 8.015 2.810 8.185 3.990 ;
        RECT 9.990 3.160 10.290 3.990 ;
        RECT 10.850 3.160 11.150 3.990 ;
        RECT 12.750 2.830 13.050 3.990 ;
        RECT 14.210 2.830 14.510 3.990 ;
        RECT 0.000 3.390 15.170 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.370 1.145 ;
        RECT 1.200 0.975 1.370 2.430 ;
        RECT 1.200 1.705 1.380 2.430 ;
        RECT 0.105 2.260 1.380 2.430 ;
        RECT 1.200 1.705 1.480 2.005 ;
        RECT 1.550 0.945 1.830 1.245 ;
        RECT 1.660 0.945 1.830 2.730 ;
        RECT 1.560 2.215 1.830 2.730 ;
        RECT 3.585 1.775 3.755 2.730 ;
        RECT 1.560 2.550 3.755 2.730 ;
        RECT 3.210 1.110 3.380 2.370 ;
        RECT 2.910 2.200 3.380 2.370 ;
        RECT 2.910 1.110 4.070 1.280 ;
        RECT 3.900 1.110 4.070 1.650 ;
        RECT 3.945 1.480 4.115 3.060 ;
        RECT 3.900 1.480 4.300 1.650 ;
        RECT 3.945 2.890 4.750 3.060 ;
        RECT 5.025 1.110 5.195 2.360 ;
        RECT 5.025 1.110 6.040 1.280 ;
        RECT 5.025 2.190 6.040 2.360 ;
        RECT 4.295 1.890 4.465 2.710 ;
        RECT 4.260 1.110 4.650 1.280 ;
        RECT 4.480 1.110 4.650 2.070 ;
        RECT 4.295 1.890 4.650 2.070 ;
        RECT 4.295 2.540 6.760 2.710 ;
        RECT 6.590 2.540 6.760 2.915 ;
        RECT 6.590 2.745 7.815 2.915 ;
        RECT 7.645 2.745 7.815 3.045 ;
        RECT 9.105 0.955 9.275 2.280 ;
        RECT 9.040 0.955 9.340 1.125 ;
        RECT 9.105 1.675 10.540 1.845 ;
        RECT 10.450 1.125 10.750 1.495 ;
        RECT 9.760 1.325 11.260 1.495 ;
        RECT 11.090 1.325 11.260 2.215 ;
        RECT 10.420 2.045 11.260 2.215 ;
        RECT 6.250 1.125 7.110 1.295 ;
        RECT 6.250 2.190 7.110 2.360 ;
        RECT 6.940 1.125 7.110 2.565 ;
        RECT 6.940 1.525 7.175 1.825 ;
        RECT 6.940 2.395 8.555 2.565 ;
        RECT 8.385 2.395 8.555 2.980 ;
        RECT 8.385 2.810 11.730 2.980 ;
        RECT 7.355 1.060 7.525 2.215 ;
        RECT 7.355 1.325 8.090 1.495 ;
        RECT 7.355 2.045 8.905 2.215 ;
        RECT 8.735 1.655 8.905 2.630 ;
        RECT 11.440 1.310 11.610 2.630 ;
        RECT 11.440 1.310 11.840 1.480 ;
        RECT 8.735 2.460 12.295 2.630 ;
        RECT 12.125 2.460 12.295 2.795 ;
        RECT 2.305 0.750 2.475 1.650 ;
        RECT 2.175 1.480 2.475 1.650 ;
        RECT 6.040 0.700 6.220 0.930 ;
        RECT 2.305 0.750 6.220 0.930 ;
        RECT 6.040 0.700 7.885 0.880 ;
        RECT 7.705 0.700 7.885 1.090 ;
        RECT 8.575 0.595 8.745 1.090 ;
        RECT 7.705 0.910 8.745 1.090 ;
        RECT 9.520 0.595 9.690 0.945 ;
        RECT 8.575 0.595 9.690 0.775 ;
        RECT 11.395 0.575 11.565 0.945 ;
        RECT 9.520 0.765 11.565 0.945 ;
        RECT 11.395 0.575 12.400 0.760 ;
        RECT 12.660 0.940 12.780 1.480 ;
        RECT 12.660 0.940 13.605 1.110 ;
        RECT 13.435 0.940 13.605 2.215 ;
        RECT 13.180 2.045 13.605 2.215 ;
        RECT 13.435 1.650 13.830 1.820 ;
        RECT 12.480 0.590 12.490 1.480 ;
        RECT 12.490 0.600 12.500 1.480 ;
        RECT 12.500 0.610 12.510 1.480 ;
        RECT 12.510 0.620 12.520 1.480 ;
        RECT 12.520 0.630 12.530 1.480 ;
        RECT 12.530 0.640 12.540 1.480 ;
        RECT 12.540 0.650 12.550 1.480 ;
        RECT 12.550 0.660 12.560 1.480 ;
        RECT 12.560 0.670 12.570 1.480 ;
        RECT 12.570 0.680 12.580 1.480 ;
        RECT 12.580 0.690 12.590 1.480 ;
        RECT 12.590 0.700 12.600 1.480 ;
        RECT 12.600 0.710 12.610 1.480 ;
        RECT 12.610 0.720 12.620 1.480 ;
        RECT 12.620 0.730 12.630 1.480 ;
        RECT 12.630 0.740 12.640 1.480 ;
        RECT 12.640 0.750 12.650 1.480 ;
        RECT 12.650 0.760 12.660 1.480 ;
        RECT 12.475 0.580 12.481 0.834 ;
        RECT 12.400 0.575 12.410 0.759 ;
        RECT 12.410 0.575 12.420 0.769 ;
        RECT 12.420 0.575 12.430 0.779 ;
        RECT 12.430 0.575 12.440 0.789 ;
        RECT 12.440 0.575 12.450 0.799 ;
        RECT 12.450 0.575 12.460 0.809 ;
        RECT 12.460 0.575 12.470 0.819 ;
        RECT 12.470 0.575 12.476 0.829 ;
        RECT 11.790 0.940 12.190 1.110 ;
        RECT 12.020 0.940 12.190 2.215 ;
        RECT 11.800 2.045 12.190 2.215 ;
        RECT 12.830 1.675 13.000 2.650 ;
        RECT 12.020 1.675 13.255 1.845 ;
        RECT 14.475 1.520 14.645 2.650 ;
        RECT 12.830 2.480 14.645 2.650 ;
        RECT 14.475 1.520 14.665 1.820 ;
  END 
END FFSEDHDLXHT

MACRO FFSEDHD2XHT
  CLASS  CORE ;
  FOREIGN FFSEDHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.810 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 15.940 0.720 16.110 1.405 ;
        RECT 15.940 1.235 16.300 1.405 ;
        RECT 16.090 0.720 16.110 2.960 ;
        RECT 15.940 1.960 16.110 2.960 ;
        RECT 16.090 1.235 16.300 2.130 ;
        RECT 15.940 1.960 16.300 2.130 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.860 0.720 15.070 1.405 ;
        RECT 14.860 1.235 15.340 1.405 ;
        RECT 15.170 1.235 15.340 2.235 ;
        RECT 14.835 2.065 15.340 2.235 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.820 1.325 1.130 2.020 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.575 0.580 2.010 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.805 1.545 3.180 2.020 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.675 -0.300 0.975 0.775 ;
        RECT 2.555 -0.300 2.855 0.570 ;
        RECT 3.540 -0.300 3.840 0.570 ;
        RECT 5.310 -0.300 5.610 0.570 ;
        RECT 6.800 -0.300 7.100 0.520 ;
        RECT 8.095 -0.300 8.265 0.730 ;
        RECT 10.020 -0.300 10.320 0.585 ;
        RECT 11.105 -0.300 11.405 0.565 ;
        RECT 13.235 -0.300 13.535 0.470 ;
        RECT 14.315 -0.300 14.615 1.055 ;
        RECT 15.355 -0.300 15.655 1.055 ;
        RECT 16.395 -0.300 16.695 1.055 ;
        RECT 0.000 -0.300 16.810 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 6.250 1.525 6.730 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.565 1.530 6.050 2.010 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.685 2.640 0.985 3.990 ;
        RECT 2.555 2.910 2.855 3.990 ;
        RECT 3.420 2.910 3.720 3.990 ;
        RECT 5.310 2.890 5.610 3.990 ;
        RECT 6.800 3.160 7.100 3.990 ;
        RECT 8.065 2.810 8.235 3.990 ;
        RECT 10.020 3.160 10.320 3.990 ;
        RECT 11.010 3.160 11.310 3.990 ;
        RECT 13.205 2.765 13.505 3.990 ;
        RECT 14.315 2.975 14.615 3.990 ;
        RECT 15.355 2.975 15.655 3.990 ;
        RECT 16.395 2.295 16.695 3.990 ;
        RECT 0.000 3.390 16.810 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.975 0.340 1.345 ;
        RECT 0.170 0.975 1.500 1.145 ;
        RECT 1.330 0.975 1.500 2.375 ;
        RECT 0.105 2.205 1.500 2.375 ;
        RECT 1.330 1.705 1.670 2.005 ;
        RECT 1.680 1.045 2.020 1.345 ;
        RECT 1.850 1.045 2.020 2.875 ;
        RECT 1.680 2.235 2.020 2.875 ;
        RECT 3.710 1.775 3.880 2.730 ;
        RECT 1.680 2.550 3.880 2.730 ;
        RECT 3.360 1.110 3.530 2.370 ;
        RECT 3.030 2.200 3.530 2.370 ;
        RECT 3.030 1.110 4.190 1.280 ;
        RECT 4.020 1.110 4.190 1.650 ;
        RECT 4.065 1.480 4.235 3.060 ;
        RECT 4.020 1.480 4.420 1.650 ;
        RECT 4.065 2.890 4.920 3.060 ;
        RECT 5.115 1.110 5.285 2.360 ;
        RECT 5.115 1.110 6.040 1.280 ;
        RECT 5.115 2.190 6.040 2.360 ;
        RECT 4.415 1.890 4.585 2.710 ;
        RECT 4.370 1.110 4.770 1.280 ;
        RECT 4.600 1.110 4.770 2.070 ;
        RECT 4.415 1.890 4.770 2.070 ;
        RECT 4.415 2.540 6.760 2.710 ;
        RECT 6.590 2.540 6.760 2.980 ;
        RECT 6.590 2.810 7.865 2.980 ;
        RECT 7.695 2.810 7.865 3.110 ;
        RECT 9.135 0.955 9.305 2.280 ;
        RECT 9.070 0.955 9.370 1.125 ;
        RECT 9.135 1.675 10.690 1.845 ;
        RECT 10.600 1.125 10.900 1.495 ;
        RECT 9.790 1.325 11.500 1.495 ;
        RECT 11.330 1.325 11.500 2.215 ;
        RECT 10.570 2.045 11.500 2.215 ;
        RECT 7.355 1.060 7.525 2.150 ;
        RECT 7.415 1.980 7.585 2.280 ;
        RECT 7.355 1.270 7.960 1.440 ;
        RECT 7.355 1.980 8.935 2.150 ;
        RECT 8.765 1.655 8.935 2.630 ;
        RECT 8.765 2.460 12.560 2.630 ;
        RECT 12.390 2.460 12.560 2.795 ;
        RECT 6.250 1.125 7.175 1.295 ;
        RECT 6.250 2.190 7.175 2.360 ;
        RECT 7.005 1.125 7.175 2.630 ;
        RECT 7.005 2.460 8.585 2.630 ;
        RECT 8.415 2.460 8.585 2.980 ;
        RECT 8.415 2.810 12.105 2.980 ;
        RECT 11.935 2.810 12.105 3.210 ;
        RECT 12.475 1.350 12.920 1.520 ;
        RECT 12.740 1.350 12.920 3.210 ;
        RECT 11.935 3.040 12.920 3.210 ;
        RECT 2.360 0.750 2.530 1.825 ;
        RECT 6.745 0.700 6.950 0.930 ;
        RECT 2.360 0.750 6.950 0.930 ;
        RECT 6.745 0.700 7.915 0.880 ;
        RECT 7.735 0.700 7.915 1.090 ;
        RECT 8.620 0.595 8.790 1.090 ;
        RECT 7.735 0.910 8.790 1.090 ;
        RECT 9.600 0.595 9.770 0.945 ;
        RECT 8.620 0.595 9.770 0.775 ;
        RECT 9.600 0.765 11.535 0.945 ;
        RECT 11.735 0.610 13.095 0.820 ;
        RECT 11.735 0.650 14.115 0.820 ;
        RECT 13.785 1.125 14.115 1.295 ;
        RECT 13.945 0.650 14.115 2.225 ;
        RECT 13.755 2.055 14.115 2.225 ;
        RECT 13.945 1.585 14.990 1.885 ;
        RECT 11.690 0.610 11.700 0.854 ;
        RECT 11.700 0.610 11.710 0.844 ;
        RECT 11.710 0.610 11.720 0.834 ;
        RECT 11.720 0.610 11.730 0.824 ;
        RECT 11.730 0.610 11.736 0.820 ;
        RECT 11.610 0.690 11.620 0.934 ;
        RECT 11.620 0.680 11.630 0.924 ;
        RECT 11.630 0.670 11.640 0.914 ;
        RECT 11.640 0.660 11.650 0.904 ;
        RECT 11.650 0.650 11.660 0.894 ;
        RECT 11.660 0.640 11.670 0.884 ;
        RECT 11.670 0.630 11.680 0.874 ;
        RECT 11.680 0.620 11.690 0.864 ;
        RECT 11.535 0.765 11.545 0.945 ;
        RECT 11.545 0.755 11.555 0.945 ;
        RECT 11.555 0.745 11.565 0.945 ;
        RECT 11.565 0.735 11.575 0.945 ;
        RECT 11.575 0.725 11.585 0.945 ;
        RECT 11.585 0.715 11.595 0.945 ;
        RECT 11.595 0.705 11.605 0.945 ;
        RECT 11.605 0.695 11.611 0.945 ;
        RECT 11.915 1.000 12.095 2.240 ;
        RECT 11.915 2.070 12.335 2.240 ;
        RECT 11.915 1.000 13.575 1.170 ;
        RECT 13.405 1.000 13.575 2.585 ;
        RECT 13.405 1.675 13.765 1.845 ;
        RECT 15.590 1.585 15.760 2.585 ;
        RECT 13.405 2.415 15.760 2.585 ;
        RECT 15.590 1.585 15.910 1.755 ;
  END 
END FFSEDHD2XHT

MACRO FFSEDHD1XHT
  CLASS  CORE ;
  FOREIGN FFSEDHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.580 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 15.225 0.720 15.485 1.360 ;
        RECT 15.270 0.720 15.485 2.960 ;
        RECT 15.225 1.980 15.485 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.185 2.000 14.355 2.300 ;
        RECT 14.185 0.720 14.420 1.470 ;
        RECT 14.185 1.265 14.660 1.470 ;
        RECT 14.450 1.265 14.660 2.170 ;
        RECT 14.185 2.000 14.660 2.170 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 1.325 1.220 1.920 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.605 0.640 2.010 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.905 1.500 3.205 2.020 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.775 -0.300 1.075 0.775 ;
        RECT 2.560 -0.300 2.880 0.570 ;
        RECT 3.640 -0.300 3.960 0.570 ;
        RECT 5.410 -0.300 5.710 0.570 ;
        RECT 7.040 -0.300 7.360 0.520 ;
        RECT 8.305 -0.300 8.475 0.730 ;
        RECT 10.110 -0.300 10.410 0.525 ;
        RECT 11.140 -0.300 11.440 0.565 ;
        RECT 13.030 -0.300 13.330 0.695 ;
        RECT 14.640 -0.300 14.940 1.055 ;
        RECT 0.000 -0.300 15.580 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 6.485 1.525 6.935 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.715 1.465 6.130 2.010 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.785 2.640 1.085 3.990 ;
        RECT 2.655 2.910 2.955 3.990 ;
        RECT 3.520 2.910 3.820 3.990 ;
        RECT 5.410 2.890 5.710 3.990 ;
        RECT 7.070 3.095 7.370 3.990 ;
        RECT 8.275 2.810 8.445 3.990 ;
        RECT 10.325 3.160 11.305 3.990 ;
        RECT 13.040 2.830 13.340 3.990 ;
        RECT 14.640 2.975 14.940 3.990 ;
        RECT 0.000 3.390 15.580 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.270 0.975 0.440 1.345 ;
        RECT 0.270 0.975 1.600 1.145 ;
        RECT 1.430 0.975 1.600 2.375 ;
        RECT 0.205 2.205 1.600 2.375 ;
        RECT 1.430 1.705 1.770 2.005 ;
        RECT 1.780 1.045 2.145 1.345 ;
        RECT 1.975 1.045 2.145 2.875 ;
        RECT 1.780 2.235 2.145 2.875 ;
        RECT 3.805 1.775 3.975 2.730 ;
        RECT 1.780 2.550 3.975 2.730 ;
        RECT 3.430 1.110 3.600 2.370 ;
        RECT 3.130 2.200 3.600 2.370 ;
        RECT 3.130 1.110 4.290 1.280 ;
        RECT 4.120 1.110 4.290 1.650 ;
        RECT 4.165 1.480 4.335 3.060 ;
        RECT 4.120 1.480 4.520 1.650 ;
        RECT 4.165 2.890 5.020 3.060 ;
        RECT 5.265 1.110 5.435 2.360 ;
        RECT 5.265 1.110 6.280 1.280 ;
        RECT 5.265 2.190 6.280 2.360 ;
        RECT 4.515 1.890 4.685 2.710 ;
        RECT 4.470 1.110 4.870 1.280 ;
        RECT 4.700 1.110 4.870 2.070 ;
        RECT 4.515 1.890 4.870 2.070 ;
        RECT 4.515 2.540 7.000 2.710 ;
        RECT 6.830 2.540 7.000 2.915 ;
        RECT 6.830 2.745 8.075 2.915 ;
        RECT 7.905 2.745 8.075 3.045 ;
        RECT 9.345 0.955 9.515 2.280 ;
        RECT 9.280 0.955 9.580 1.125 ;
        RECT 9.345 1.675 10.780 1.845 ;
        RECT 10.690 1.125 10.990 1.495 ;
        RECT 10.000 1.325 11.550 1.495 ;
        RECT 11.380 1.325 11.550 2.215 ;
        RECT 10.660 2.045 11.550 2.215 ;
        RECT 6.490 1.125 7.415 1.295 ;
        RECT 6.490 2.190 7.415 2.360 ;
        RECT 7.245 1.125 7.415 2.565 ;
        RECT 7.245 2.395 8.795 2.565 ;
        RECT 8.625 2.395 8.795 2.980 ;
        RECT 8.625 2.810 12.130 2.980 ;
        RECT 7.595 1.060 7.765 2.215 ;
        RECT 7.595 1.325 8.330 1.495 ;
        RECT 7.595 2.045 9.145 2.215 ;
        RECT 8.975 1.655 9.145 2.630 ;
        RECT 11.730 1.310 11.900 2.630 ;
        RECT 11.730 1.310 12.130 1.480 ;
        RECT 8.975 2.460 12.585 2.630 ;
        RECT 12.415 2.460 12.585 2.945 ;
        RECT 2.460 0.750 2.630 1.825 ;
        RECT 6.535 0.700 6.715 0.930 ;
        RECT 2.460 0.750 6.715 0.930 ;
        RECT 6.535 0.700 8.125 0.880 ;
        RECT 7.945 0.700 8.125 1.090 ;
        RECT 8.800 0.595 8.970 1.090 ;
        RECT 7.945 0.910 8.970 1.090 ;
        RECT 8.800 0.595 9.795 0.775 ;
        RECT 10.090 0.765 11.740 0.945 ;
        RECT 12.000 0.575 12.565 0.760 ;
        RECT 12.940 0.935 13.070 1.480 ;
        RECT 12.940 0.935 14.005 1.110 ;
        RECT 13.835 0.935 14.005 2.215 ;
        RECT 13.580 2.045 14.005 2.215 ;
        RECT 13.835 1.650 14.270 1.820 ;
        RECT 12.770 0.715 12.780 1.479 ;
        RECT 12.780 0.725 12.790 1.479 ;
        RECT 12.790 0.735 12.800 1.479 ;
        RECT 12.800 0.745 12.810 1.479 ;
        RECT 12.810 0.755 12.820 1.479 ;
        RECT 12.820 0.765 12.830 1.479 ;
        RECT 12.830 0.775 12.840 1.479 ;
        RECT 12.840 0.785 12.850 1.479 ;
        RECT 12.850 0.795 12.860 1.479 ;
        RECT 12.860 0.805 12.870 1.479 ;
        RECT 12.870 0.815 12.880 1.479 ;
        RECT 12.880 0.825 12.890 1.479 ;
        RECT 12.890 0.835 12.900 1.479 ;
        RECT 12.900 0.845 12.910 1.479 ;
        RECT 12.910 0.855 12.920 1.479 ;
        RECT 12.920 0.865 12.930 1.479 ;
        RECT 12.930 0.875 12.940 1.479 ;
        RECT 12.640 0.585 12.650 0.835 ;
        RECT 12.650 0.595 12.660 0.845 ;
        RECT 12.660 0.605 12.670 0.855 ;
        RECT 12.670 0.615 12.680 0.865 ;
        RECT 12.680 0.625 12.690 0.875 ;
        RECT 12.690 0.635 12.700 0.885 ;
        RECT 12.700 0.645 12.710 0.895 ;
        RECT 12.710 0.655 12.720 0.905 ;
        RECT 12.720 0.665 12.730 0.915 ;
        RECT 12.730 0.675 12.740 0.925 ;
        RECT 12.740 0.685 12.750 0.935 ;
        RECT 12.750 0.695 12.760 0.945 ;
        RECT 12.760 0.705 12.770 0.955 ;
        RECT 12.565 0.575 12.575 0.759 ;
        RECT 12.575 0.575 12.585 0.769 ;
        RECT 12.585 0.575 12.595 0.779 ;
        RECT 12.595 0.575 12.605 0.789 ;
        RECT 12.605 0.575 12.615 0.799 ;
        RECT 12.615 0.575 12.625 0.809 ;
        RECT 12.625 0.575 12.635 0.819 ;
        RECT 12.635 0.575 12.641 0.829 ;
        RECT 11.930 0.575 11.940 0.819 ;
        RECT 11.940 0.575 11.950 0.809 ;
        RECT 11.950 0.575 11.960 0.799 ;
        RECT 11.960 0.575 11.970 0.789 ;
        RECT 11.970 0.575 11.980 0.779 ;
        RECT 11.980 0.575 11.990 0.769 ;
        RECT 11.990 0.575 12.000 0.759 ;
        RECT 11.815 0.690 11.825 0.934 ;
        RECT 11.825 0.680 11.835 0.924 ;
        RECT 11.835 0.670 11.845 0.914 ;
        RECT 11.845 0.660 11.855 0.904 ;
        RECT 11.855 0.650 11.865 0.894 ;
        RECT 11.865 0.640 11.875 0.884 ;
        RECT 11.875 0.630 11.885 0.874 ;
        RECT 11.885 0.620 11.895 0.864 ;
        RECT 11.895 0.610 11.905 0.854 ;
        RECT 11.905 0.600 11.915 0.844 ;
        RECT 11.915 0.590 11.925 0.834 ;
        RECT 11.925 0.580 11.931 0.830 ;
        RECT 11.740 0.765 11.750 0.945 ;
        RECT 11.750 0.755 11.760 0.945 ;
        RECT 11.760 0.745 11.770 0.945 ;
        RECT 11.770 0.735 11.780 0.945 ;
        RECT 11.780 0.725 11.790 0.945 ;
        RECT 11.790 0.715 11.800 0.945 ;
        RECT 11.800 0.705 11.810 0.945 ;
        RECT 11.810 0.695 11.816 0.945 ;
        RECT 9.965 0.650 9.975 0.944 ;
        RECT 9.975 0.660 9.985 0.944 ;
        RECT 9.985 0.670 9.995 0.944 ;
        RECT 9.995 0.680 10.005 0.944 ;
        RECT 10.005 0.690 10.015 0.944 ;
        RECT 10.015 0.700 10.025 0.944 ;
        RECT 10.025 0.710 10.035 0.944 ;
        RECT 10.035 0.720 10.045 0.944 ;
        RECT 10.045 0.730 10.055 0.944 ;
        RECT 10.055 0.740 10.065 0.944 ;
        RECT 10.065 0.750 10.075 0.944 ;
        RECT 10.075 0.760 10.085 0.944 ;
        RECT 10.085 0.765 10.091 0.945 ;
        RECT 9.920 0.605 9.930 0.899 ;
        RECT 9.930 0.615 9.940 0.909 ;
        RECT 9.940 0.625 9.950 0.919 ;
        RECT 9.950 0.635 9.960 0.929 ;
        RECT 9.960 0.640 9.966 0.940 ;
        RECT 9.795 0.595 9.805 0.775 ;
        RECT 9.805 0.595 9.815 0.785 ;
        RECT 9.815 0.595 9.825 0.795 ;
        RECT 9.825 0.595 9.835 0.805 ;
        RECT 9.835 0.595 9.845 0.815 ;
        RECT 9.845 0.595 9.855 0.825 ;
        RECT 9.855 0.595 9.865 0.835 ;
        RECT 9.865 0.595 9.875 0.845 ;
        RECT 9.875 0.595 9.885 0.855 ;
        RECT 9.885 0.595 9.895 0.865 ;
        RECT 9.895 0.595 9.905 0.875 ;
        RECT 9.905 0.595 9.915 0.885 ;
        RECT 9.915 0.595 9.921 0.895 ;
        RECT 12.080 0.940 12.480 1.110 ;
        RECT 12.310 0.940 12.480 2.215 ;
        RECT 12.080 2.045 12.480 2.215 ;
        RECT 13.230 1.675 13.400 2.650 ;
        RECT 12.310 1.675 13.655 1.845 ;
        RECT 14.875 1.520 15.045 2.650 ;
        RECT 13.230 2.480 15.045 2.650 ;
        RECT 14.875 1.520 15.090 1.820 ;
  END 
END FFSEDHD1XHT

MACRO FFSEDCRHDMXHT
  CLASS  CORE ;
  FOREIGN FFSEDCRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.400 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 16.055 1.060 16.300 2.280 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.950 1.125 15.480 1.295 ;
        RECT 15.270 1.125 15.480 2.215 ;
        RECT 14.950 2.045 15.480 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.115 1.265 2.425 1.795 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 2.560 0.990 2.770 ;
        RECT 0.820 2.560 0.990 3.105 ;
        RECT 0.820 2.935 1.525 3.105 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.620 1.590 2.800 2.430 ;
        RECT 2.560 2.085 2.800 2.430 ;
        RECT 2.620 1.590 3.035 1.760 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.775 1.675 6.955 2.360 ;
        RECT 6.550 2.150 6.955 2.360 ;
        RECT 6.775 1.675 7.125 1.975 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.685 ;
        RECT 2.425 -0.300 2.725 0.665 ;
        RECT 3.555 -0.300 3.855 0.550 ;
        RECT 4.615 -0.300 4.915 0.550 ;
        RECT 6.640 -0.300 6.940 0.595 ;
        RECT 8.230 -0.300 8.530 0.595 ;
        RECT 11.100 -0.300 11.400 0.575 ;
        RECT 12.080 -0.300 12.250 1.360 ;
        RECT 13.875 -0.300 14.175 0.770 ;
        RECT 15.500 -0.300 15.800 0.600 ;
        RECT 0.000 -0.300 16.400 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 7.790 1.545 8.220 1.965 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.170 1.515 6.595 1.950 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.405 2.960 0.640 3.990 ;
        RECT 2.545 2.970 3.525 3.990 ;
        RECT 4.780 2.455 5.080 3.990 ;
        RECT 6.690 2.995 6.990 3.990 ;
        RECT 8.230 2.895 8.530 3.990 ;
        RECT 10.945 2.900 11.245 3.990 ;
        RECT 12.015 2.900 12.315 3.990 ;
        RECT 13.885 2.745 14.185 3.990 ;
        RECT 15.500 2.925 15.800 3.990 ;
        RECT 0.000 3.390 16.400 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.010 0.340 2.300 ;
        RECT 0.170 1.585 1.340 1.755 ;
        RECT 1.170 0.605 1.340 2.755 ;
        RECT 1.170 0.605 1.525 0.775 ;
        RECT 1.170 2.585 1.940 2.755 ;
        RECT 1.770 2.585 1.940 2.920 ;
        RECT 2.980 1.125 3.770 1.295 ;
        RECT 3.600 1.125 3.770 2.300 ;
        RECT 2.980 2.000 3.770 2.300 ;
        RECT 1.550 1.010 1.720 2.405 ;
        RECT 1.550 2.225 2.330 2.405 ;
        RECT 2.160 2.225 2.330 2.780 ;
        RECT 2.160 2.610 4.020 2.780 ;
        RECT 3.850 2.610 4.020 3.030 ;
        RECT 3.850 2.860 4.365 3.030 ;
        RECT 4.055 1.125 4.355 1.295 ;
        RECT 4.185 1.125 4.355 1.950 ;
        RECT 4.310 1.780 4.480 2.455 ;
        RECT 5.025 1.645 5.195 1.950 ;
        RECT 4.185 1.780 5.195 1.950 ;
        RECT 5.410 0.830 5.555 3.085 ;
        RECT 5.410 0.830 5.930 1.000 ;
        RECT 5.410 2.915 6.250 3.085 ;
        RECT 6.315 1.125 7.475 1.295 ;
        RECT 7.305 1.125 7.475 2.415 ;
        RECT 7.135 2.245 7.475 2.415 ;
        RECT 6.225 1.045 6.235 1.295 ;
        RECT 6.235 1.055 6.245 1.295 ;
        RECT 6.245 1.065 6.255 1.295 ;
        RECT 6.255 1.075 6.265 1.295 ;
        RECT 6.265 1.085 6.275 1.295 ;
        RECT 6.275 1.095 6.285 1.295 ;
        RECT 6.285 1.105 6.295 1.295 ;
        RECT 6.295 1.115 6.305 1.295 ;
        RECT 6.305 1.125 6.315 1.295 ;
        RECT 6.020 0.840 6.030 1.090 ;
        RECT 6.030 0.850 6.040 1.100 ;
        RECT 6.040 0.860 6.050 1.110 ;
        RECT 6.050 0.870 6.060 1.120 ;
        RECT 6.060 0.880 6.070 1.130 ;
        RECT 6.070 0.890 6.080 1.140 ;
        RECT 6.080 0.900 6.090 1.150 ;
        RECT 6.090 0.910 6.100 1.160 ;
        RECT 6.100 0.920 6.110 1.170 ;
        RECT 6.110 0.930 6.120 1.180 ;
        RECT 6.120 0.940 6.130 1.190 ;
        RECT 6.130 0.950 6.140 1.200 ;
        RECT 6.140 0.960 6.150 1.210 ;
        RECT 6.150 0.970 6.160 1.220 ;
        RECT 6.160 0.980 6.170 1.230 ;
        RECT 6.170 0.990 6.180 1.240 ;
        RECT 6.180 1.000 6.190 1.250 ;
        RECT 6.190 1.010 6.200 1.260 ;
        RECT 6.200 1.020 6.210 1.270 ;
        RECT 6.210 1.030 6.220 1.280 ;
        RECT 6.220 1.035 6.226 1.289 ;
        RECT 5.930 0.830 5.940 1.000 ;
        RECT 5.940 0.830 5.950 1.010 ;
        RECT 5.950 0.830 5.960 1.020 ;
        RECT 5.960 0.830 5.970 1.030 ;
        RECT 5.970 0.830 5.980 1.040 ;
        RECT 5.980 0.830 5.990 1.050 ;
        RECT 5.990 0.830 6.000 1.060 ;
        RECT 6.000 0.830 6.010 1.070 ;
        RECT 6.010 0.830 6.020 1.080 ;
        RECT 5.385 0.855 5.395 3.085 ;
        RECT 5.395 0.845 5.405 3.085 ;
        RECT 5.405 0.835 5.411 3.085 ;
        RECT 7.655 1.125 8.580 1.295 ;
        RECT 8.400 1.125 8.580 2.335 ;
        RECT 7.675 2.165 8.580 2.335 ;
        RECT 8.400 1.535 8.685 1.835 ;
        RECT 8.865 1.125 9.035 2.365 ;
        RECT 8.805 1.125 9.105 1.295 ;
        RECT 5.735 1.235 5.905 2.735 ;
        RECT 6.350 2.605 7.935 2.745 ;
        RECT 6.360 2.605 7.935 2.755 ;
        RECT 6.370 2.605 7.935 2.765 ;
        RECT 5.735 2.565 6.445 2.735 ;
        RECT 5.735 2.575 6.455 2.735 ;
        RECT 5.735 2.585 6.465 2.735 ;
        RECT 5.735 2.595 6.475 2.735 ;
        RECT 7.745 2.545 7.935 2.775 ;
        RECT 6.380 2.605 7.935 2.775 ;
        RECT 9.380 1.135 9.585 1.435 ;
        RECT 7.745 2.545 9.585 2.715 ;
        RECT 9.415 1.135 9.585 2.715 ;
        RECT 10.180 1.200 10.350 2.445 ;
        RECT 10.115 1.200 10.415 1.370 ;
        RECT 10.180 1.930 11.205 2.100 ;
        RECT 11.410 1.685 11.550 1.985 ;
        RECT 11.315 1.685 11.325 2.069 ;
        RECT 11.325 1.685 11.335 2.059 ;
        RECT 11.335 1.685 11.345 2.049 ;
        RECT 11.345 1.685 11.355 2.039 ;
        RECT 11.355 1.685 11.365 2.029 ;
        RECT 11.365 1.685 11.375 2.019 ;
        RECT 11.375 1.685 11.385 2.009 ;
        RECT 11.385 1.685 11.395 1.999 ;
        RECT 11.395 1.685 11.405 1.989 ;
        RECT 11.405 1.685 11.411 1.985 ;
        RECT 11.295 1.840 11.305 2.090 ;
        RECT 11.305 1.830 11.315 2.080 ;
        RECT 11.205 1.930 11.215 2.100 ;
        RECT 11.215 1.920 11.225 2.100 ;
        RECT 11.225 1.910 11.235 2.100 ;
        RECT 11.235 1.900 11.245 2.100 ;
        RECT 11.245 1.890 11.255 2.100 ;
        RECT 11.255 1.880 11.265 2.100 ;
        RECT 11.265 1.870 11.275 2.100 ;
        RECT 11.275 1.860 11.285 2.100 ;
        RECT 11.285 1.850 11.295 2.100 ;
        RECT 3.070 0.490 3.370 0.945 ;
        RECT 3.070 0.775 4.945 0.945 ;
        RECT 5.325 0.480 6.105 0.650 ;
        RECT 6.490 0.775 9.405 0.945 ;
        RECT 9.785 0.480 10.605 0.650 ;
        RECT 11.600 0.510 11.900 0.935 ;
        RECT 10.985 0.765 11.900 0.935 ;
        RECT 10.890 0.680 10.900 0.934 ;
        RECT 10.900 0.690 10.910 0.934 ;
        RECT 10.910 0.700 10.920 0.934 ;
        RECT 10.920 0.710 10.930 0.934 ;
        RECT 10.930 0.720 10.940 0.934 ;
        RECT 10.940 0.730 10.950 0.934 ;
        RECT 10.950 0.740 10.960 0.934 ;
        RECT 10.960 0.750 10.970 0.934 ;
        RECT 10.970 0.760 10.980 0.934 ;
        RECT 10.980 0.765 10.986 0.935 ;
        RECT 10.700 0.490 10.710 0.744 ;
        RECT 10.710 0.500 10.720 0.754 ;
        RECT 10.720 0.510 10.730 0.764 ;
        RECT 10.730 0.520 10.740 0.774 ;
        RECT 10.740 0.530 10.750 0.784 ;
        RECT 10.750 0.540 10.760 0.794 ;
        RECT 10.760 0.550 10.770 0.804 ;
        RECT 10.770 0.560 10.780 0.814 ;
        RECT 10.780 0.570 10.790 0.824 ;
        RECT 10.790 0.580 10.800 0.834 ;
        RECT 10.800 0.590 10.810 0.844 ;
        RECT 10.810 0.600 10.820 0.854 ;
        RECT 10.820 0.610 10.830 0.864 ;
        RECT 10.830 0.620 10.840 0.874 ;
        RECT 10.840 0.630 10.850 0.884 ;
        RECT 10.850 0.640 10.860 0.894 ;
        RECT 10.860 0.650 10.870 0.904 ;
        RECT 10.870 0.660 10.880 0.914 ;
        RECT 10.880 0.670 10.890 0.924 ;
        RECT 10.605 0.480 10.615 0.650 ;
        RECT 10.615 0.480 10.625 0.660 ;
        RECT 10.625 0.480 10.635 0.670 ;
        RECT 10.635 0.480 10.645 0.680 ;
        RECT 10.645 0.480 10.655 0.690 ;
        RECT 10.655 0.480 10.665 0.700 ;
        RECT 10.665 0.480 10.675 0.710 ;
        RECT 10.675 0.480 10.685 0.720 ;
        RECT 10.685 0.480 10.695 0.730 ;
        RECT 10.695 0.480 10.701 0.740 ;
        RECT 9.700 0.480 9.710 0.724 ;
        RECT 9.710 0.480 9.720 0.714 ;
        RECT 9.720 0.480 9.730 0.704 ;
        RECT 9.730 0.480 9.740 0.694 ;
        RECT 9.740 0.480 9.750 0.684 ;
        RECT 9.750 0.480 9.760 0.674 ;
        RECT 9.760 0.480 9.770 0.664 ;
        RECT 9.770 0.480 9.780 0.654 ;
        RECT 9.780 0.480 9.786 0.650 ;
        RECT 9.490 0.690 9.500 0.934 ;
        RECT 9.500 0.680 9.510 0.924 ;
        RECT 9.510 0.670 9.520 0.914 ;
        RECT 9.520 0.660 9.530 0.904 ;
        RECT 9.530 0.650 9.540 0.894 ;
        RECT 9.540 0.640 9.550 0.884 ;
        RECT 9.550 0.630 9.560 0.874 ;
        RECT 9.560 0.620 9.570 0.864 ;
        RECT 9.570 0.610 9.580 0.854 ;
        RECT 9.580 0.600 9.590 0.844 ;
        RECT 9.590 0.590 9.600 0.834 ;
        RECT 9.600 0.580 9.610 0.824 ;
        RECT 9.610 0.570 9.620 0.814 ;
        RECT 9.620 0.560 9.630 0.804 ;
        RECT 9.630 0.550 9.640 0.794 ;
        RECT 9.640 0.540 9.650 0.784 ;
        RECT 9.650 0.530 9.660 0.774 ;
        RECT 9.660 0.520 9.670 0.764 ;
        RECT 9.670 0.510 9.680 0.754 ;
        RECT 9.680 0.500 9.690 0.744 ;
        RECT 9.690 0.490 9.700 0.734 ;
        RECT 9.405 0.775 9.415 0.945 ;
        RECT 9.415 0.765 9.425 0.945 ;
        RECT 9.425 0.755 9.435 0.945 ;
        RECT 9.435 0.745 9.445 0.945 ;
        RECT 9.445 0.735 9.455 0.945 ;
        RECT 9.455 0.725 9.465 0.945 ;
        RECT 9.465 0.715 9.475 0.945 ;
        RECT 9.475 0.705 9.485 0.945 ;
        RECT 9.485 0.695 9.491 0.945 ;
        RECT 6.400 0.695 6.410 0.945 ;
        RECT 6.410 0.705 6.420 0.945 ;
        RECT 6.420 0.715 6.430 0.945 ;
        RECT 6.430 0.725 6.440 0.945 ;
        RECT 6.440 0.735 6.450 0.945 ;
        RECT 6.450 0.745 6.460 0.945 ;
        RECT 6.460 0.755 6.470 0.945 ;
        RECT 6.470 0.765 6.480 0.945 ;
        RECT 6.480 0.775 6.490 0.945 ;
        RECT 6.195 0.490 6.205 0.740 ;
        RECT 6.205 0.500 6.215 0.750 ;
        RECT 6.215 0.510 6.225 0.760 ;
        RECT 6.225 0.520 6.235 0.770 ;
        RECT 6.235 0.530 6.245 0.780 ;
        RECT 6.245 0.540 6.255 0.790 ;
        RECT 6.255 0.550 6.265 0.800 ;
        RECT 6.265 0.560 6.275 0.810 ;
        RECT 6.275 0.570 6.285 0.820 ;
        RECT 6.285 0.580 6.295 0.830 ;
        RECT 6.295 0.590 6.305 0.840 ;
        RECT 6.305 0.600 6.315 0.850 ;
        RECT 6.315 0.610 6.325 0.860 ;
        RECT 6.325 0.620 6.335 0.870 ;
        RECT 6.335 0.630 6.345 0.880 ;
        RECT 6.345 0.640 6.355 0.890 ;
        RECT 6.355 0.650 6.365 0.900 ;
        RECT 6.365 0.660 6.375 0.910 ;
        RECT 6.375 0.670 6.385 0.920 ;
        RECT 6.385 0.680 6.395 0.930 ;
        RECT 6.395 0.685 6.401 0.939 ;
        RECT 6.105 0.480 6.115 0.650 ;
        RECT 6.115 0.480 6.125 0.660 ;
        RECT 6.125 0.480 6.135 0.670 ;
        RECT 6.135 0.480 6.145 0.680 ;
        RECT 6.145 0.480 6.155 0.690 ;
        RECT 6.155 0.480 6.165 0.700 ;
        RECT 6.165 0.480 6.175 0.710 ;
        RECT 6.175 0.480 6.185 0.720 ;
        RECT 6.185 0.480 6.195 0.730 ;
        RECT 5.240 0.480 5.250 0.724 ;
        RECT 5.250 0.480 5.260 0.714 ;
        RECT 5.260 0.480 5.270 0.704 ;
        RECT 5.270 0.480 5.280 0.694 ;
        RECT 5.280 0.480 5.290 0.684 ;
        RECT 5.290 0.480 5.300 0.674 ;
        RECT 5.300 0.480 5.310 0.664 ;
        RECT 5.310 0.480 5.320 0.654 ;
        RECT 5.320 0.480 5.326 0.650 ;
        RECT 5.030 0.690 5.040 0.934 ;
        RECT 5.040 0.680 5.050 0.924 ;
        RECT 5.050 0.670 5.060 0.914 ;
        RECT 5.060 0.660 5.070 0.904 ;
        RECT 5.070 0.650 5.080 0.894 ;
        RECT 5.080 0.640 5.090 0.884 ;
        RECT 5.090 0.630 5.100 0.874 ;
        RECT 5.100 0.620 5.110 0.864 ;
        RECT 5.110 0.610 5.120 0.854 ;
        RECT 5.120 0.600 5.130 0.844 ;
        RECT 5.130 0.590 5.140 0.834 ;
        RECT 5.140 0.580 5.150 0.824 ;
        RECT 5.150 0.570 5.160 0.814 ;
        RECT 5.160 0.560 5.170 0.804 ;
        RECT 5.170 0.550 5.180 0.794 ;
        RECT 5.180 0.540 5.190 0.784 ;
        RECT 5.190 0.530 5.200 0.774 ;
        RECT 5.200 0.520 5.210 0.764 ;
        RECT 5.210 0.510 5.220 0.754 ;
        RECT 5.220 0.500 5.230 0.744 ;
        RECT 5.230 0.490 5.240 0.734 ;
        RECT 4.945 0.775 4.955 0.945 ;
        RECT 4.955 0.765 4.965 0.945 ;
        RECT 4.965 0.755 4.975 0.945 ;
        RECT 4.975 0.745 4.985 0.945 ;
        RECT 4.985 0.735 4.995 0.945 ;
        RECT 4.995 0.725 5.005 0.945 ;
        RECT 5.005 0.715 5.015 0.945 ;
        RECT 5.015 0.705 5.025 0.945 ;
        RECT 5.025 0.695 5.031 0.945 ;
        RECT 10.955 1.125 11.125 1.750 ;
        RECT 10.825 1.580 11.125 1.750 ;
        RECT 10.955 1.125 11.900 1.295 ;
        RECT 11.730 1.125 11.900 2.340 ;
        RECT 11.495 2.170 11.900 2.340 ;
        RECT 11.730 1.610 12.445 1.780 ;
        RECT 8.850 2.895 9.765 3.065 ;
        RECT 10.060 0.830 10.525 1.000 ;
        RECT 10.530 2.530 10.700 2.795 ;
        RECT 9.935 2.625 10.700 2.795 ;
        RECT 10.530 2.530 12.825 2.700 ;
        RECT 12.655 0.710 12.825 2.820 ;
        RECT 12.655 0.710 13.025 0.880 ;
        RECT 12.655 2.650 13.445 2.820 ;
        RECT 9.985 0.830 9.995 1.064 ;
        RECT 9.995 0.830 10.005 1.054 ;
        RECT 10.005 0.830 10.015 1.044 ;
        RECT 10.015 0.830 10.025 1.034 ;
        RECT 10.025 0.830 10.035 1.024 ;
        RECT 10.035 0.830 10.045 1.014 ;
        RECT 10.045 0.830 10.055 1.004 ;
        RECT 10.055 0.830 10.061 1.000 ;
        RECT 9.935 0.880 9.945 1.114 ;
        RECT 9.945 0.870 9.955 1.104 ;
        RECT 9.955 0.860 9.965 1.094 ;
        RECT 9.965 0.850 9.975 1.084 ;
        RECT 9.975 0.840 9.985 1.074 ;
        RECT 9.765 1.050 9.775 3.064 ;
        RECT 9.775 1.040 9.785 3.064 ;
        RECT 9.785 1.030 9.795 3.064 ;
        RECT 9.795 1.020 9.805 3.064 ;
        RECT 9.805 1.010 9.815 3.064 ;
        RECT 9.815 1.000 9.825 3.064 ;
        RECT 9.825 0.990 9.835 3.064 ;
        RECT 9.835 0.980 9.845 3.064 ;
        RECT 9.845 0.970 9.855 3.064 ;
        RECT 9.855 0.960 9.865 3.064 ;
        RECT 9.865 0.950 9.875 3.064 ;
        RECT 9.875 0.940 9.885 3.064 ;
        RECT 9.885 0.930 9.895 3.064 ;
        RECT 9.895 0.920 9.905 3.064 ;
        RECT 9.905 0.910 9.915 3.064 ;
        RECT 9.915 0.900 9.925 3.064 ;
        RECT 9.925 0.890 9.935 3.064 ;
        RECT 14.420 1.125 14.760 1.295 ;
        RECT 14.590 0.480 14.760 2.215 ;
        RECT 14.420 2.045 14.760 2.215 ;
        RECT 14.590 0.480 14.780 0.780 ;
        RECT 14.590 1.665 15.090 1.835 ;
        RECT 13.025 1.060 13.205 2.395 ;
        RECT 13.025 1.060 13.210 1.775 ;
        RECT 13.980 1.605 14.150 2.565 ;
        RECT 13.025 1.605 14.380 1.775 ;
        RECT 15.705 1.530 15.875 2.565 ;
        RECT 13.980 2.395 15.875 2.565 ;
  END 
END FFSEDCRHDMXHT

MACRO FFSEDCRHDLXHT
  CLASS  CORE ;
  FOREIGN FFSEDCRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.400 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 16.055 1.060 16.300 2.280 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.950 1.125 15.480 1.295 ;
        RECT 15.270 1.125 15.480 2.215 ;
        RECT 14.950 2.045 15.480 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.115 1.265 2.440 1.870 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 2.560 0.990 2.770 ;
        RECT 0.820 2.560 0.990 3.105 ;
        RECT 0.820 2.935 1.415 3.105 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.620 1.590 2.800 2.430 ;
        RECT 2.560 2.085 2.800 2.430 ;
        RECT 2.620 1.590 3.015 1.760 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.775 1.675 6.955 2.360 ;
        RECT 6.550 2.150 6.955 2.360 ;
        RECT 6.775 1.675 7.125 1.975 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.685 ;
        RECT 2.425 -0.300 2.725 0.775 ;
        RECT 3.555 -0.300 3.855 0.550 ;
        RECT 4.615 -0.300 4.915 0.550 ;
        RECT 6.640 -0.300 6.940 0.595 ;
        RECT 8.225 -0.300 8.525 0.595 ;
        RECT 11.130 -0.300 11.430 0.575 ;
        RECT 12.200 -0.300 12.370 0.860 ;
        RECT 13.915 -0.300 14.215 0.735 ;
        RECT 15.500 -0.300 15.800 0.750 ;
        RECT 0.000 -0.300 16.400 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 7.790 1.545 8.220 1.965 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.170 1.585 6.595 1.950 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.470 2.950 0.640 3.990 ;
        RECT 2.545 2.970 3.525 3.990 ;
        RECT 4.780 2.360 5.080 3.990 ;
        RECT 6.690 2.995 6.990 3.990 ;
        RECT 8.230 2.895 8.530 3.990 ;
        RECT 11.005 2.900 11.305 3.990 ;
        RECT 12.015 2.900 12.315 3.990 ;
        RECT 13.870 2.745 14.170 3.990 ;
        RECT 15.500 2.745 15.800 3.990 ;
        RECT 0.000 3.390 16.400 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.010 0.340 2.300 ;
        RECT 0.170 1.585 1.340 1.755 ;
        RECT 1.170 0.660 1.340 2.755 ;
        RECT 1.170 0.660 1.525 0.830 ;
        RECT 1.170 2.585 1.940 2.755 ;
        RECT 1.770 2.585 1.940 2.885 ;
        RECT 2.980 1.125 3.770 1.295 ;
        RECT 3.600 1.125 3.770 2.300 ;
        RECT 2.980 2.000 3.770 2.300 ;
        RECT 1.520 1.010 1.690 2.405 ;
        RECT 1.520 1.010 1.720 1.310 ;
        RECT 1.520 2.225 2.330 2.405 ;
        RECT 2.160 2.225 2.330 2.780 ;
        RECT 2.160 2.610 4.020 2.780 ;
        RECT 3.850 2.610 4.020 3.030 ;
        RECT 3.850 2.860 4.365 3.030 ;
        RECT 4.055 1.125 4.355 1.295 ;
        RECT 4.185 1.125 4.355 2.150 ;
        RECT 4.310 1.980 4.480 2.455 ;
        RECT 5.025 1.645 5.195 2.150 ;
        RECT 4.185 1.980 5.195 2.150 ;
        RECT 5.410 0.830 5.555 3.085 ;
        RECT 5.410 0.830 5.930 1.000 ;
        RECT 5.410 2.915 6.250 3.085 ;
        RECT 6.315 1.125 7.475 1.295 ;
        RECT 7.305 1.125 7.475 2.415 ;
        RECT 7.135 2.245 7.475 2.415 ;
        RECT 6.225 1.045 6.235 1.295 ;
        RECT 6.235 1.055 6.245 1.295 ;
        RECT 6.245 1.065 6.255 1.295 ;
        RECT 6.255 1.075 6.265 1.295 ;
        RECT 6.265 1.085 6.275 1.295 ;
        RECT 6.275 1.095 6.285 1.295 ;
        RECT 6.285 1.105 6.295 1.295 ;
        RECT 6.295 1.115 6.305 1.295 ;
        RECT 6.305 1.125 6.315 1.295 ;
        RECT 6.020 0.840 6.030 1.090 ;
        RECT 6.030 0.850 6.040 1.100 ;
        RECT 6.040 0.860 6.050 1.110 ;
        RECT 6.050 0.870 6.060 1.120 ;
        RECT 6.060 0.880 6.070 1.130 ;
        RECT 6.070 0.890 6.080 1.140 ;
        RECT 6.080 0.900 6.090 1.150 ;
        RECT 6.090 0.910 6.100 1.160 ;
        RECT 6.100 0.920 6.110 1.170 ;
        RECT 6.110 0.930 6.120 1.180 ;
        RECT 6.120 0.940 6.130 1.190 ;
        RECT 6.130 0.950 6.140 1.200 ;
        RECT 6.140 0.960 6.150 1.210 ;
        RECT 6.150 0.970 6.160 1.220 ;
        RECT 6.160 0.980 6.170 1.230 ;
        RECT 6.170 0.990 6.180 1.240 ;
        RECT 6.180 1.000 6.190 1.250 ;
        RECT 6.190 1.010 6.200 1.260 ;
        RECT 6.200 1.020 6.210 1.270 ;
        RECT 6.210 1.030 6.220 1.280 ;
        RECT 6.220 1.035 6.226 1.289 ;
        RECT 5.930 0.830 5.940 1.000 ;
        RECT 5.940 0.830 5.950 1.010 ;
        RECT 5.950 0.830 5.960 1.020 ;
        RECT 5.960 0.830 5.970 1.030 ;
        RECT 5.970 0.830 5.980 1.040 ;
        RECT 5.980 0.830 5.990 1.050 ;
        RECT 5.990 0.830 6.000 1.060 ;
        RECT 6.000 0.830 6.010 1.070 ;
        RECT 6.010 0.830 6.020 1.080 ;
        RECT 5.385 0.855 5.395 3.085 ;
        RECT 5.395 0.845 5.405 3.085 ;
        RECT 5.405 0.835 5.411 3.085 ;
        RECT 7.675 1.125 8.580 1.295 ;
        RECT 8.400 1.125 8.580 2.335 ;
        RECT 7.675 2.165 8.580 2.335 ;
        RECT 8.400 1.535 8.685 1.835 ;
        RECT 8.865 1.125 9.035 2.365 ;
        RECT 8.865 2.055 9.045 2.365 ;
        RECT 8.865 2.065 9.055 2.365 ;
        RECT 8.805 1.125 9.105 1.295 ;
        RECT 5.735 1.235 5.905 2.735 ;
        RECT 6.350 2.605 7.935 2.745 ;
        RECT 6.360 2.605 7.935 2.755 ;
        RECT 6.370 2.605 7.935 2.765 ;
        RECT 5.735 2.565 6.445 2.735 ;
        RECT 5.735 2.575 6.455 2.735 ;
        RECT 5.735 2.585 6.465 2.735 ;
        RECT 5.735 2.595 6.475 2.735 ;
        RECT 7.745 2.545 7.935 2.775 ;
        RECT 6.380 2.605 7.935 2.775 ;
        RECT 9.315 1.200 9.615 1.370 ;
        RECT 7.745 2.545 9.615 2.715 ;
        RECT 9.445 1.200 9.615 2.715 ;
        RECT 10.180 1.200 10.350 2.445 ;
        RECT 10.145 1.200 10.445 1.370 ;
        RECT 10.180 1.930 11.210 2.100 ;
        RECT 11.410 1.685 11.550 1.985 ;
        RECT 11.380 1.685 11.390 2.005 ;
        RECT 11.390 1.685 11.400 1.995 ;
        RECT 11.400 1.685 11.410 1.985 ;
        RECT 11.295 1.845 11.305 2.089 ;
        RECT 11.305 1.835 11.315 2.079 ;
        RECT 11.315 1.825 11.325 2.069 ;
        RECT 11.325 1.815 11.335 2.059 ;
        RECT 11.335 1.805 11.345 2.049 ;
        RECT 11.345 1.795 11.355 2.039 ;
        RECT 11.355 1.785 11.365 2.029 ;
        RECT 11.365 1.775 11.375 2.019 ;
        RECT 11.375 1.765 11.381 2.015 ;
        RECT 11.210 1.930 11.220 2.100 ;
        RECT 11.220 1.920 11.230 2.100 ;
        RECT 11.230 1.910 11.240 2.100 ;
        RECT 11.240 1.900 11.250 2.100 ;
        RECT 11.250 1.890 11.260 2.100 ;
        RECT 11.260 1.880 11.270 2.100 ;
        RECT 11.270 1.870 11.280 2.100 ;
        RECT 11.280 1.860 11.290 2.100 ;
        RECT 11.290 1.850 11.296 2.100 ;
        RECT 3.070 0.490 3.370 0.945 ;
        RECT 3.070 0.775 4.945 0.945 ;
        RECT 5.325 0.480 6.105 0.650 ;
        RECT 6.490 0.775 9.545 0.945 ;
        RECT 9.930 0.480 10.665 0.650 ;
        RECT 11.720 0.510 12.020 0.935 ;
        RECT 11.045 0.765 12.020 0.935 ;
        RECT 10.950 0.680 10.960 0.934 ;
        RECT 10.960 0.690 10.970 0.934 ;
        RECT 10.970 0.700 10.980 0.934 ;
        RECT 10.980 0.710 10.990 0.934 ;
        RECT 10.990 0.720 11.000 0.934 ;
        RECT 11.000 0.730 11.010 0.934 ;
        RECT 11.010 0.740 11.020 0.934 ;
        RECT 11.020 0.750 11.030 0.934 ;
        RECT 11.030 0.760 11.040 0.934 ;
        RECT 11.040 0.765 11.046 0.935 ;
        RECT 10.760 0.490 10.770 0.744 ;
        RECT 10.770 0.500 10.780 0.754 ;
        RECT 10.780 0.510 10.790 0.764 ;
        RECT 10.790 0.520 10.800 0.774 ;
        RECT 10.800 0.530 10.810 0.784 ;
        RECT 10.810 0.540 10.820 0.794 ;
        RECT 10.820 0.550 10.830 0.804 ;
        RECT 10.830 0.560 10.840 0.814 ;
        RECT 10.840 0.570 10.850 0.824 ;
        RECT 10.850 0.580 10.860 0.834 ;
        RECT 10.860 0.590 10.870 0.844 ;
        RECT 10.870 0.600 10.880 0.854 ;
        RECT 10.880 0.610 10.890 0.864 ;
        RECT 10.890 0.620 10.900 0.874 ;
        RECT 10.900 0.630 10.910 0.884 ;
        RECT 10.910 0.640 10.920 0.894 ;
        RECT 10.920 0.650 10.930 0.904 ;
        RECT 10.930 0.660 10.940 0.914 ;
        RECT 10.940 0.670 10.950 0.924 ;
        RECT 10.665 0.480 10.675 0.650 ;
        RECT 10.675 0.480 10.685 0.660 ;
        RECT 10.685 0.480 10.695 0.670 ;
        RECT 10.695 0.480 10.705 0.680 ;
        RECT 10.705 0.480 10.715 0.690 ;
        RECT 10.715 0.480 10.725 0.700 ;
        RECT 10.725 0.480 10.735 0.710 ;
        RECT 10.735 0.480 10.745 0.720 ;
        RECT 10.745 0.480 10.755 0.730 ;
        RECT 10.755 0.480 10.761 0.740 ;
        RECT 9.840 0.480 9.850 0.730 ;
        RECT 9.850 0.480 9.860 0.720 ;
        RECT 9.860 0.480 9.870 0.710 ;
        RECT 9.870 0.480 9.880 0.700 ;
        RECT 9.880 0.480 9.890 0.690 ;
        RECT 9.890 0.480 9.900 0.680 ;
        RECT 9.900 0.480 9.910 0.670 ;
        RECT 9.910 0.480 9.920 0.660 ;
        RECT 9.920 0.480 9.930 0.650 ;
        RECT 9.635 0.685 9.645 0.935 ;
        RECT 9.645 0.675 9.655 0.925 ;
        RECT 9.655 0.665 9.665 0.915 ;
        RECT 9.665 0.655 9.675 0.905 ;
        RECT 9.675 0.645 9.685 0.895 ;
        RECT 9.685 0.635 9.695 0.885 ;
        RECT 9.695 0.625 9.705 0.875 ;
        RECT 9.705 0.615 9.715 0.865 ;
        RECT 9.715 0.605 9.725 0.855 ;
        RECT 9.725 0.595 9.735 0.845 ;
        RECT 9.735 0.585 9.745 0.835 ;
        RECT 9.745 0.575 9.755 0.825 ;
        RECT 9.755 0.565 9.765 0.815 ;
        RECT 9.765 0.555 9.775 0.805 ;
        RECT 9.775 0.545 9.785 0.795 ;
        RECT 9.785 0.535 9.795 0.785 ;
        RECT 9.795 0.525 9.805 0.775 ;
        RECT 9.805 0.515 9.815 0.765 ;
        RECT 9.815 0.505 9.825 0.755 ;
        RECT 9.825 0.495 9.835 0.745 ;
        RECT 9.835 0.485 9.841 0.739 ;
        RECT 9.545 0.775 9.555 0.945 ;
        RECT 9.555 0.765 9.565 0.945 ;
        RECT 9.565 0.755 9.575 0.945 ;
        RECT 9.575 0.745 9.585 0.945 ;
        RECT 9.585 0.735 9.595 0.945 ;
        RECT 9.595 0.725 9.605 0.945 ;
        RECT 9.605 0.715 9.615 0.945 ;
        RECT 9.615 0.705 9.625 0.945 ;
        RECT 9.625 0.695 9.635 0.945 ;
        RECT 6.400 0.695 6.410 0.945 ;
        RECT 6.410 0.705 6.420 0.945 ;
        RECT 6.420 0.715 6.430 0.945 ;
        RECT 6.430 0.725 6.440 0.945 ;
        RECT 6.440 0.735 6.450 0.945 ;
        RECT 6.450 0.745 6.460 0.945 ;
        RECT 6.460 0.755 6.470 0.945 ;
        RECT 6.470 0.765 6.480 0.945 ;
        RECT 6.480 0.775 6.490 0.945 ;
        RECT 6.195 0.490 6.205 0.740 ;
        RECT 6.205 0.500 6.215 0.750 ;
        RECT 6.215 0.510 6.225 0.760 ;
        RECT 6.225 0.520 6.235 0.770 ;
        RECT 6.235 0.530 6.245 0.780 ;
        RECT 6.245 0.540 6.255 0.790 ;
        RECT 6.255 0.550 6.265 0.800 ;
        RECT 6.265 0.560 6.275 0.810 ;
        RECT 6.275 0.570 6.285 0.820 ;
        RECT 6.285 0.580 6.295 0.830 ;
        RECT 6.295 0.590 6.305 0.840 ;
        RECT 6.305 0.600 6.315 0.850 ;
        RECT 6.315 0.610 6.325 0.860 ;
        RECT 6.325 0.620 6.335 0.870 ;
        RECT 6.335 0.630 6.345 0.880 ;
        RECT 6.345 0.640 6.355 0.890 ;
        RECT 6.355 0.650 6.365 0.900 ;
        RECT 6.365 0.660 6.375 0.910 ;
        RECT 6.375 0.670 6.385 0.920 ;
        RECT 6.385 0.680 6.395 0.930 ;
        RECT 6.395 0.685 6.401 0.939 ;
        RECT 6.105 0.480 6.115 0.650 ;
        RECT 6.115 0.480 6.125 0.660 ;
        RECT 6.125 0.480 6.135 0.670 ;
        RECT 6.135 0.480 6.145 0.680 ;
        RECT 6.145 0.480 6.155 0.690 ;
        RECT 6.155 0.480 6.165 0.700 ;
        RECT 6.165 0.480 6.175 0.710 ;
        RECT 6.175 0.480 6.185 0.720 ;
        RECT 6.185 0.480 6.195 0.730 ;
        RECT 5.240 0.480 5.250 0.724 ;
        RECT 5.250 0.480 5.260 0.714 ;
        RECT 5.260 0.480 5.270 0.704 ;
        RECT 5.270 0.480 5.280 0.694 ;
        RECT 5.280 0.480 5.290 0.684 ;
        RECT 5.290 0.480 5.300 0.674 ;
        RECT 5.300 0.480 5.310 0.664 ;
        RECT 5.310 0.480 5.320 0.654 ;
        RECT 5.320 0.480 5.326 0.650 ;
        RECT 5.030 0.690 5.040 0.934 ;
        RECT 5.040 0.680 5.050 0.924 ;
        RECT 5.050 0.670 5.060 0.914 ;
        RECT 5.060 0.660 5.070 0.904 ;
        RECT 5.070 0.650 5.080 0.894 ;
        RECT 5.080 0.640 5.090 0.884 ;
        RECT 5.090 0.630 5.100 0.874 ;
        RECT 5.100 0.620 5.110 0.864 ;
        RECT 5.110 0.610 5.120 0.854 ;
        RECT 5.120 0.600 5.130 0.844 ;
        RECT 5.130 0.590 5.140 0.834 ;
        RECT 5.140 0.580 5.150 0.824 ;
        RECT 5.150 0.570 5.160 0.814 ;
        RECT 5.160 0.560 5.170 0.804 ;
        RECT 5.170 0.550 5.180 0.794 ;
        RECT 5.180 0.540 5.190 0.784 ;
        RECT 5.190 0.530 5.200 0.774 ;
        RECT 5.200 0.520 5.210 0.764 ;
        RECT 5.210 0.510 5.220 0.754 ;
        RECT 5.220 0.500 5.230 0.744 ;
        RECT 5.230 0.490 5.240 0.734 ;
        RECT 4.945 0.775 4.955 0.945 ;
        RECT 4.955 0.765 4.965 0.945 ;
        RECT 4.965 0.755 4.975 0.945 ;
        RECT 4.975 0.745 4.985 0.945 ;
        RECT 4.985 0.735 4.995 0.945 ;
        RECT 4.995 0.725 5.005 0.945 ;
        RECT 5.005 0.715 5.015 0.945 ;
        RECT 5.015 0.705 5.025 0.945 ;
        RECT 5.025 0.695 5.031 0.945 ;
        RECT 10.965 1.125 11.135 1.750 ;
        RECT 10.835 1.580 11.135 1.750 ;
        RECT 10.965 1.125 11.900 1.295 ;
        RECT 11.730 1.125 11.900 2.340 ;
        RECT 11.555 2.170 11.900 2.340 ;
        RECT 11.730 1.605 12.445 1.775 ;
        RECT 8.850 2.895 9.795 3.065 ;
        RECT 10.085 0.830 10.585 1.000 ;
        RECT 10.530 2.530 10.700 2.795 ;
        RECT 9.965 2.625 10.700 2.795 ;
        RECT 12.655 0.710 12.825 2.745 ;
        RECT 10.530 2.530 12.825 2.700 ;
        RECT 12.655 0.710 13.025 0.880 ;
        RECT 12.655 2.575 13.475 2.745 ;
        RECT 10.010 0.830 10.020 1.064 ;
        RECT 10.020 0.830 10.030 1.054 ;
        RECT 10.030 0.830 10.040 1.044 ;
        RECT 10.040 0.830 10.050 1.034 ;
        RECT 10.050 0.830 10.060 1.024 ;
        RECT 10.060 0.830 10.070 1.014 ;
        RECT 10.070 0.830 10.080 1.004 ;
        RECT 10.080 0.830 10.086 1.000 ;
        RECT 9.965 0.875 9.975 1.109 ;
        RECT 9.975 0.865 9.985 1.099 ;
        RECT 9.985 0.855 9.995 1.089 ;
        RECT 9.995 0.845 10.005 1.079 ;
        RECT 10.005 0.835 10.011 1.075 ;
        RECT 9.795 1.045 9.805 3.065 ;
        RECT 9.805 1.035 9.815 3.065 ;
        RECT 9.815 1.025 9.825 3.065 ;
        RECT 9.825 1.015 9.835 3.065 ;
        RECT 9.835 1.005 9.845 3.065 ;
        RECT 9.845 0.995 9.855 3.065 ;
        RECT 9.855 0.985 9.865 3.065 ;
        RECT 9.865 0.975 9.875 3.065 ;
        RECT 9.875 0.965 9.885 3.065 ;
        RECT 9.885 0.955 9.895 3.065 ;
        RECT 9.895 0.945 9.905 3.065 ;
        RECT 9.905 0.935 9.915 3.065 ;
        RECT 9.915 0.925 9.925 3.065 ;
        RECT 9.925 0.915 9.935 3.065 ;
        RECT 9.935 0.905 9.945 3.065 ;
        RECT 9.945 0.895 9.955 3.065 ;
        RECT 9.955 0.885 9.965 3.065 ;
        RECT 14.440 1.125 14.760 1.295 ;
        RECT 14.590 0.480 14.760 2.215 ;
        RECT 14.420 2.045 14.760 2.215 ;
        RECT 14.590 0.480 14.780 0.780 ;
        RECT 14.590 1.590 15.090 1.760 ;
        RECT 13.025 1.060 13.205 2.395 ;
        RECT 13.960 1.605 14.130 2.565 ;
        RECT 13.025 1.605 14.380 1.775 ;
        RECT 15.705 1.530 15.875 2.565 ;
        RECT 13.960 2.395 15.875 2.565 ;
  END 
END FFSEDCRHDLXHT

MACRO HAHD2XHT
  CLASS  CORE ;
  FOREIGN HAHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.380 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.240 2.560 0.475 3.020 ;
        RECT 0.240 2.560 0.785 2.915 ;
        RECT 0.240 2.745 4.125 2.915 ;
        RECT 3.955 2.745 4.125 3.100 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.220 1.265 3.590 1.820 ;
    END
  END B
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.365 0.720 5.600 1.360 ;
        RECT 5.430 0.720 5.600 2.215 ;
        RECT 5.430 1.660 5.640 2.215 ;
        RECT 5.300 2.045 5.640 2.215 ;
    END
  END S
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.205 ;
        RECT 3.160 -0.300 3.460 0.595 ;
        RECT 4.845 -0.300 5.020 1.120 ;
        RECT 5.820 -0.300 6.120 1.055 ;
        RECT 6.865 -0.300 7.165 1.055 ;
        RECT 0.000 -0.300 7.380 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 3.095 0.955 3.990 ;
        RECT 3.160 3.095 3.460 3.990 ;
        RECT 4.325 2.835 4.500 3.990 ;
        RECT 4.780 2.975 5.080 3.990 ;
        RECT 5.825 2.975 6.125 3.990 ;
        RECT 6.865 2.295 7.165 3.990 ;
        RECT 0.000 3.390 7.380 3.990 ;
    END
  END VDD
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 6.250 2.085 6.580 2.425 ;
        RECT 6.410 0.720 6.580 2.960 ;
    END
  END CO
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.335 1.755 ;
        RECT 1.165 1.585 1.335 2.565 ;
        RECT 2.165 0.950 2.335 2.565 ;
        RECT 1.165 2.395 2.335 2.565 ;
        RECT 2.515 1.125 2.685 2.215 ;
        RECT 2.515 1.125 2.910 1.295 ;
        RECT 2.515 2.045 2.910 2.215 ;
        RECT 1.640 0.600 1.810 2.215 ;
        RECT 1.575 2.045 1.875 2.215 ;
        RECT 1.640 0.600 2.695 0.770 ;
        RECT 2.525 0.600 2.695 0.945 ;
        RECT 3.735 0.710 3.960 0.945 ;
        RECT 2.525 0.775 3.960 0.945 ;
        RECT 3.735 0.710 4.665 0.880 ;
        RECT 4.495 0.710 4.665 1.755 ;
        RECT 4.495 1.585 5.250 1.755 ;
        RECT 3.710 2.045 4.010 2.555 ;
        RECT 4.145 1.060 4.315 2.215 ;
        RECT 3.710 2.045 4.615 2.215 ;
        RECT 4.445 2.045 4.615 2.620 ;
        RECT 5.895 1.520 6.065 2.620 ;
        RECT 4.445 2.450 6.065 2.620 ;
        RECT 5.895 1.520 6.230 1.820 ;
  END 
END HAHD2XHT

MACRO FFSEDCRHD1XHT
  CLASS  CORE ;
  FOREIGN FFSEDCRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.400 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 16.055 0.720 16.300 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.965 0.720 15.185 1.435 ;
        RECT 14.965 1.265 15.480 1.435 ;
        RECT 15.270 1.265 15.480 2.215 ;
        RECT 14.950 2.045 15.480 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.115 1.265 2.425 1.795 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 2.560 0.990 2.770 ;
        RECT 0.820 2.560 0.990 3.105 ;
        RECT 0.820 2.935 1.525 3.105 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.620 1.590 2.800 2.430 ;
        RECT 2.560 2.085 2.800 2.430 ;
        RECT 2.620 1.590 3.015 1.760 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.775 1.675 6.955 2.360 ;
        RECT 6.550 2.150 6.955 2.360 ;
        RECT 6.775 1.675 7.125 1.975 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.685 ;
        RECT 2.425 -0.300 2.725 1.085 ;
        RECT 3.555 -0.300 3.855 0.550 ;
        RECT 4.615 -0.300 4.915 0.550 ;
        RECT 6.640 -0.300 6.940 0.595 ;
        RECT 8.240 -0.300 8.540 0.595 ;
        RECT 11.100 -0.300 11.400 0.575 ;
        RECT 12.080 -0.300 12.250 1.220 ;
        RECT 13.885 -0.300 14.185 0.735 ;
        RECT 15.470 -0.300 15.770 1.055 ;
        RECT 0.000 -0.300 16.400 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 7.790 1.545 8.220 1.965 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.170 1.515 6.595 1.950 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.405 2.960 0.640 3.990 ;
        RECT 2.545 2.970 3.525 3.990 ;
        RECT 4.780 2.350 5.080 3.990 ;
        RECT 6.690 2.995 6.990 3.990 ;
        RECT 8.230 2.965 8.530 3.990 ;
        RECT 10.945 2.960 11.245 3.990 ;
        RECT 12.015 2.960 12.315 3.990 ;
        RECT 13.885 2.745 14.185 3.990 ;
        RECT 15.470 2.975 15.770 3.990 ;
        RECT 0.000 3.390 16.400 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.010 0.340 2.300 ;
        RECT 0.170 1.585 1.340 1.755 ;
        RECT 1.170 0.605 1.340 2.755 ;
        RECT 1.170 0.605 1.525 0.775 ;
        RECT 1.170 2.585 1.940 2.755 ;
        RECT 1.770 2.585 1.940 3.170 ;
        RECT 2.980 1.125 3.770 1.295 ;
        RECT 3.600 1.125 3.770 2.300 ;
        RECT 2.980 2.000 3.770 2.300 ;
        RECT 1.520 1.010 1.690 2.405 ;
        RECT 1.520 2.225 2.330 2.405 ;
        RECT 2.160 2.225 2.330 2.780 ;
        RECT 2.160 2.610 4.020 2.780 ;
        RECT 3.850 2.610 4.020 3.030 ;
        RECT 3.850 2.860 4.365 3.030 ;
        RECT 4.055 1.125 4.355 1.295 ;
        RECT 4.185 1.125 4.355 2.150 ;
        RECT 4.310 1.980 4.480 2.455 ;
        RECT 5.025 1.645 5.195 2.150 ;
        RECT 4.185 1.980 5.195 2.150 ;
        RECT 5.410 0.830 5.555 3.085 ;
        RECT 5.410 0.830 5.930 1.000 ;
        RECT 5.410 2.915 6.250 3.085 ;
        RECT 6.315 1.125 7.475 1.295 ;
        RECT 7.305 1.125 7.475 2.415 ;
        RECT 7.135 2.245 7.475 2.415 ;
        RECT 6.225 1.045 6.235 1.295 ;
        RECT 6.235 1.055 6.245 1.295 ;
        RECT 6.245 1.065 6.255 1.295 ;
        RECT 6.255 1.075 6.265 1.295 ;
        RECT 6.265 1.085 6.275 1.295 ;
        RECT 6.275 1.095 6.285 1.295 ;
        RECT 6.285 1.105 6.295 1.295 ;
        RECT 6.295 1.115 6.305 1.295 ;
        RECT 6.305 1.125 6.315 1.295 ;
        RECT 6.020 0.840 6.030 1.090 ;
        RECT 6.030 0.850 6.040 1.100 ;
        RECT 6.040 0.860 6.050 1.110 ;
        RECT 6.050 0.870 6.060 1.120 ;
        RECT 6.060 0.880 6.070 1.130 ;
        RECT 6.070 0.890 6.080 1.140 ;
        RECT 6.080 0.900 6.090 1.150 ;
        RECT 6.090 0.910 6.100 1.160 ;
        RECT 6.100 0.920 6.110 1.170 ;
        RECT 6.110 0.930 6.120 1.180 ;
        RECT 6.120 0.940 6.130 1.190 ;
        RECT 6.130 0.950 6.140 1.200 ;
        RECT 6.140 0.960 6.150 1.210 ;
        RECT 6.150 0.970 6.160 1.220 ;
        RECT 6.160 0.980 6.170 1.230 ;
        RECT 6.170 0.990 6.180 1.240 ;
        RECT 6.180 1.000 6.190 1.250 ;
        RECT 6.190 1.010 6.200 1.260 ;
        RECT 6.200 1.020 6.210 1.270 ;
        RECT 6.210 1.030 6.220 1.280 ;
        RECT 6.220 1.035 6.226 1.289 ;
        RECT 5.930 0.830 5.940 1.000 ;
        RECT 5.940 0.830 5.950 1.010 ;
        RECT 5.950 0.830 5.960 1.020 ;
        RECT 5.960 0.830 5.970 1.030 ;
        RECT 5.970 0.830 5.980 1.040 ;
        RECT 5.980 0.830 5.990 1.050 ;
        RECT 5.990 0.830 6.000 1.060 ;
        RECT 6.000 0.830 6.010 1.070 ;
        RECT 6.010 0.830 6.020 1.080 ;
        RECT 5.385 0.855 5.395 3.085 ;
        RECT 5.395 0.845 5.405 3.085 ;
        RECT 5.405 0.835 5.411 3.085 ;
        RECT 7.675 1.125 8.580 1.295 ;
        RECT 8.400 1.125 8.580 2.335 ;
        RECT 7.675 2.165 8.580 2.335 ;
        RECT 8.400 1.535 8.685 1.835 ;
        RECT 8.865 1.125 9.035 2.400 ;
        RECT 8.805 1.125 9.105 1.295 ;
        RECT 5.735 1.235 5.905 2.735 ;
        RECT 6.350 2.605 9.615 2.745 ;
        RECT 6.360 2.605 7.935 2.755 ;
        RECT 6.370 2.605 7.935 2.765 ;
        RECT 5.735 2.565 6.445 2.735 ;
        RECT 5.735 2.575 6.455 2.735 ;
        RECT 5.735 2.585 6.465 2.735 ;
        RECT 5.735 2.595 6.475 2.735 ;
        RECT 7.745 2.580 7.935 2.775 ;
        RECT 6.380 2.605 7.935 2.775 ;
        RECT 9.315 1.220 9.615 1.390 ;
        RECT 7.745 2.580 9.615 2.750 ;
        RECT 9.445 1.220 9.615 2.750 ;
        RECT 10.180 1.220 10.350 2.465 ;
        RECT 10.145 1.220 10.445 1.390 ;
        RECT 10.180 1.950 11.215 2.120 ;
        RECT 11.410 1.715 11.550 2.015 ;
        RECT 11.315 1.715 11.325 2.099 ;
        RECT 11.325 1.715 11.335 2.089 ;
        RECT 11.335 1.715 11.345 2.079 ;
        RECT 11.345 1.715 11.355 2.069 ;
        RECT 11.355 1.715 11.365 2.059 ;
        RECT 11.365 1.715 11.375 2.049 ;
        RECT 11.375 1.715 11.385 2.039 ;
        RECT 11.385 1.715 11.395 2.029 ;
        RECT 11.395 1.715 11.405 2.019 ;
        RECT 11.405 1.715 11.411 2.015 ;
        RECT 11.305 1.860 11.315 2.110 ;
        RECT 11.215 1.950 11.225 2.120 ;
        RECT 11.225 1.940 11.235 2.120 ;
        RECT 11.235 1.930 11.245 2.120 ;
        RECT 11.245 1.920 11.255 2.120 ;
        RECT 11.255 1.910 11.265 2.120 ;
        RECT 11.265 1.900 11.275 2.120 ;
        RECT 11.275 1.890 11.285 2.120 ;
        RECT 11.285 1.880 11.295 2.120 ;
        RECT 11.295 1.870 11.305 2.120 ;
        RECT 3.070 0.490 3.370 0.945 ;
        RECT 3.070 0.775 4.945 0.945 ;
        RECT 5.325 0.480 6.105 0.650 ;
        RECT 9.315 0.500 9.485 0.945 ;
        RECT 6.490 0.775 9.485 0.945 ;
        RECT 9.315 0.500 10.655 0.670 ;
        RECT 11.600 0.510 11.900 0.935 ;
        RECT 11.015 0.765 11.900 0.935 ;
        RECT 10.920 0.680 10.930 0.934 ;
        RECT 10.930 0.690 10.940 0.934 ;
        RECT 10.940 0.700 10.950 0.934 ;
        RECT 10.950 0.710 10.960 0.934 ;
        RECT 10.960 0.720 10.970 0.934 ;
        RECT 10.970 0.730 10.980 0.934 ;
        RECT 10.980 0.740 10.990 0.934 ;
        RECT 10.990 0.750 11.000 0.934 ;
        RECT 11.000 0.760 11.010 0.934 ;
        RECT 11.010 0.765 11.016 0.935 ;
        RECT 10.750 0.510 10.760 0.764 ;
        RECT 10.760 0.520 10.770 0.774 ;
        RECT 10.770 0.530 10.780 0.784 ;
        RECT 10.780 0.540 10.790 0.794 ;
        RECT 10.790 0.550 10.800 0.804 ;
        RECT 10.800 0.560 10.810 0.814 ;
        RECT 10.810 0.570 10.820 0.824 ;
        RECT 10.820 0.580 10.830 0.834 ;
        RECT 10.830 0.590 10.840 0.844 ;
        RECT 10.840 0.600 10.850 0.854 ;
        RECT 10.850 0.610 10.860 0.864 ;
        RECT 10.860 0.620 10.870 0.874 ;
        RECT 10.870 0.630 10.880 0.884 ;
        RECT 10.880 0.640 10.890 0.894 ;
        RECT 10.890 0.650 10.900 0.904 ;
        RECT 10.900 0.660 10.910 0.914 ;
        RECT 10.910 0.670 10.920 0.924 ;
        RECT 10.655 0.500 10.665 0.670 ;
        RECT 10.665 0.500 10.675 0.680 ;
        RECT 10.675 0.500 10.685 0.690 ;
        RECT 10.685 0.500 10.695 0.700 ;
        RECT 10.695 0.500 10.705 0.710 ;
        RECT 10.705 0.500 10.715 0.720 ;
        RECT 10.715 0.500 10.725 0.730 ;
        RECT 10.725 0.500 10.735 0.740 ;
        RECT 10.735 0.500 10.745 0.750 ;
        RECT 10.745 0.500 10.751 0.760 ;
        RECT 6.400 0.695 6.410 0.945 ;
        RECT 6.410 0.705 6.420 0.945 ;
        RECT 6.420 0.715 6.430 0.945 ;
        RECT 6.430 0.725 6.440 0.945 ;
        RECT 6.440 0.735 6.450 0.945 ;
        RECT 6.450 0.745 6.460 0.945 ;
        RECT 6.460 0.755 6.470 0.945 ;
        RECT 6.470 0.765 6.480 0.945 ;
        RECT 6.480 0.775 6.490 0.945 ;
        RECT 6.195 0.490 6.205 0.740 ;
        RECT 6.205 0.500 6.215 0.750 ;
        RECT 6.215 0.510 6.225 0.760 ;
        RECT 6.225 0.520 6.235 0.770 ;
        RECT 6.235 0.530 6.245 0.780 ;
        RECT 6.245 0.540 6.255 0.790 ;
        RECT 6.255 0.550 6.265 0.800 ;
        RECT 6.265 0.560 6.275 0.810 ;
        RECT 6.275 0.570 6.285 0.820 ;
        RECT 6.285 0.580 6.295 0.830 ;
        RECT 6.295 0.590 6.305 0.840 ;
        RECT 6.305 0.600 6.315 0.850 ;
        RECT 6.315 0.610 6.325 0.860 ;
        RECT 6.325 0.620 6.335 0.870 ;
        RECT 6.335 0.630 6.345 0.880 ;
        RECT 6.345 0.640 6.355 0.890 ;
        RECT 6.355 0.650 6.365 0.900 ;
        RECT 6.365 0.660 6.375 0.910 ;
        RECT 6.375 0.670 6.385 0.920 ;
        RECT 6.385 0.680 6.395 0.930 ;
        RECT 6.395 0.685 6.401 0.939 ;
        RECT 6.105 0.480 6.115 0.650 ;
        RECT 6.115 0.480 6.125 0.660 ;
        RECT 6.125 0.480 6.135 0.670 ;
        RECT 6.135 0.480 6.145 0.680 ;
        RECT 6.145 0.480 6.155 0.690 ;
        RECT 6.155 0.480 6.165 0.700 ;
        RECT 6.165 0.480 6.175 0.710 ;
        RECT 6.175 0.480 6.185 0.720 ;
        RECT 6.185 0.480 6.195 0.730 ;
        RECT 5.240 0.480 5.250 0.724 ;
        RECT 5.250 0.480 5.260 0.714 ;
        RECT 5.260 0.480 5.270 0.704 ;
        RECT 5.270 0.480 5.280 0.694 ;
        RECT 5.280 0.480 5.290 0.684 ;
        RECT 5.290 0.480 5.300 0.674 ;
        RECT 5.300 0.480 5.310 0.664 ;
        RECT 5.310 0.480 5.320 0.654 ;
        RECT 5.320 0.480 5.326 0.650 ;
        RECT 5.030 0.690 5.040 0.934 ;
        RECT 5.040 0.680 5.050 0.924 ;
        RECT 5.050 0.670 5.060 0.914 ;
        RECT 5.060 0.660 5.070 0.904 ;
        RECT 5.070 0.650 5.080 0.894 ;
        RECT 5.080 0.640 5.090 0.884 ;
        RECT 5.090 0.630 5.100 0.874 ;
        RECT 5.100 0.620 5.110 0.864 ;
        RECT 5.110 0.610 5.120 0.854 ;
        RECT 5.120 0.600 5.130 0.844 ;
        RECT 5.130 0.590 5.140 0.834 ;
        RECT 5.140 0.580 5.150 0.824 ;
        RECT 5.150 0.570 5.160 0.814 ;
        RECT 5.160 0.560 5.170 0.804 ;
        RECT 5.170 0.550 5.180 0.794 ;
        RECT 5.180 0.540 5.190 0.784 ;
        RECT 5.190 0.530 5.200 0.774 ;
        RECT 5.200 0.520 5.210 0.764 ;
        RECT 5.210 0.510 5.220 0.754 ;
        RECT 5.220 0.500 5.230 0.744 ;
        RECT 5.230 0.490 5.240 0.734 ;
        RECT 4.945 0.775 4.955 0.945 ;
        RECT 4.955 0.765 4.965 0.945 ;
        RECT 4.965 0.755 4.975 0.945 ;
        RECT 4.975 0.745 4.985 0.945 ;
        RECT 4.985 0.735 4.995 0.945 ;
        RECT 4.995 0.725 5.005 0.945 ;
        RECT 5.005 0.715 5.015 0.945 ;
        RECT 5.015 0.705 5.025 0.945 ;
        RECT 5.025 0.695 5.031 0.945 ;
        RECT 10.955 1.125 11.125 1.760 ;
        RECT 10.825 1.590 11.125 1.760 ;
        RECT 10.955 1.125 11.900 1.295 ;
        RECT 11.730 1.125 11.900 2.400 ;
        RECT 11.495 2.230 11.900 2.400 ;
        RECT 11.730 1.570 12.445 1.740 ;
        RECT 9.795 0.850 9.965 3.100 ;
        RECT 8.850 2.930 9.965 3.100 ;
        RECT 9.795 0.850 10.555 1.020 ;
        RECT 10.530 2.590 10.700 2.815 ;
        RECT 9.795 2.645 10.700 2.815 ;
        RECT 10.530 2.590 12.825 2.760 ;
        RECT 12.655 0.615 12.825 3.020 ;
        RECT 12.655 0.615 13.025 0.785 ;
        RECT 12.655 2.850 13.445 3.020 ;
        RECT 14.420 1.125 14.760 1.295 ;
        RECT 14.590 0.480 14.760 2.215 ;
        RECT 14.420 2.045 14.760 2.215 ;
        RECT 14.590 0.480 14.780 0.780 ;
        RECT 14.590 1.665 15.090 1.835 ;
        RECT 13.025 1.060 13.205 2.395 ;
        RECT 13.990 1.605 14.160 2.565 ;
        RECT 13.025 1.605 14.380 1.775 ;
        RECT 15.705 1.530 15.875 2.565 ;
        RECT 13.990 2.395 15.875 2.565 ;
  END 
END FFSEDCRHD1XHT

MACRO FFSDSRHQHDMXHT
  CLASS  CORE ;
  FOREIGN FFSDSRHQHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.170 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.815 1.045 15.070 2.870 ;
        RECT 14.765 1.980 15.070 2.870 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 1.290 1.605 1.540 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.060 1.615 7.510 2.045 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.520 1.735 0.690 2.100 ;
        RECT 0.815 1.930 1.230 2.360 ;
        RECT 1.400 1.735 1.570 2.100 ;
        RECT 0.520 1.930 1.570 2.100 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.995 ;
        RECT 2.435 -0.300 2.735 0.785 ;
        RECT 3.350 -0.300 3.650 0.945 ;
        RECT 7.135 -0.300 7.435 1.130 ;
        RECT 10.390 -0.300 10.560 1.160 ;
        RECT 12.220 -0.300 12.520 0.795 ;
        RECT 14.290 -0.300 14.460 1.345 ;
        RECT 0.000 -0.300 15.170 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.845 1.550 3.275 2.015 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.145 1.415 2.535 2.015 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 13.545 1.540 14.170 1.960 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.905 0.895 3.990 ;
        RECT 2.490 2.895 3.470 3.990 ;
        RECT 4.395 2.895 4.695 3.990 ;
        RECT 7.310 3.025 8.290 3.990 ;
        RECT 10.200 3.025 10.500 3.990 ;
        RECT 12.325 2.315 12.625 3.990 ;
        RECT 14.180 2.895 14.480 3.990 ;
        RECT 0.000 3.390 15.170 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.170 0.340 2.470 ;
        RECT 0.105 0.825 0.275 2.470 ;
        RECT 0.170 2.170 0.340 2.725 ;
        RECT 0.105 0.825 0.405 0.995 ;
        RECT 0.170 2.555 1.305 2.725 ;
        RECT 1.135 2.555 1.305 3.210 ;
        RECT 1.135 3.040 1.995 3.210 ;
        RECT 2.780 1.125 3.770 1.295 ;
        RECT 3.600 1.125 3.770 2.365 ;
        RECT 2.825 2.195 3.770 2.365 ;
        RECT 4.860 0.975 5.430 1.145 ;
        RECT 5.260 0.975 5.430 2.295 ;
        RECT 1.580 0.725 1.750 1.055 ;
        RECT 1.580 0.885 1.965 1.055 ;
        RECT 1.795 0.885 1.965 2.715 ;
        RECT 1.580 2.370 1.965 2.715 ;
        RECT 1.580 2.545 5.780 2.715 ;
        RECT 5.610 0.895 5.780 2.790 ;
        RECT 7.720 0.960 7.920 2.145 ;
        RECT 7.655 0.960 7.955 1.130 ;
        RECT 7.720 1.675 7.985 2.145 ;
        RECT 7.720 1.675 8.495 1.845 ;
        RECT 6.310 0.895 6.480 2.495 ;
        RECT 8.705 1.680 8.875 2.495 ;
        RECT 6.310 2.325 8.875 2.495 ;
        RECT 8.940 1.550 9.110 1.850 ;
        RECT 8.705 1.680 9.110 1.850 ;
        RECT 8.165 0.955 8.465 1.365 ;
        RECT 9.180 0.960 9.350 1.365 ;
        RECT 8.165 1.190 9.350 1.365 ;
        RECT 9.180 0.960 9.860 1.130 ;
        RECT 7.795 0.480 8.095 0.725 ;
        RECT 8.695 0.555 8.995 1.010 ;
        RECT 9.525 1.580 9.695 2.215 ;
        RECT 9.055 2.045 9.695 2.215 ;
        RECT 7.795 0.555 10.210 0.725 ;
        RECT 10.040 0.555 10.210 1.750 ;
        RECT 9.525 1.580 10.755 1.750 ;
        RECT 3.950 0.545 4.155 2.365 ;
        RECT 5.960 0.545 6.130 3.160 ;
        RECT 3.950 0.545 6.725 0.715 ;
        RECT 5.960 2.675 9.505 2.845 ;
        RECT 9.940 2.325 10.810 2.495 ;
        RECT 10.880 2.325 10.885 2.565 ;
        RECT 10.955 2.395 11.635 2.565 ;
        RECT 11.465 2.395 11.635 2.770 ;
        RECT 10.885 2.335 10.895 2.565 ;
        RECT 10.895 2.345 10.905 2.565 ;
        RECT 10.905 2.355 10.915 2.565 ;
        RECT 10.915 2.365 10.925 2.565 ;
        RECT 10.925 2.375 10.935 2.565 ;
        RECT 10.935 2.385 10.945 2.565 ;
        RECT 10.945 2.395 10.955 2.565 ;
        RECT 10.810 2.325 10.820 2.495 ;
        RECT 10.820 2.325 10.830 2.505 ;
        RECT 10.830 2.325 10.840 2.515 ;
        RECT 10.840 2.325 10.850 2.525 ;
        RECT 10.850 2.325 10.860 2.535 ;
        RECT 10.860 2.325 10.870 2.545 ;
        RECT 10.870 2.325 10.880 2.555 ;
        RECT 9.855 2.325 9.865 2.569 ;
        RECT 9.865 2.325 9.875 2.559 ;
        RECT 9.875 2.325 9.885 2.549 ;
        RECT 9.885 2.325 9.895 2.539 ;
        RECT 9.895 2.325 9.905 2.529 ;
        RECT 9.905 2.325 9.915 2.519 ;
        RECT 9.915 2.325 9.925 2.509 ;
        RECT 9.925 2.325 9.935 2.499 ;
        RECT 9.935 2.325 9.941 2.495 ;
        RECT 9.590 2.590 9.600 2.834 ;
        RECT 9.600 2.580 9.610 2.824 ;
        RECT 9.610 2.570 9.620 2.814 ;
        RECT 9.620 2.560 9.630 2.804 ;
        RECT 9.630 2.550 9.640 2.794 ;
        RECT 9.640 2.540 9.650 2.784 ;
        RECT 9.650 2.530 9.660 2.774 ;
        RECT 9.660 2.520 9.670 2.764 ;
        RECT 9.670 2.510 9.680 2.754 ;
        RECT 9.680 2.500 9.690 2.744 ;
        RECT 9.690 2.490 9.700 2.734 ;
        RECT 9.700 2.480 9.710 2.724 ;
        RECT 9.710 2.470 9.720 2.714 ;
        RECT 9.720 2.460 9.730 2.704 ;
        RECT 9.730 2.450 9.740 2.694 ;
        RECT 9.740 2.440 9.750 2.684 ;
        RECT 9.750 2.430 9.760 2.674 ;
        RECT 9.760 2.420 9.770 2.664 ;
        RECT 9.770 2.410 9.780 2.654 ;
        RECT 9.780 2.400 9.790 2.644 ;
        RECT 9.790 2.390 9.800 2.634 ;
        RECT 9.800 2.380 9.810 2.624 ;
        RECT 9.810 2.370 9.820 2.614 ;
        RECT 9.820 2.360 9.830 2.604 ;
        RECT 9.830 2.350 9.840 2.594 ;
        RECT 9.840 2.340 9.850 2.584 ;
        RECT 9.850 2.330 9.856 2.580 ;
        RECT 9.505 2.675 9.515 2.845 ;
        RECT 9.515 2.665 9.525 2.845 ;
        RECT 9.525 2.655 9.535 2.845 ;
        RECT 9.535 2.645 9.545 2.845 ;
        RECT 9.545 2.635 9.555 2.845 ;
        RECT 9.555 2.625 9.565 2.845 ;
        RECT 9.565 2.615 9.575 2.845 ;
        RECT 9.575 2.605 9.585 2.845 ;
        RECT 9.585 2.595 9.591 2.845 ;
        RECT 9.135 3.025 9.680 3.195 ;
        RECT 10.120 2.675 10.585 2.845 ;
        RECT 10.655 2.675 10.675 2.915 ;
        RECT 10.745 2.745 11.195 2.915 ;
        RECT 11.025 2.745 11.195 3.120 ;
        RECT 11.530 1.270 11.830 1.440 ;
        RECT 11.660 1.270 11.830 1.825 ;
        RECT 11.660 1.655 12.030 1.825 ;
        RECT 11.860 1.655 12.030 3.120 ;
        RECT 11.025 2.950 12.030 3.120 ;
        RECT 10.675 2.685 10.685 2.915 ;
        RECT 10.685 2.695 10.695 2.915 ;
        RECT 10.695 2.705 10.705 2.915 ;
        RECT 10.705 2.715 10.715 2.915 ;
        RECT 10.715 2.725 10.725 2.915 ;
        RECT 10.725 2.735 10.735 2.915 ;
        RECT 10.735 2.745 10.745 2.915 ;
        RECT 10.585 2.675 10.595 2.845 ;
        RECT 10.595 2.675 10.605 2.855 ;
        RECT 10.605 2.675 10.615 2.865 ;
        RECT 10.615 2.675 10.625 2.875 ;
        RECT 10.625 2.675 10.635 2.885 ;
        RECT 10.635 2.675 10.645 2.895 ;
        RECT 10.645 2.675 10.655 2.905 ;
        RECT 10.030 2.675 10.040 2.925 ;
        RECT 10.040 2.675 10.050 2.915 ;
        RECT 10.050 2.675 10.060 2.905 ;
        RECT 10.060 2.675 10.070 2.895 ;
        RECT 10.070 2.675 10.080 2.885 ;
        RECT 10.080 2.675 10.090 2.875 ;
        RECT 10.090 2.675 10.100 2.865 ;
        RECT 10.100 2.675 10.110 2.855 ;
        RECT 10.110 2.675 10.120 2.845 ;
        RECT 9.770 2.935 9.780 3.185 ;
        RECT 9.780 2.925 9.790 3.175 ;
        RECT 9.790 2.915 9.800 3.165 ;
        RECT 9.800 2.905 9.810 3.155 ;
        RECT 9.810 2.895 9.820 3.145 ;
        RECT 9.820 2.885 9.830 3.135 ;
        RECT 9.830 2.875 9.840 3.125 ;
        RECT 9.840 2.865 9.850 3.115 ;
        RECT 9.850 2.855 9.860 3.105 ;
        RECT 9.860 2.845 9.870 3.095 ;
        RECT 9.870 2.835 9.880 3.085 ;
        RECT 9.880 2.825 9.890 3.075 ;
        RECT 9.890 2.815 9.900 3.065 ;
        RECT 9.900 2.805 9.910 3.055 ;
        RECT 9.910 2.795 9.920 3.045 ;
        RECT 9.920 2.785 9.930 3.035 ;
        RECT 9.930 2.775 9.940 3.025 ;
        RECT 9.940 2.765 9.950 3.015 ;
        RECT 9.950 2.755 9.960 3.005 ;
        RECT 9.960 2.745 9.970 2.995 ;
        RECT 9.970 2.735 9.980 2.985 ;
        RECT 9.980 2.725 9.990 2.975 ;
        RECT 9.990 2.715 10.000 2.965 ;
        RECT 10.000 2.705 10.010 2.955 ;
        RECT 10.010 2.695 10.020 2.945 ;
        RECT 10.020 2.685 10.030 2.935 ;
        RECT 9.680 3.025 9.690 3.195 ;
        RECT 9.690 3.015 9.700 3.195 ;
        RECT 9.700 3.005 9.710 3.195 ;
        RECT 9.710 2.995 9.720 3.195 ;
        RECT 9.720 2.985 9.730 3.195 ;
        RECT 9.730 2.975 9.740 3.195 ;
        RECT 9.740 2.965 9.750 3.195 ;
        RECT 9.750 2.955 9.760 3.195 ;
        RECT 9.760 2.945 9.770 3.195 ;
        RECT 12.560 1.460 12.730 1.760 ;
        RECT 13.170 1.110 13.345 1.630 ;
        RECT 12.560 1.460 13.345 1.630 ;
        RECT 13.175 1.110 13.345 2.335 ;
        RECT 13.170 1.110 13.470 1.280 ;
        RECT 13.175 2.165 13.870 2.335 ;
        RECT 12.780 0.760 12.950 1.280 ;
        RECT 12.650 1.110 12.950 1.280 ;
        RECT 12.780 0.760 13.860 0.930 ;
        RECT 13.690 0.760 13.860 1.280 ;
        RECT 13.690 1.110 13.990 1.280 ;
        RECT 11.120 0.900 11.290 2.215 ;
        RECT 11.120 2.045 11.420 2.215 ;
        RECT 11.120 0.900 11.905 1.070 ;
        RECT 12.140 1.060 12.380 1.230 ;
        RECT 12.210 1.060 12.380 2.110 ;
        RECT 12.210 1.940 12.975 2.110 ;
        RECT 12.805 1.940 12.975 2.715 ;
        RECT 14.390 1.540 14.560 2.715 ;
        RECT 12.805 2.545 14.560 2.715 ;
        RECT 14.390 1.540 14.635 1.840 ;
        RECT 12.065 0.995 12.075 1.229 ;
        RECT 12.075 1.005 12.085 1.229 ;
        RECT 12.085 1.015 12.095 1.229 ;
        RECT 12.095 1.025 12.105 1.229 ;
        RECT 12.105 1.035 12.115 1.229 ;
        RECT 12.115 1.045 12.125 1.229 ;
        RECT 12.125 1.055 12.135 1.229 ;
        RECT 12.135 1.060 12.141 1.230 ;
        RECT 11.980 0.910 11.990 1.144 ;
        RECT 11.990 0.920 12.000 1.154 ;
        RECT 12.000 0.930 12.010 1.164 ;
        RECT 12.010 0.940 12.020 1.174 ;
        RECT 12.020 0.950 12.030 1.184 ;
        RECT 12.030 0.960 12.040 1.194 ;
        RECT 12.040 0.970 12.050 1.204 ;
        RECT 12.050 0.980 12.060 1.214 ;
        RECT 12.060 0.985 12.066 1.225 ;
        RECT 11.905 0.900 11.915 1.070 ;
        RECT 11.915 0.900 11.925 1.080 ;
        RECT 11.925 0.900 11.935 1.090 ;
        RECT 11.935 0.900 11.945 1.100 ;
        RECT 11.945 0.900 11.955 1.110 ;
        RECT 11.955 0.900 11.965 1.120 ;
        RECT 11.965 0.900 11.975 1.130 ;
        RECT 11.975 0.900 11.981 1.140 ;
  END 
END FFSDSRHQHDMXHT

MACRO FFSDSRHQHD3XHT
  CLASS  CORE ;
  FOREIGN FFSDSRHQHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.910 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 19.530 1.045 19.700 1.390 ;
        RECT 19.530 1.980 19.700 2.960 ;
        RECT 19.530 1.220 20.815 1.390 ;
        RECT 19.530 1.980 20.815 2.335 ;
        RECT 20.570 1.045 20.815 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.445 1.560 1.040 1.955 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.460 1.615 7.910 2.045 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.180 0.755 0.480 0.945 ;
        RECT 1.160 0.550 1.330 0.945 ;
        RECT 0.180 0.775 1.330 0.945 ;
        RECT 1.160 0.550 2.095 0.720 ;
        RECT 0.235 2.555 0.405 2.855 ;
        RECT 0.830 2.145 1.305 2.725 ;
        RECT 0.235 2.555 1.305 2.725 ;
        RECT 1.135 2.145 1.305 3.210 ;
        RECT 1.135 3.040 2.130 3.210 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 -0.300 0.895 0.595 ;
        RECT 2.485 -0.300 2.785 0.620 ;
        RECT 3.475 -0.300 3.775 0.945 ;
        RECT 5.535 -0.300 5.855 0.465 ;
        RECT 7.515 -0.300 7.815 1.130 ;
        RECT 11.495 -0.300 11.665 0.730 ;
        RECT 12.535 -0.300 12.705 0.730 ;
        RECT 14.340 -0.300 14.980 0.665 ;
        RECT 16.985 -0.300 17.285 0.795 ;
        RECT 18.980 -0.300 19.150 0.780 ;
        RECT 19.985 -0.300 20.285 0.990 ;
        RECT 0.000 -0.300 20.910 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.965 1.550 3.465 2.015 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.540 1.490 2.780 2.015 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 18.355 1.525 18.930 1.960 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.975 0.895 3.990 ;
        RECT 2.590 3.075 3.595 3.990 ;
        RECT 4.660 2.985 4.830 3.990 ;
        RECT 7.515 2.995 7.815 3.990 ;
        RECT 8.525 2.995 8.825 3.990 ;
        RECT 10.460 2.920 10.695 3.990 ;
        RECT 11.760 3.010 12.060 3.990 ;
        RECT 17.090 2.315 17.390 3.990 ;
        RECT 18.915 2.895 19.215 3.990 ;
        RECT 19.985 2.635 20.285 3.990 ;
        RECT 0.000 3.390 20.910 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.095 1.125 0.265 2.335 ;
        RECT 0.095 1.125 0.405 1.350 ;
        RECT 0.095 2.160 0.405 2.335 ;
        RECT 0.095 1.180 1.395 1.350 ;
        RECT 1.225 1.180 1.395 1.625 ;
        RECT 1.225 1.455 1.930 1.625 ;
        RECT 1.760 1.455 1.930 1.910 ;
        RECT 2.875 1.125 3.930 1.295 ;
        RECT 3.760 1.125 3.930 2.365 ;
        RECT 2.985 2.195 3.930 2.365 ;
        RECT 4.985 1.055 5.795 1.225 ;
        RECT 5.625 1.055 5.795 2.305 ;
        RECT 5.420 2.135 5.795 2.305 ;
        RECT 1.580 0.950 1.750 1.250 ;
        RECT 1.580 2.275 1.750 2.715 ;
        RECT 1.580 1.075 2.350 1.250 ;
        RECT 2.180 1.075 2.350 2.715 ;
        RECT 3.845 2.600 6.160 2.725 ;
        RECT 3.855 2.600 6.160 2.735 ;
        RECT 3.865 2.600 6.160 2.745 ;
        RECT 3.875 2.600 6.160 2.755 ;
        RECT 3.885 2.600 6.160 2.765 ;
        RECT 3.895 2.600 6.160 2.775 ;
        RECT 3.905 2.600 6.160 2.785 ;
        RECT 1.580 2.545 3.911 2.715 ;
        RECT 1.580 2.555 3.920 2.715 ;
        RECT 1.580 2.565 3.930 2.715 ;
        RECT 1.580 2.575 3.940 2.715 ;
        RECT 1.580 2.585 3.950 2.715 ;
        RECT 3.910 2.600 6.160 2.789 ;
        RECT 1.580 2.595 3.960 2.715 ;
        RECT 5.990 0.995 6.160 2.790 ;
        RECT 3.960 2.600 6.160 2.790 ;
        RECT 6.690 0.895 6.860 2.465 ;
        RECT 9.095 1.975 9.265 2.465 ;
        RECT 6.690 2.295 9.265 2.465 ;
        RECT 9.095 1.975 9.515 2.145 ;
        RECT 8.100 0.895 8.280 1.195 ;
        RECT 8.110 0.895 8.280 2.115 ;
        RECT 8.110 1.615 8.415 2.115 ;
        RECT 8.110 1.615 10.550 1.785 ;
        RECT 10.250 1.615 10.550 1.855 ;
        RECT 8.815 0.510 8.985 1.080 ;
        RECT 9.855 0.510 10.025 1.080 ;
        RECT 8.815 0.510 11.065 0.680 ;
        RECT 10.895 0.510 11.065 1.080 ;
        RECT 10.895 0.910 12.280 1.080 ;
        RECT 8.335 0.480 8.635 0.650 ;
        RECT 8.465 0.480 8.635 1.435 ;
        RECT 9.335 0.890 9.505 1.435 ;
        RECT 9.445 2.395 9.740 2.565 ;
        RECT 10.375 0.890 10.545 1.435 ;
        RECT 10.215 2.045 11.045 2.215 ;
        RECT 8.465 1.265 11.225 1.435 ;
        RECT 11.160 1.265 11.225 2.215 ;
        RECT 11.330 1.265 11.365 1.745 ;
        RECT 11.330 1.575 12.155 1.745 ;
        RECT 12.665 1.140 13.915 1.310 ;
        RECT 14.020 1.140 14.050 1.415 ;
        RECT 14.155 1.245 14.860 1.415 ;
        RECT 14.050 1.150 14.060 1.414 ;
        RECT 14.060 1.160 14.070 1.414 ;
        RECT 14.070 1.170 14.080 1.414 ;
        RECT 14.080 1.180 14.090 1.414 ;
        RECT 14.090 1.190 14.100 1.414 ;
        RECT 14.100 1.200 14.110 1.414 ;
        RECT 14.110 1.210 14.120 1.414 ;
        RECT 14.120 1.220 14.130 1.414 ;
        RECT 14.130 1.230 14.140 1.414 ;
        RECT 14.140 1.240 14.150 1.414 ;
        RECT 14.150 1.245 14.156 1.415 ;
        RECT 13.915 1.140 13.925 1.310 ;
        RECT 13.925 1.140 13.935 1.320 ;
        RECT 13.935 1.140 13.945 1.330 ;
        RECT 13.945 1.140 13.955 1.340 ;
        RECT 13.955 1.140 13.965 1.350 ;
        RECT 13.965 1.140 13.975 1.360 ;
        RECT 13.975 1.140 13.985 1.370 ;
        RECT 13.985 1.140 13.995 1.380 ;
        RECT 13.995 1.140 14.005 1.390 ;
        RECT 14.005 1.140 14.015 1.400 ;
        RECT 14.015 1.140 14.021 1.410 ;
        RECT 12.590 1.140 12.600 1.374 ;
        RECT 12.600 1.140 12.610 1.364 ;
        RECT 12.610 1.140 12.620 1.354 ;
        RECT 12.620 1.140 12.630 1.344 ;
        RECT 12.630 1.140 12.640 1.334 ;
        RECT 12.640 1.140 12.650 1.324 ;
        RECT 12.650 1.140 12.660 1.314 ;
        RECT 12.660 1.140 12.666 1.310 ;
        RECT 12.390 1.340 12.400 1.574 ;
        RECT 12.400 1.330 12.410 1.564 ;
        RECT 12.410 1.320 12.420 1.554 ;
        RECT 12.420 1.310 12.430 1.544 ;
        RECT 12.430 1.300 12.440 1.534 ;
        RECT 12.440 1.290 12.450 1.524 ;
        RECT 12.450 1.280 12.460 1.514 ;
        RECT 12.460 1.270 12.470 1.504 ;
        RECT 12.470 1.260 12.480 1.494 ;
        RECT 12.480 1.250 12.490 1.484 ;
        RECT 12.490 1.240 12.500 1.474 ;
        RECT 12.500 1.230 12.510 1.464 ;
        RECT 12.510 1.220 12.520 1.454 ;
        RECT 12.520 1.210 12.530 1.444 ;
        RECT 12.530 1.200 12.540 1.434 ;
        RECT 12.540 1.190 12.550 1.424 ;
        RECT 12.550 1.180 12.560 1.414 ;
        RECT 12.560 1.170 12.570 1.404 ;
        RECT 12.570 1.160 12.580 1.394 ;
        RECT 12.580 1.150 12.590 1.384 ;
        RECT 12.220 1.510 12.230 1.810 ;
        RECT 12.230 1.500 12.240 1.810 ;
        RECT 12.240 1.490 12.250 1.810 ;
        RECT 12.250 1.480 12.260 1.810 ;
        RECT 12.260 1.470 12.270 1.810 ;
        RECT 12.270 1.460 12.280 1.810 ;
        RECT 12.280 1.450 12.290 1.810 ;
        RECT 12.290 1.440 12.300 1.810 ;
        RECT 12.300 1.430 12.310 1.810 ;
        RECT 12.310 1.420 12.320 1.810 ;
        RECT 12.320 1.410 12.330 1.810 ;
        RECT 12.330 1.400 12.340 1.810 ;
        RECT 12.340 1.390 12.350 1.810 ;
        RECT 12.350 1.380 12.360 1.810 ;
        RECT 12.360 1.370 12.370 1.810 ;
        RECT 12.370 1.360 12.380 1.810 ;
        RECT 12.380 1.350 12.390 1.810 ;
        RECT 12.155 1.575 12.165 1.745 ;
        RECT 12.165 1.565 12.175 1.745 ;
        RECT 12.175 1.555 12.185 1.745 ;
        RECT 12.185 1.545 12.195 1.745 ;
        RECT 12.195 1.535 12.205 1.745 ;
        RECT 12.205 1.525 12.215 1.745 ;
        RECT 12.215 1.515 12.221 1.745 ;
        RECT 11.225 1.265 11.235 2.099 ;
        RECT 11.235 1.265 11.245 2.089 ;
        RECT 11.245 1.265 11.255 2.079 ;
        RECT 11.255 1.265 11.265 2.069 ;
        RECT 11.265 1.265 11.275 2.059 ;
        RECT 11.275 1.265 11.285 2.049 ;
        RECT 11.285 1.265 11.295 2.039 ;
        RECT 11.295 1.265 11.305 2.029 ;
        RECT 11.305 1.265 11.315 2.019 ;
        RECT 11.315 1.265 11.325 2.009 ;
        RECT 11.325 1.265 11.331 2.005 ;
        RECT 11.045 2.045 11.055 2.215 ;
        RECT 11.055 2.035 11.065 2.215 ;
        RECT 11.065 2.025 11.075 2.215 ;
        RECT 11.075 2.015 11.085 2.215 ;
        RECT 11.085 2.005 11.095 2.215 ;
        RECT 11.095 1.995 11.105 2.215 ;
        RECT 11.105 1.985 11.115 2.215 ;
        RECT 11.115 1.975 11.125 2.215 ;
        RECT 11.125 1.965 11.135 2.215 ;
        RECT 11.135 1.955 11.145 2.215 ;
        RECT 11.145 1.945 11.155 2.215 ;
        RECT 11.155 1.935 11.161 2.215 ;
        RECT 10.090 2.045 10.100 2.329 ;
        RECT 10.100 2.045 10.110 2.319 ;
        RECT 10.110 2.045 10.120 2.309 ;
        RECT 10.120 2.045 10.130 2.299 ;
        RECT 10.130 2.045 10.140 2.289 ;
        RECT 10.140 2.045 10.150 2.279 ;
        RECT 10.150 2.045 10.160 2.269 ;
        RECT 10.160 2.045 10.170 2.259 ;
        RECT 10.170 2.045 10.180 2.249 ;
        RECT 10.180 2.045 10.190 2.239 ;
        RECT 10.190 2.045 10.200 2.229 ;
        RECT 10.200 2.045 10.210 2.219 ;
        RECT 10.210 2.045 10.216 2.215 ;
        RECT 9.865 2.270 9.875 2.554 ;
        RECT 9.875 2.260 9.885 2.544 ;
        RECT 9.885 2.250 9.895 2.534 ;
        RECT 9.895 2.240 9.905 2.524 ;
        RECT 9.905 2.230 9.915 2.514 ;
        RECT 9.915 2.220 9.925 2.504 ;
        RECT 9.925 2.210 9.935 2.494 ;
        RECT 9.935 2.200 9.945 2.484 ;
        RECT 9.945 2.190 9.955 2.474 ;
        RECT 9.955 2.180 9.965 2.464 ;
        RECT 9.965 2.170 9.975 2.454 ;
        RECT 9.975 2.160 9.985 2.444 ;
        RECT 9.985 2.150 9.995 2.434 ;
        RECT 9.995 2.140 10.005 2.424 ;
        RECT 10.005 2.130 10.015 2.414 ;
        RECT 10.015 2.120 10.025 2.404 ;
        RECT 10.025 2.110 10.035 2.394 ;
        RECT 10.035 2.100 10.045 2.384 ;
        RECT 10.045 2.090 10.055 2.374 ;
        RECT 10.055 2.080 10.065 2.364 ;
        RECT 10.065 2.070 10.075 2.354 ;
        RECT 10.075 2.060 10.085 2.344 ;
        RECT 10.085 2.050 10.091 2.340 ;
        RECT 9.740 2.395 9.750 2.565 ;
        RECT 9.750 2.385 9.760 2.565 ;
        RECT 9.760 2.375 9.770 2.565 ;
        RECT 9.770 2.365 9.780 2.565 ;
        RECT 9.780 2.355 9.790 2.565 ;
        RECT 9.790 2.345 9.800 2.565 ;
        RECT 9.800 2.335 9.810 2.565 ;
        RECT 9.810 2.325 9.820 2.565 ;
        RECT 9.820 2.315 9.830 2.565 ;
        RECT 9.830 2.305 9.840 2.565 ;
        RECT 9.840 2.295 9.850 2.565 ;
        RECT 9.850 2.285 9.860 2.565 ;
        RECT 9.860 2.275 9.866 2.565 ;
        RECT 12.970 1.850 13.270 2.115 ;
        RECT 12.970 1.945 15.730 2.115 ;
        RECT 4.110 0.645 4.280 2.370 ;
        RECT 4.110 0.645 6.510 0.815 ;
        RECT 6.340 0.545 6.510 3.150 ;
        RECT 5.240 2.980 6.510 3.150 ;
        RECT 6.340 0.545 7.105 0.715 ;
        RECT 6.805 0.510 7.105 0.715 ;
        RECT 6.340 2.645 8.930 2.815 ;
        RECT 9.180 2.815 9.950 2.985 ;
        RECT 10.455 2.435 11.260 2.605 ;
        RECT 11.465 2.305 12.575 2.475 ;
        RECT 12.900 1.490 13.745 1.660 ;
        RECT 15.565 1.340 15.735 1.765 ;
        RECT 13.940 1.595 15.735 1.765 ;
        RECT 12.990 2.645 16.440 2.815 ;
        RECT 13.850 1.515 13.860 1.765 ;
        RECT 13.860 1.525 13.870 1.765 ;
        RECT 13.870 1.535 13.880 1.765 ;
        RECT 13.880 1.545 13.890 1.765 ;
        RECT 13.890 1.555 13.900 1.765 ;
        RECT 13.900 1.565 13.910 1.765 ;
        RECT 13.910 1.575 13.920 1.765 ;
        RECT 13.920 1.585 13.930 1.765 ;
        RECT 13.930 1.595 13.940 1.765 ;
        RECT 13.835 1.500 13.845 1.750 ;
        RECT 13.845 1.505 13.851 1.759 ;
        RECT 13.745 1.490 13.755 1.660 ;
        RECT 13.755 1.490 13.765 1.670 ;
        RECT 13.765 1.490 13.775 1.680 ;
        RECT 13.775 1.490 13.785 1.690 ;
        RECT 13.785 1.490 13.795 1.700 ;
        RECT 13.795 1.490 13.805 1.710 ;
        RECT 13.805 1.490 13.815 1.720 ;
        RECT 13.815 1.490 13.825 1.730 ;
        RECT 13.825 1.490 13.835 1.740 ;
        RECT 12.915 2.580 12.925 2.814 ;
        RECT 12.925 2.590 12.935 2.814 ;
        RECT 12.935 2.600 12.945 2.814 ;
        RECT 12.945 2.610 12.955 2.814 ;
        RECT 12.955 2.620 12.965 2.814 ;
        RECT 12.965 2.630 12.975 2.814 ;
        RECT 12.975 2.640 12.985 2.814 ;
        RECT 12.985 2.645 12.991 2.815 ;
        RECT 12.785 2.450 12.795 2.684 ;
        RECT 12.795 2.460 12.805 2.694 ;
        RECT 12.805 2.470 12.815 2.704 ;
        RECT 12.815 2.480 12.825 2.714 ;
        RECT 12.825 2.490 12.835 2.724 ;
        RECT 12.835 2.500 12.845 2.734 ;
        RECT 12.845 2.510 12.855 2.744 ;
        RECT 12.855 2.520 12.865 2.754 ;
        RECT 12.865 2.530 12.875 2.764 ;
        RECT 12.875 2.540 12.885 2.774 ;
        RECT 12.885 2.550 12.895 2.784 ;
        RECT 12.895 2.560 12.905 2.794 ;
        RECT 12.905 2.570 12.915 2.804 ;
        RECT 12.820 1.490 12.830 1.730 ;
        RECT 12.830 1.490 12.840 1.720 ;
        RECT 12.840 1.490 12.850 1.710 ;
        RECT 12.850 1.490 12.860 1.700 ;
        RECT 12.860 1.490 12.870 1.690 ;
        RECT 12.870 1.490 12.880 1.680 ;
        RECT 12.880 1.490 12.890 1.670 ;
        RECT 12.890 1.490 12.900 1.660 ;
        RECT 12.785 1.525 12.795 1.765 ;
        RECT 12.795 1.515 12.805 1.755 ;
        RECT 12.805 1.505 12.815 1.745 ;
        RECT 12.815 1.495 12.821 1.739 ;
        RECT 12.615 1.695 12.625 2.515 ;
        RECT 12.625 1.685 12.635 2.525 ;
        RECT 12.635 1.675 12.645 2.535 ;
        RECT 12.645 1.665 12.655 2.545 ;
        RECT 12.655 1.655 12.665 2.555 ;
        RECT 12.665 1.645 12.675 2.565 ;
        RECT 12.675 1.635 12.685 2.575 ;
        RECT 12.685 1.625 12.695 2.585 ;
        RECT 12.695 1.615 12.705 2.595 ;
        RECT 12.705 1.605 12.715 2.605 ;
        RECT 12.715 1.595 12.725 2.615 ;
        RECT 12.725 1.585 12.735 2.625 ;
        RECT 12.735 1.575 12.745 2.635 ;
        RECT 12.745 1.565 12.755 2.645 ;
        RECT 12.755 1.555 12.765 2.655 ;
        RECT 12.765 1.545 12.775 2.665 ;
        RECT 12.775 1.535 12.785 2.675 ;
        RECT 12.575 2.305 12.585 2.475 ;
        RECT 12.585 2.305 12.595 2.485 ;
        RECT 12.595 2.305 12.605 2.495 ;
        RECT 12.605 2.305 12.615 2.505 ;
        RECT 11.390 2.305 11.400 2.539 ;
        RECT 11.400 2.305 11.410 2.529 ;
        RECT 11.410 2.305 11.420 2.519 ;
        RECT 11.420 2.305 11.430 2.509 ;
        RECT 11.430 2.305 11.440 2.499 ;
        RECT 11.440 2.305 11.450 2.489 ;
        RECT 11.450 2.305 11.460 2.479 ;
        RECT 11.460 2.305 11.466 2.475 ;
        RECT 11.335 2.360 11.345 2.594 ;
        RECT 11.345 2.350 11.355 2.584 ;
        RECT 11.355 2.340 11.365 2.574 ;
        RECT 11.365 2.330 11.375 2.564 ;
        RECT 11.375 2.320 11.385 2.554 ;
        RECT 11.385 2.310 11.391 2.550 ;
        RECT 11.260 2.435 11.270 2.605 ;
        RECT 11.270 2.425 11.280 2.605 ;
        RECT 11.280 2.415 11.290 2.605 ;
        RECT 11.290 2.405 11.300 2.605 ;
        RECT 11.300 2.395 11.310 2.605 ;
        RECT 11.310 2.385 11.320 2.605 ;
        RECT 11.320 2.375 11.330 2.605 ;
        RECT 11.330 2.365 11.336 2.605 ;
        RECT 10.330 2.435 10.340 2.719 ;
        RECT 10.340 2.435 10.350 2.709 ;
        RECT 10.350 2.435 10.360 2.699 ;
        RECT 10.360 2.435 10.370 2.689 ;
        RECT 10.370 2.435 10.380 2.679 ;
        RECT 10.380 2.435 10.390 2.669 ;
        RECT 10.390 2.435 10.400 2.659 ;
        RECT 10.400 2.435 10.410 2.649 ;
        RECT 10.410 2.435 10.420 2.639 ;
        RECT 10.420 2.435 10.430 2.629 ;
        RECT 10.430 2.435 10.440 2.619 ;
        RECT 10.440 2.435 10.450 2.609 ;
        RECT 10.450 2.435 10.456 2.605 ;
        RECT 10.075 2.690 10.085 2.974 ;
        RECT 10.085 2.680 10.095 2.964 ;
        RECT 10.095 2.670 10.105 2.954 ;
        RECT 10.105 2.660 10.115 2.944 ;
        RECT 10.115 2.650 10.125 2.934 ;
        RECT 10.125 2.640 10.135 2.924 ;
        RECT 10.135 2.630 10.145 2.914 ;
        RECT 10.145 2.620 10.155 2.904 ;
        RECT 10.155 2.610 10.165 2.894 ;
        RECT 10.165 2.600 10.175 2.884 ;
        RECT 10.175 2.590 10.185 2.874 ;
        RECT 10.185 2.580 10.195 2.864 ;
        RECT 10.195 2.570 10.205 2.854 ;
        RECT 10.205 2.560 10.215 2.844 ;
        RECT 10.215 2.550 10.225 2.834 ;
        RECT 10.225 2.540 10.235 2.824 ;
        RECT 10.235 2.530 10.245 2.814 ;
        RECT 10.245 2.520 10.255 2.804 ;
        RECT 10.255 2.510 10.265 2.794 ;
        RECT 10.265 2.500 10.275 2.784 ;
        RECT 10.275 2.490 10.285 2.774 ;
        RECT 10.285 2.480 10.295 2.764 ;
        RECT 10.295 2.470 10.305 2.754 ;
        RECT 10.305 2.460 10.315 2.744 ;
        RECT 10.315 2.450 10.325 2.734 ;
        RECT 10.325 2.440 10.331 2.730 ;
        RECT 9.950 2.815 9.960 2.985 ;
        RECT 9.960 2.805 9.970 2.985 ;
        RECT 9.970 2.795 9.980 2.985 ;
        RECT 9.980 2.785 9.990 2.985 ;
        RECT 9.990 2.775 10.000 2.985 ;
        RECT 10.000 2.765 10.010 2.985 ;
        RECT 10.010 2.755 10.020 2.985 ;
        RECT 10.020 2.745 10.030 2.985 ;
        RECT 10.030 2.735 10.040 2.985 ;
        RECT 10.040 2.725 10.050 2.985 ;
        RECT 10.050 2.715 10.060 2.985 ;
        RECT 10.060 2.705 10.070 2.985 ;
        RECT 10.070 2.695 10.076 2.985 ;
        RECT 9.100 2.745 9.110 2.985 ;
        RECT 9.110 2.755 9.120 2.985 ;
        RECT 9.120 2.765 9.130 2.985 ;
        RECT 9.130 2.775 9.140 2.985 ;
        RECT 9.140 2.785 9.150 2.985 ;
        RECT 9.150 2.795 9.160 2.985 ;
        RECT 9.160 2.805 9.170 2.985 ;
        RECT 9.170 2.815 9.180 2.985 ;
        RECT 9.010 2.655 9.020 2.895 ;
        RECT 9.020 2.665 9.030 2.905 ;
        RECT 9.030 2.675 9.040 2.915 ;
        RECT 9.040 2.685 9.050 2.925 ;
        RECT 9.050 2.695 9.060 2.935 ;
        RECT 9.060 2.705 9.070 2.945 ;
        RECT 9.070 2.715 9.080 2.955 ;
        RECT 9.080 2.725 9.090 2.965 ;
        RECT 9.090 2.735 9.100 2.975 ;
        RECT 8.930 2.645 8.940 2.815 ;
        RECT 8.940 2.645 8.950 2.825 ;
        RECT 8.950 2.645 8.960 2.835 ;
        RECT 8.960 2.645 8.970 2.845 ;
        RECT 8.970 2.645 8.980 2.855 ;
        RECT 8.980 2.645 8.990 2.865 ;
        RECT 8.990 2.645 9.000 2.875 ;
        RECT 9.000 2.645 9.010 2.885 ;
        RECT 10.930 2.995 11.200 3.165 ;
        RECT 11.615 2.655 12.415 2.825 ;
        RECT 12.245 2.655 12.415 3.190 ;
        RECT 16.360 1.320 16.530 1.825 ;
        RECT 16.360 1.655 16.795 1.825 ;
        RECT 16.625 1.655 16.795 3.190 ;
        RECT 12.245 3.020 16.795 3.190 ;
        RECT 11.540 2.655 11.550 2.889 ;
        RECT 11.550 2.655 11.560 2.879 ;
        RECT 11.560 2.655 11.570 2.869 ;
        RECT 11.570 2.655 11.580 2.859 ;
        RECT 11.580 2.655 11.590 2.849 ;
        RECT 11.590 2.655 11.600 2.839 ;
        RECT 11.600 2.655 11.610 2.829 ;
        RECT 11.610 2.655 11.616 2.825 ;
        RECT 11.375 2.820 11.385 3.054 ;
        RECT 11.385 2.810 11.395 3.044 ;
        RECT 11.395 2.800 11.405 3.034 ;
        RECT 11.405 2.790 11.415 3.024 ;
        RECT 11.415 2.780 11.425 3.014 ;
        RECT 11.425 2.770 11.435 3.004 ;
        RECT 11.435 2.760 11.445 2.994 ;
        RECT 11.445 2.750 11.455 2.984 ;
        RECT 11.455 2.740 11.465 2.974 ;
        RECT 11.465 2.730 11.475 2.964 ;
        RECT 11.475 2.720 11.485 2.954 ;
        RECT 11.485 2.710 11.495 2.944 ;
        RECT 11.495 2.700 11.505 2.934 ;
        RECT 11.505 2.690 11.515 2.924 ;
        RECT 11.515 2.680 11.525 2.914 ;
        RECT 11.525 2.670 11.535 2.904 ;
        RECT 11.535 2.660 11.541 2.900 ;
        RECT 11.200 2.995 11.210 3.165 ;
        RECT 11.210 2.985 11.220 3.165 ;
        RECT 11.220 2.975 11.230 3.165 ;
        RECT 11.230 2.965 11.240 3.165 ;
        RECT 11.240 2.955 11.250 3.165 ;
        RECT 11.250 2.945 11.260 3.165 ;
        RECT 11.260 2.935 11.270 3.165 ;
        RECT 11.270 2.925 11.280 3.165 ;
        RECT 11.280 2.915 11.290 3.165 ;
        RECT 11.290 2.905 11.300 3.165 ;
        RECT 11.300 2.895 11.310 3.165 ;
        RECT 11.310 2.885 11.320 3.165 ;
        RECT 11.320 2.875 11.330 3.165 ;
        RECT 11.330 2.865 11.340 3.165 ;
        RECT 11.340 2.855 11.350 3.165 ;
        RECT 11.350 2.845 11.360 3.165 ;
        RECT 11.360 2.835 11.370 3.165 ;
        RECT 11.370 2.825 11.376 3.165 ;
        RECT 17.325 1.460 17.495 1.760 ;
        RECT 18.000 1.110 18.175 1.630 ;
        RECT 17.325 1.460 18.175 1.630 ;
        RECT 18.005 1.110 18.175 2.335 ;
        RECT 17.935 1.110 18.235 1.280 ;
        RECT 18.005 2.165 18.635 2.335 ;
        RECT 17.545 0.760 17.715 1.280 ;
        RECT 17.415 1.110 17.715 1.280 ;
        RECT 17.545 0.760 18.625 0.930 ;
        RECT 18.455 0.760 18.625 1.280 ;
        RECT 18.455 1.110 18.755 1.280 ;
        RECT 13.390 0.785 14.120 0.955 ;
        RECT 14.180 0.785 14.200 1.015 ;
        RECT 16.010 0.845 16.180 2.465 ;
        RECT 13.180 2.295 16.180 2.465 ;
        RECT 15.905 0.845 16.205 1.135 ;
        RECT 16.010 2.115 16.320 2.285 ;
        RECT 14.260 0.845 16.615 1.015 ;
        RECT 16.905 1.060 17.145 1.230 ;
        RECT 16.975 1.060 17.145 2.110 ;
        RECT 16.975 1.940 17.755 2.110 ;
        RECT 17.585 1.940 17.755 2.715 ;
        RECT 19.155 1.570 19.325 2.715 ;
        RECT 17.585 2.545 19.325 2.715 ;
        RECT 19.155 1.570 20.355 1.740 ;
        RECT 16.830 0.995 16.840 1.229 ;
        RECT 16.840 1.005 16.850 1.229 ;
        RECT 16.850 1.015 16.860 1.229 ;
        RECT 16.860 1.025 16.870 1.229 ;
        RECT 16.870 1.035 16.880 1.229 ;
        RECT 16.880 1.045 16.890 1.229 ;
        RECT 16.890 1.055 16.900 1.229 ;
        RECT 16.900 1.060 16.906 1.230 ;
        RECT 16.690 0.855 16.700 1.089 ;
        RECT 16.700 0.865 16.710 1.099 ;
        RECT 16.710 0.875 16.720 1.109 ;
        RECT 16.720 0.885 16.730 1.119 ;
        RECT 16.730 0.895 16.740 1.129 ;
        RECT 16.740 0.905 16.750 1.139 ;
        RECT 16.750 0.915 16.760 1.149 ;
        RECT 16.760 0.925 16.770 1.159 ;
        RECT 16.770 0.935 16.780 1.169 ;
        RECT 16.780 0.945 16.790 1.179 ;
        RECT 16.790 0.955 16.800 1.189 ;
        RECT 16.800 0.965 16.810 1.199 ;
        RECT 16.810 0.975 16.820 1.209 ;
        RECT 16.820 0.985 16.830 1.219 ;
        RECT 16.615 0.845 16.625 1.015 ;
        RECT 16.625 0.845 16.635 1.025 ;
        RECT 16.635 0.845 16.645 1.035 ;
        RECT 16.645 0.845 16.655 1.045 ;
        RECT 16.655 0.845 16.665 1.055 ;
        RECT 16.665 0.845 16.675 1.065 ;
        RECT 16.675 0.845 16.685 1.075 ;
        RECT 16.685 0.845 16.691 1.085 ;
        RECT 14.200 0.795 14.210 1.015 ;
        RECT 14.210 0.805 14.220 1.015 ;
        RECT 14.220 0.815 14.230 1.015 ;
        RECT 14.230 0.825 14.240 1.015 ;
        RECT 14.240 0.835 14.250 1.015 ;
        RECT 14.250 0.845 14.260 1.015 ;
        RECT 14.120 0.785 14.130 0.955 ;
        RECT 14.130 0.785 14.140 0.965 ;
        RECT 14.140 0.785 14.150 0.975 ;
        RECT 14.150 0.785 14.160 0.985 ;
        RECT 14.160 0.785 14.170 0.995 ;
        RECT 14.170 0.785 14.180 1.005 ;
  END 
END FFSDSRHQHD3XHT

MACRO FFSDSRHQHD2XHT
  CLASS  CORE ;
  FOREIGN FFSDSRHQHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.860 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 17.935 0.725 18.320 1.300 ;
        RECT 18.050 0.725 18.235 2.965 ;
        RECT 18.000 1.985 18.235 2.965 ;
        RECT 18.050 0.725 18.320 2.425 ;
        RECT 18.000 1.985 18.350 2.425 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.445 1.560 1.040 1.955 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.060 1.615 7.605 2.045 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.235 2.555 0.405 2.855 ;
        RECT 0.830 2.145 1.305 2.725 ;
        RECT 0.235 2.555 1.305 2.725 ;
        RECT 1.135 2.145 1.305 3.210 ;
        RECT 1.135 3.040 2.130 3.210 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.995 ;
        RECT 2.435 -0.300 2.735 0.785 ;
        RECT 3.400 -0.300 3.700 0.945 ;
        RECT 7.210 -0.300 7.510 1.130 ;
        RECT 12.020 -0.300 12.190 0.730 ;
        RECT 15.455 -0.300 15.755 0.800 ;
        RECT 17.480 -0.300 17.650 0.780 ;
        RECT 18.520 -0.300 18.690 1.120 ;
        RECT 0.000 -0.300 18.860 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.965 1.550 3.390 2.015 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.490 1.475 2.780 2.015 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 16.825 1.530 17.400 1.965 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.945 0.895 3.990 ;
        RECT 2.540 2.950 3.520 3.990 ;
        RECT 4.480 2.950 4.780 3.990 ;
        RECT 7.210 3.025 7.510 3.990 ;
        RECT 8.195 3.025 8.495 3.990 ;
        RECT 10.040 3.025 10.340 3.990 ;
        RECT 11.390 3.015 11.690 3.990 ;
        RECT 15.560 2.320 15.860 3.990 ;
        RECT 17.415 2.975 17.715 3.990 ;
        RECT 18.520 2.570 18.690 3.990 ;
        RECT 0.000 3.390 18.860 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.095 0.825 0.265 2.335 ;
        RECT 0.095 0.825 0.405 0.995 ;
        RECT 0.095 2.160 0.405 2.335 ;
        RECT 0.095 1.180 1.395 1.350 ;
        RECT 1.225 1.180 1.395 1.560 ;
        RECT 1.225 1.390 1.930 1.560 ;
        RECT 1.760 1.390 1.930 1.690 ;
        RECT 2.830 1.125 3.855 1.295 ;
        RECT 3.685 1.125 3.855 2.365 ;
        RECT 2.910 2.195 3.855 2.365 ;
        RECT 4.910 1.200 5.210 1.515 ;
        RECT 5.345 1.345 5.515 2.355 ;
        RECT 4.910 1.345 5.580 1.515 ;
        RECT 1.580 0.725 1.750 1.195 ;
        RECT 1.580 2.175 1.750 2.770 ;
        RECT 1.580 1.025 2.300 1.195 ;
        RECT 2.130 1.025 2.300 2.770 ;
        RECT 4.505 0.850 4.675 2.770 ;
        RECT 4.505 0.850 5.845 1.020 ;
        RECT 1.580 2.600 5.845 2.770 ;
        RECT 5.675 0.850 5.845 1.150 ;
        RECT 5.675 2.565 5.845 2.865 ;
        RECT 7.795 0.970 7.965 2.125 ;
        RECT 7.795 1.675 8.115 2.125 ;
        RECT 7.795 1.675 8.575 1.845 ;
        RECT 6.385 0.895 6.555 2.475 ;
        RECT 8.765 1.675 8.935 2.475 ;
        RECT 6.385 2.305 8.935 2.475 ;
        RECT 8.765 1.675 10.485 1.845 ;
        RECT 8.500 0.580 8.670 1.140 ;
        RECT 9.550 0.580 9.720 1.140 ;
        RECT 10.590 0.580 10.760 1.140 ;
        RECT 8.500 0.580 11.800 0.750 ;
        RECT 11.630 0.580 11.800 1.235 ;
        RECT 7.910 0.485 8.320 0.655 ;
        RECT 8.150 0.485 8.320 1.490 ;
        RECT 9.030 0.950 9.200 1.490 ;
        RECT 10.070 0.950 10.240 1.490 ;
        RECT 9.120 2.045 10.720 2.215 ;
        RECT 8.150 1.320 10.900 1.490 ;
        RECT 10.830 1.320 10.900 2.215 ;
        RECT 11.000 1.320 11.035 1.750 ;
        RECT 11.000 1.580 11.730 1.750 ;
        RECT 12.390 0.725 12.560 1.200 ;
        RECT 12.185 1.030 12.560 1.200 ;
        RECT 12.390 0.725 14.280 0.895 ;
        RECT 14.110 0.725 14.280 1.025 ;
        RECT 12.015 1.030 12.025 1.544 ;
        RECT 12.025 1.030 12.035 1.534 ;
        RECT 12.035 1.030 12.045 1.524 ;
        RECT 12.045 1.030 12.055 1.514 ;
        RECT 12.055 1.030 12.065 1.504 ;
        RECT 12.065 1.030 12.075 1.494 ;
        RECT 12.075 1.030 12.085 1.484 ;
        RECT 12.085 1.030 12.095 1.474 ;
        RECT 12.095 1.030 12.105 1.464 ;
        RECT 12.105 1.030 12.115 1.454 ;
        RECT 12.115 1.030 12.125 1.444 ;
        RECT 12.125 1.030 12.135 1.434 ;
        RECT 12.135 1.030 12.145 1.424 ;
        RECT 12.145 1.030 12.155 1.414 ;
        RECT 12.155 1.030 12.165 1.404 ;
        RECT 12.165 1.030 12.175 1.394 ;
        RECT 12.175 1.030 12.185 1.384 ;
        RECT 12.010 1.300 12.016 1.554 ;
        RECT 11.730 1.580 11.740 1.750 ;
        RECT 11.740 1.570 11.750 1.750 ;
        RECT 11.750 1.560 11.760 1.750 ;
        RECT 11.760 1.550 11.770 1.750 ;
        RECT 11.770 1.540 11.780 1.750 ;
        RECT 11.780 1.530 11.790 1.750 ;
        RECT 11.790 1.520 11.800 1.750 ;
        RECT 11.800 1.510 11.810 1.750 ;
        RECT 11.810 1.500 11.820 1.750 ;
        RECT 11.820 1.490 11.830 1.750 ;
        RECT 11.830 1.480 11.840 1.750 ;
        RECT 11.840 1.470 11.850 1.750 ;
        RECT 11.850 1.460 11.860 1.750 ;
        RECT 11.860 1.450 11.870 1.750 ;
        RECT 11.870 1.440 11.880 1.750 ;
        RECT 11.880 1.430 11.890 1.750 ;
        RECT 11.890 1.420 11.900 1.750 ;
        RECT 11.900 1.410 11.910 1.750 ;
        RECT 11.910 1.400 11.920 1.750 ;
        RECT 11.920 1.390 11.930 1.750 ;
        RECT 11.930 1.380 11.940 1.750 ;
        RECT 11.940 1.370 11.950 1.750 ;
        RECT 11.950 1.360 11.960 1.750 ;
        RECT 11.960 1.350 11.970 1.750 ;
        RECT 11.970 1.340 11.980 1.750 ;
        RECT 11.980 1.330 11.990 1.750 ;
        RECT 11.990 1.320 12.000 1.750 ;
        RECT 12.000 1.310 12.010 1.750 ;
        RECT 10.900 1.320 10.910 2.100 ;
        RECT 10.910 1.320 10.920 2.090 ;
        RECT 10.920 1.320 10.930 2.080 ;
        RECT 10.930 1.320 10.940 2.070 ;
        RECT 10.940 1.320 10.950 2.060 ;
        RECT 10.950 1.320 10.960 2.050 ;
        RECT 10.960 1.320 10.970 2.040 ;
        RECT 10.970 1.320 10.980 2.030 ;
        RECT 10.980 1.320 10.990 2.020 ;
        RECT 10.990 1.320 11.000 2.010 ;
        RECT 10.720 2.045 10.730 2.215 ;
        RECT 10.730 2.035 10.740 2.215 ;
        RECT 10.740 2.025 10.750 2.215 ;
        RECT 10.750 2.015 10.760 2.215 ;
        RECT 10.760 2.005 10.770 2.215 ;
        RECT 10.770 1.995 10.780 2.215 ;
        RECT 10.780 1.985 10.790 2.215 ;
        RECT 10.790 1.975 10.800 2.215 ;
        RECT 10.800 1.965 10.810 2.215 ;
        RECT 10.810 1.955 10.820 2.215 ;
        RECT 10.820 1.945 10.830 2.215 ;
        RECT 12.570 1.835 12.870 2.025 ;
        RECT 14.000 1.835 14.300 2.025 ;
        RECT 12.570 1.855 14.300 2.025 ;
        RECT 4.035 0.500 4.205 2.365 ;
        RECT 6.035 0.500 6.205 3.210 ;
        RECT 6.035 2.670 6.270 3.210 ;
        RECT 4.035 0.500 6.800 0.670 ;
        RECT 6.035 2.670 9.500 2.840 ;
        RECT 9.775 2.485 10.900 2.655 ;
        RECT 11.145 2.315 12.190 2.485 ;
        RECT 12.495 1.470 13.355 1.640 ;
        RECT 13.055 1.470 13.355 1.665 ;
        RECT 12.595 2.645 14.910 2.815 ;
        RECT 12.520 2.580 12.530 2.814 ;
        RECT 12.530 2.590 12.540 2.814 ;
        RECT 12.540 2.600 12.550 2.814 ;
        RECT 12.550 2.610 12.560 2.814 ;
        RECT 12.560 2.620 12.570 2.814 ;
        RECT 12.570 2.630 12.580 2.814 ;
        RECT 12.580 2.640 12.590 2.814 ;
        RECT 12.590 2.645 12.596 2.815 ;
        RECT 12.390 2.450 12.400 2.684 ;
        RECT 12.400 2.460 12.410 2.694 ;
        RECT 12.410 2.470 12.420 2.704 ;
        RECT 12.420 2.480 12.430 2.714 ;
        RECT 12.430 2.490 12.440 2.724 ;
        RECT 12.440 2.500 12.450 2.734 ;
        RECT 12.450 2.510 12.460 2.744 ;
        RECT 12.460 2.520 12.470 2.754 ;
        RECT 12.470 2.530 12.480 2.764 ;
        RECT 12.480 2.540 12.490 2.774 ;
        RECT 12.490 2.550 12.500 2.784 ;
        RECT 12.500 2.560 12.510 2.794 ;
        RECT 12.510 2.570 12.520 2.804 ;
        RECT 12.420 1.470 12.430 1.704 ;
        RECT 12.430 1.470 12.440 1.694 ;
        RECT 12.440 1.470 12.450 1.684 ;
        RECT 12.450 1.470 12.460 1.674 ;
        RECT 12.460 1.470 12.470 1.664 ;
        RECT 12.470 1.470 12.480 1.654 ;
        RECT 12.480 1.470 12.490 1.644 ;
        RECT 12.490 1.470 12.496 1.640 ;
        RECT 12.390 1.500 12.400 1.734 ;
        RECT 12.400 1.490 12.410 1.724 ;
        RECT 12.410 1.480 12.420 1.714 ;
        RECT 12.220 1.670 12.230 2.514 ;
        RECT 12.230 1.660 12.240 2.524 ;
        RECT 12.240 1.650 12.250 2.534 ;
        RECT 12.250 1.640 12.260 2.544 ;
        RECT 12.260 1.630 12.270 2.554 ;
        RECT 12.270 1.620 12.280 2.564 ;
        RECT 12.280 1.610 12.290 2.574 ;
        RECT 12.290 1.600 12.300 2.584 ;
        RECT 12.300 1.590 12.310 2.594 ;
        RECT 12.310 1.580 12.320 2.604 ;
        RECT 12.320 1.570 12.330 2.614 ;
        RECT 12.330 1.560 12.340 2.624 ;
        RECT 12.340 1.550 12.350 2.634 ;
        RECT 12.350 1.540 12.360 2.644 ;
        RECT 12.360 1.530 12.370 2.654 ;
        RECT 12.370 1.520 12.380 2.664 ;
        RECT 12.380 1.510 12.390 2.674 ;
        RECT 12.190 2.315 12.200 2.485 ;
        RECT 12.200 2.315 12.210 2.495 ;
        RECT 12.210 2.315 12.220 2.505 ;
        RECT 11.070 2.315 11.080 2.549 ;
        RECT 11.080 2.315 11.090 2.539 ;
        RECT 11.090 2.315 11.100 2.529 ;
        RECT 11.100 2.315 11.110 2.519 ;
        RECT 11.110 2.315 11.120 2.509 ;
        RECT 11.120 2.315 11.130 2.499 ;
        RECT 11.130 2.315 11.140 2.489 ;
        RECT 11.140 2.315 11.146 2.485 ;
        RECT 10.975 2.410 10.985 2.644 ;
        RECT 10.985 2.400 10.995 2.634 ;
        RECT 10.995 2.390 11.005 2.624 ;
        RECT 11.005 2.380 11.015 2.614 ;
        RECT 11.015 2.370 11.025 2.604 ;
        RECT 11.025 2.360 11.035 2.594 ;
        RECT 11.035 2.350 11.045 2.584 ;
        RECT 11.045 2.340 11.055 2.574 ;
        RECT 11.055 2.330 11.065 2.564 ;
        RECT 11.065 2.320 11.071 2.560 ;
        RECT 10.900 2.485 10.910 2.655 ;
        RECT 10.910 2.475 10.920 2.655 ;
        RECT 10.920 2.465 10.930 2.655 ;
        RECT 10.930 2.455 10.940 2.655 ;
        RECT 10.940 2.445 10.950 2.655 ;
        RECT 10.950 2.435 10.960 2.655 ;
        RECT 10.960 2.425 10.970 2.655 ;
        RECT 10.970 2.415 10.976 2.655 ;
        RECT 9.685 2.485 9.695 2.735 ;
        RECT 9.695 2.485 9.705 2.725 ;
        RECT 9.705 2.485 9.715 2.715 ;
        RECT 9.715 2.485 9.725 2.705 ;
        RECT 9.725 2.485 9.735 2.695 ;
        RECT 9.735 2.485 9.745 2.685 ;
        RECT 9.745 2.485 9.755 2.675 ;
        RECT 9.755 2.485 9.765 2.665 ;
        RECT 9.765 2.485 9.775 2.655 ;
        RECT 9.590 2.580 9.600 2.830 ;
        RECT 9.600 2.570 9.610 2.820 ;
        RECT 9.610 2.560 9.620 2.810 ;
        RECT 9.620 2.550 9.630 2.800 ;
        RECT 9.630 2.540 9.640 2.790 ;
        RECT 9.640 2.530 9.650 2.780 ;
        RECT 9.650 2.520 9.660 2.770 ;
        RECT 9.660 2.510 9.670 2.760 ;
        RECT 9.670 2.500 9.680 2.750 ;
        RECT 9.680 2.490 9.686 2.744 ;
        RECT 9.500 2.670 9.510 2.840 ;
        RECT 9.510 2.660 9.520 2.840 ;
        RECT 9.520 2.650 9.530 2.840 ;
        RECT 9.530 2.640 9.540 2.840 ;
        RECT 9.540 2.630 9.550 2.840 ;
        RECT 9.550 2.620 9.560 2.840 ;
        RECT 9.560 2.610 9.570 2.840 ;
        RECT 9.570 2.600 9.580 2.840 ;
        RECT 9.580 2.590 9.590 2.840 ;
        RECT 10.520 2.940 10.950 3.110 ;
        RECT 11.300 2.665 12.040 2.835 ;
        RECT 11.870 2.665 12.040 3.190 ;
        RECT 14.830 1.325 15.000 1.830 ;
        RECT 14.830 1.660 15.265 1.830 ;
        RECT 15.095 1.660 15.265 3.190 ;
        RECT 11.870 3.020 15.265 3.190 ;
        RECT 11.225 2.665 11.235 2.899 ;
        RECT 11.235 2.665 11.245 2.889 ;
        RECT 11.245 2.665 11.255 2.879 ;
        RECT 11.255 2.665 11.265 2.869 ;
        RECT 11.265 2.665 11.275 2.859 ;
        RECT 11.275 2.665 11.285 2.849 ;
        RECT 11.285 2.665 11.295 2.839 ;
        RECT 11.295 2.665 11.301 2.835 ;
        RECT 11.025 2.865 11.035 3.099 ;
        RECT 11.035 2.855 11.045 3.089 ;
        RECT 11.045 2.845 11.055 3.079 ;
        RECT 11.055 2.835 11.065 3.069 ;
        RECT 11.065 2.825 11.075 3.059 ;
        RECT 11.075 2.815 11.085 3.049 ;
        RECT 11.085 2.805 11.095 3.039 ;
        RECT 11.095 2.795 11.105 3.029 ;
        RECT 11.105 2.785 11.115 3.019 ;
        RECT 11.115 2.775 11.125 3.009 ;
        RECT 11.125 2.765 11.135 2.999 ;
        RECT 11.135 2.755 11.145 2.989 ;
        RECT 11.145 2.745 11.155 2.979 ;
        RECT 11.155 2.735 11.165 2.969 ;
        RECT 11.165 2.725 11.175 2.959 ;
        RECT 11.175 2.715 11.185 2.949 ;
        RECT 11.185 2.705 11.195 2.939 ;
        RECT 11.195 2.695 11.205 2.929 ;
        RECT 11.205 2.685 11.215 2.919 ;
        RECT 11.215 2.675 11.225 2.909 ;
        RECT 10.950 2.940 10.960 3.110 ;
        RECT 10.960 2.930 10.970 3.110 ;
        RECT 10.970 2.920 10.980 3.110 ;
        RECT 10.980 2.910 10.990 3.110 ;
        RECT 10.990 2.900 11.000 3.110 ;
        RECT 11.000 2.890 11.010 3.110 ;
        RECT 11.010 2.880 11.020 3.110 ;
        RECT 11.020 2.870 11.026 3.110 ;
        RECT 15.795 1.465 15.965 1.765 ;
        RECT 16.470 1.115 16.645 1.635 ;
        RECT 15.795 1.465 16.645 1.635 ;
        RECT 16.475 1.115 16.645 2.340 ;
        RECT 16.405 1.115 16.705 1.285 ;
        RECT 16.475 2.170 17.105 2.340 ;
        RECT 16.015 0.765 16.185 1.285 ;
        RECT 15.885 1.115 16.185 1.285 ;
        RECT 16.015 0.765 17.095 0.935 ;
        RECT 16.925 0.765 17.095 1.285 ;
        RECT 16.925 1.115 17.225 1.285 ;
        RECT 13.665 1.075 13.835 1.415 ;
        RECT 12.875 1.075 13.835 1.245 ;
        RECT 13.665 1.245 14.650 1.415 ;
        RECT 14.480 0.860 14.650 2.460 ;
        RECT 12.780 2.290 14.650 2.460 ;
        RECT 14.480 0.860 14.725 1.160 ;
        RECT 14.480 2.050 14.790 2.220 ;
        RECT 14.480 0.860 15.095 1.030 ;
        RECT 15.375 1.065 15.615 1.235 ;
        RECT 15.445 1.065 15.615 2.115 ;
        RECT 15.445 1.945 16.240 2.115 ;
        RECT 16.070 1.945 16.240 2.720 ;
        RECT 17.625 1.510 17.795 2.720 ;
        RECT 16.070 2.550 17.795 2.720 ;
        RECT 17.625 1.510 17.870 1.810 ;
        RECT 15.300 1.000 15.310 1.234 ;
        RECT 15.310 1.010 15.320 1.234 ;
        RECT 15.320 1.020 15.330 1.234 ;
        RECT 15.330 1.030 15.340 1.234 ;
        RECT 15.340 1.040 15.350 1.234 ;
        RECT 15.350 1.050 15.360 1.234 ;
        RECT 15.360 1.060 15.370 1.234 ;
        RECT 15.370 1.065 15.376 1.235 ;
        RECT 15.170 0.870 15.180 1.104 ;
        RECT 15.180 0.880 15.190 1.114 ;
        RECT 15.190 0.890 15.200 1.124 ;
        RECT 15.200 0.900 15.210 1.134 ;
        RECT 15.210 0.910 15.220 1.144 ;
        RECT 15.220 0.920 15.230 1.154 ;
        RECT 15.230 0.930 15.240 1.164 ;
        RECT 15.240 0.940 15.250 1.174 ;
        RECT 15.250 0.950 15.260 1.184 ;
        RECT 15.260 0.960 15.270 1.194 ;
        RECT 15.270 0.970 15.280 1.204 ;
        RECT 15.280 0.980 15.290 1.214 ;
        RECT 15.290 0.990 15.300 1.224 ;
        RECT 15.095 0.860 15.105 1.030 ;
        RECT 15.105 0.860 15.115 1.040 ;
        RECT 15.115 0.860 15.125 1.050 ;
        RECT 15.125 0.860 15.135 1.060 ;
        RECT 15.135 0.860 15.145 1.070 ;
        RECT 15.145 0.860 15.155 1.080 ;
        RECT 15.155 0.860 15.165 1.090 ;
        RECT 15.165 0.860 15.171 1.100 ;
  END 
END FFSDSRHQHD2XHT

MACRO FFSDSRHQHD1XHT
  CLASS  CORE ;
  FOREIGN FFSDSRHQHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.170 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.815 0.720 15.070 2.960 ;
        RECT 14.765 1.980 15.070 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 1.290 1.605 1.540 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.060 1.435 7.510 2.045 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.520 1.735 0.690 2.100 ;
        RECT 0.815 1.930 1.230 2.360 ;
        RECT 1.400 1.735 1.570 2.100 ;
        RECT 0.520 1.930 1.570 2.100 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.995 ;
        RECT 2.435 -0.300 2.735 0.785 ;
        RECT 3.350 -0.300 3.650 0.945 ;
        RECT 7.135 -0.300 7.435 1.130 ;
        RECT 10.390 -0.300 10.560 1.220 ;
        RECT 12.220 -0.300 12.520 0.795 ;
        RECT 14.290 -0.300 14.460 1.345 ;
        RECT 0.000 -0.300 15.170 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.825 1.550 3.275 2.015 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.145 1.395 2.535 2.015 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 13.545 1.540 14.170 1.960 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.905 0.895 3.990 ;
        RECT 2.490 2.895 3.470 3.990 ;
        RECT 4.395 2.895 4.695 3.990 ;
        RECT 7.310 3.025 8.290 3.990 ;
        RECT 10.200 3.025 10.500 3.990 ;
        RECT 12.325 2.315 12.625 3.990 ;
        RECT 14.180 2.975 14.480 3.990 ;
        RECT 0.000 3.390 15.170 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.170 0.340 2.470 ;
        RECT 0.105 0.825 0.275 2.470 ;
        RECT 0.170 2.170 0.340 2.725 ;
        RECT 0.105 0.825 0.405 0.995 ;
        RECT 0.170 2.555 1.305 2.725 ;
        RECT 1.135 2.555 1.305 3.210 ;
        RECT 1.135 3.040 1.995 3.210 ;
        RECT 2.780 1.125 3.770 1.295 ;
        RECT 3.600 1.125 3.770 2.365 ;
        RECT 2.825 2.195 3.770 2.365 ;
        RECT 4.860 0.975 5.430 1.145 ;
        RECT 5.260 0.975 5.430 2.295 ;
        RECT 1.580 0.725 1.750 1.055 ;
        RECT 1.580 0.885 1.960 1.055 ;
        RECT 1.790 0.885 1.960 2.715 ;
        RECT 1.580 2.415 1.960 2.715 ;
        RECT 1.580 2.545 5.780 2.715 ;
        RECT 5.610 0.895 5.780 2.760 ;
        RECT 5.480 2.545 5.780 2.760 ;
        RECT 7.750 0.960 7.920 2.125 ;
        RECT 7.655 0.960 7.955 1.130 ;
        RECT 7.750 1.675 7.985 2.125 ;
        RECT 7.750 1.675 8.495 1.845 ;
        RECT 6.310 0.895 6.480 2.475 ;
        RECT 8.705 1.615 8.875 2.475 ;
        RECT 6.310 2.305 8.875 2.475 ;
        RECT 8.705 1.615 9.180 1.785 ;
        RECT 8.165 0.970 8.465 1.380 ;
        RECT 9.180 0.965 9.350 1.380 ;
        RECT 8.165 1.205 9.350 1.380 ;
        RECT 9.180 0.965 9.860 1.135 ;
        RECT 7.795 0.480 8.095 0.730 ;
        RECT 8.695 0.560 8.995 1.015 ;
        RECT 9.525 1.580 9.695 2.215 ;
        RECT 9.055 2.045 9.695 2.215 ;
        RECT 7.795 0.560 10.210 0.730 ;
        RECT 10.040 0.560 10.210 1.750 ;
        RECT 9.525 1.580 10.755 1.750 ;
        RECT 3.950 0.545 4.155 2.365 ;
        RECT 5.960 0.545 6.130 3.160 ;
        RECT 3.950 0.545 6.725 0.715 ;
        RECT 5.960 2.655 9.525 2.825 ;
        RECT 9.930 2.325 10.810 2.495 ;
        RECT 10.880 2.325 10.885 2.565 ;
        RECT 10.955 2.395 11.635 2.565 ;
        RECT 11.465 2.395 11.635 2.770 ;
        RECT 10.885 2.335 10.895 2.565 ;
        RECT 10.895 2.345 10.905 2.565 ;
        RECT 10.905 2.355 10.915 2.565 ;
        RECT 10.915 2.365 10.925 2.565 ;
        RECT 10.925 2.375 10.935 2.565 ;
        RECT 10.935 2.385 10.945 2.565 ;
        RECT 10.945 2.395 10.955 2.565 ;
        RECT 10.810 2.325 10.820 2.495 ;
        RECT 10.820 2.325 10.830 2.505 ;
        RECT 10.830 2.325 10.840 2.515 ;
        RECT 10.840 2.325 10.850 2.525 ;
        RECT 10.850 2.325 10.860 2.535 ;
        RECT 10.860 2.325 10.870 2.545 ;
        RECT 10.870 2.325 10.880 2.555 ;
        RECT 9.855 2.325 9.865 2.559 ;
        RECT 9.865 2.325 9.875 2.549 ;
        RECT 9.875 2.325 9.885 2.539 ;
        RECT 9.885 2.325 9.895 2.529 ;
        RECT 9.895 2.325 9.905 2.519 ;
        RECT 9.905 2.325 9.915 2.509 ;
        RECT 9.915 2.325 9.925 2.499 ;
        RECT 9.925 2.325 9.931 2.495 ;
        RECT 9.600 2.580 9.610 2.814 ;
        RECT 9.610 2.570 9.620 2.804 ;
        RECT 9.620 2.560 9.630 2.794 ;
        RECT 9.630 2.550 9.640 2.784 ;
        RECT 9.640 2.540 9.650 2.774 ;
        RECT 9.650 2.530 9.660 2.764 ;
        RECT 9.660 2.520 9.670 2.754 ;
        RECT 9.670 2.510 9.680 2.744 ;
        RECT 9.680 2.500 9.690 2.734 ;
        RECT 9.690 2.490 9.700 2.724 ;
        RECT 9.700 2.480 9.710 2.714 ;
        RECT 9.710 2.470 9.720 2.704 ;
        RECT 9.720 2.460 9.730 2.694 ;
        RECT 9.730 2.450 9.740 2.684 ;
        RECT 9.740 2.440 9.750 2.674 ;
        RECT 9.750 2.430 9.760 2.664 ;
        RECT 9.760 2.420 9.770 2.654 ;
        RECT 9.770 2.410 9.780 2.644 ;
        RECT 9.780 2.400 9.790 2.634 ;
        RECT 9.790 2.390 9.800 2.624 ;
        RECT 9.800 2.380 9.810 2.614 ;
        RECT 9.810 2.370 9.820 2.604 ;
        RECT 9.820 2.360 9.830 2.594 ;
        RECT 9.830 2.350 9.840 2.584 ;
        RECT 9.840 2.340 9.850 2.574 ;
        RECT 9.850 2.330 9.856 2.570 ;
        RECT 9.525 2.655 9.535 2.825 ;
        RECT 9.535 2.645 9.545 2.825 ;
        RECT 9.545 2.635 9.555 2.825 ;
        RECT 9.555 2.625 9.565 2.825 ;
        RECT 9.565 2.615 9.575 2.825 ;
        RECT 9.575 2.605 9.585 2.825 ;
        RECT 9.585 2.595 9.595 2.825 ;
        RECT 9.595 2.585 9.601 2.825 ;
        RECT 9.275 3.025 9.670 3.195 ;
        RECT 10.095 2.675 10.635 2.845 ;
        RECT 10.705 2.675 10.730 2.915 ;
        RECT 10.800 2.745 11.240 2.915 ;
        RECT 11.070 2.745 11.240 3.120 ;
        RECT 11.530 1.270 11.830 1.440 ;
        RECT 11.660 1.270 11.830 1.825 ;
        RECT 11.660 1.655 12.030 1.825 ;
        RECT 11.860 1.655 12.030 3.120 ;
        RECT 11.860 2.815 12.130 3.120 ;
        RECT 11.070 2.950 12.130 3.120 ;
        RECT 10.730 2.685 10.740 2.915 ;
        RECT 10.740 2.695 10.750 2.915 ;
        RECT 10.750 2.705 10.760 2.915 ;
        RECT 10.760 2.715 10.770 2.915 ;
        RECT 10.770 2.725 10.780 2.915 ;
        RECT 10.780 2.735 10.790 2.915 ;
        RECT 10.790 2.745 10.800 2.915 ;
        RECT 10.635 2.675 10.645 2.845 ;
        RECT 10.645 2.675 10.655 2.855 ;
        RECT 10.655 2.675 10.665 2.865 ;
        RECT 10.665 2.675 10.675 2.875 ;
        RECT 10.675 2.675 10.685 2.885 ;
        RECT 10.685 2.675 10.695 2.895 ;
        RECT 10.695 2.675 10.705 2.905 ;
        RECT 10.020 2.675 10.030 2.909 ;
        RECT 10.030 2.675 10.040 2.899 ;
        RECT 10.040 2.675 10.050 2.889 ;
        RECT 10.050 2.675 10.060 2.879 ;
        RECT 10.060 2.675 10.070 2.869 ;
        RECT 10.070 2.675 10.080 2.859 ;
        RECT 10.080 2.675 10.090 2.849 ;
        RECT 10.090 2.675 10.096 2.845 ;
        RECT 9.745 2.950 9.755 3.184 ;
        RECT 9.755 2.940 9.765 3.174 ;
        RECT 9.765 2.930 9.775 3.164 ;
        RECT 9.775 2.920 9.785 3.154 ;
        RECT 9.785 2.910 9.795 3.144 ;
        RECT 9.795 2.900 9.805 3.134 ;
        RECT 9.805 2.890 9.815 3.124 ;
        RECT 9.815 2.880 9.825 3.114 ;
        RECT 9.825 2.870 9.835 3.104 ;
        RECT 9.835 2.860 9.845 3.094 ;
        RECT 9.845 2.850 9.855 3.084 ;
        RECT 9.855 2.840 9.865 3.074 ;
        RECT 9.865 2.830 9.875 3.064 ;
        RECT 9.875 2.820 9.885 3.054 ;
        RECT 9.885 2.810 9.895 3.044 ;
        RECT 9.895 2.800 9.905 3.034 ;
        RECT 9.905 2.790 9.915 3.024 ;
        RECT 9.915 2.780 9.925 3.014 ;
        RECT 9.925 2.770 9.935 3.004 ;
        RECT 9.935 2.760 9.945 2.994 ;
        RECT 9.945 2.750 9.955 2.984 ;
        RECT 9.955 2.740 9.965 2.974 ;
        RECT 9.965 2.730 9.975 2.964 ;
        RECT 9.975 2.720 9.985 2.954 ;
        RECT 9.985 2.710 9.995 2.944 ;
        RECT 9.995 2.700 10.005 2.934 ;
        RECT 10.005 2.690 10.015 2.924 ;
        RECT 10.015 2.680 10.021 2.920 ;
        RECT 9.670 3.025 9.680 3.195 ;
        RECT 9.680 3.015 9.690 3.195 ;
        RECT 9.690 3.005 9.700 3.195 ;
        RECT 9.700 2.995 9.710 3.195 ;
        RECT 9.710 2.985 9.720 3.195 ;
        RECT 9.720 2.975 9.730 3.195 ;
        RECT 9.730 2.965 9.740 3.195 ;
        RECT 9.740 2.955 9.746 3.195 ;
        RECT 12.560 1.460 12.730 1.760 ;
        RECT 13.170 1.110 13.345 1.630 ;
        RECT 12.560 1.460 13.345 1.630 ;
        RECT 13.175 1.110 13.345 2.335 ;
        RECT 13.170 1.110 13.470 1.280 ;
        RECT 13.175 2.165 13.870 2.335 ;
        RECT 12.780 0.760 12.950 1.280 ;
        RECT 12.650 1.110 12.950 1.280 ;
        RECT 12.780 0.760 13.860 0.930 ;
        RECT 13.690 0.760 13.860 1.280 ;
        RECT 13.690 1.110 13.990 1.280 ;
        RECT 11.120 0.900 11.290 2.215 ;
        RECT 11.120 2.045 11.420 2.215 ;
        RECT 11.120 0.900 11.905 1.070 ;
        RECT 12.140 1.060 12.380 1.230 ;
        RECT 12.210 1.060 12.380 2.110 ;
        RECT 12.210 1.940 12.975 2.110 ;
        RECT 12.805 1.940 12.975 2.715 ;
        RECT 14.390 1.540 14.560 2.715 ;
        RECT 12.805 2.545 14.560 2.715 ;
        RECT 14.390 1.540 14.635 1.840 ;
        RECT 12.065 0.995 12.075 1.229 ;
        RECT 12.075 1.005 12.085 1.229 ;
        RECT 12.085 1.015 12.095 1.229 ;
        RECT 12.095 1.025 12.105 1.229 ;
        RECT 12.105 1.035 12.115 1.229 ;
        RECT 12.115 1.045 12.125 1.229 ;
        RECT 12.125 1.055 12.135 1.229 ;
        RECT 12.135 1.060 12.141 1.230 ;
        RECT 11.980 0.910 11.990 1.144 ;
        RECT 11.990 0.920 12.000 1.154 ;
        RECT 12.000 0.930 12.010 1.164 ;
        RECT 12.010 0.940 12.020 1.174 ;
        RECT 12.020 0.950 12.030 1.184 ;
        RECT 12.030 0.960 12.040 1.194 ;
        RECT 12.040 0.970 12.050 1.204 ;
        RECT 12.050 0.980 12.060 1.214 ;
        RECT 12.060 0.985 12.066 1.225 ;
        RECT 11.905 0.900 11.915 1.070 ;
        RECT 11.915 0.900 11.925 1.080 ;
        RECT 11.925 0.900 11.935 1.090 ;
        RECT 11.935 0.900 11.945 1.100 ;
        RECT 11.945 0.900 11.955 1.110 ;
        RECT 11.955 0.900 11.965 1.120 ;
        RECT 11.965 0.900 11.975 1.130 ;
        RECT 11.975 0.900 11.981 1.140 ;
  END 
END FFSDSRHQHD1XHT

MACRO FFSDSRHDLXHT
  CLASS  CORE ;
  FOREIGN FFSDSRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.760 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.410 0.995 14.580 2.845 ;
        RECT 14.410 2.490 14.660 2.845 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.145 0.920 13.680 1.230 ;
        RECT 13.510 0.920 13.680 2.215 ;
        RECT 13.245 2.045 13.680 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.835 1.290 1.605 1.540 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.980 1.740 6.525 2.055 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.520 1.735 0.690 2.050 ;
        RECT 0.815 1.880 1.230 2.360 ;
        RECT 1.400 1.735 1.570 2.050 ;
        RECT 0.520 1.880 1.570 2.050 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.090 ;
        RECT 2.525 -0.300 2.825 0.785 ;
        RECT 3.330 -0.300 3.630 0.745 ;
        RECT 6.020 -0.300 6.320 0.460 ;
        RECT 8.950 -0.300 9.120 0.860 ;
        RECT 10.790 -0.300 11.090 0.770 ;
        RECT 12.825 -0.300 13.125 0.715 ;
        RECT 13.860 -0.300 14.030 1.295 ;
        RECT 0.000 -0.300 14.760 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.965 1.550 3.370 2.015 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.290 1.550 2.775 2.015 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 12.315 1.355 12.680 1.950 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.905 0.895 3.990 ;
        RECT 2.540 2.935 3.520 3.990 ;
        RECT 6.190 2.995 7.170 3.990 ;
        RECT 8.835 2.995 9.135 3.990 ;
        RECT 10.860 2.315 11.160 3.990 ;
        RECT 12.735 2.930 13.035 3.990 ;
        RECT 13.795 2.790 14.095 3.990 ;
        RECT 0.000 3.390 14.760 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.920 0.275 2.725 ;
        RECT 0.105 2.290 0.340 2.725 ;
        RECT 0.105 0.920 0.405 1.090 ;
        RECT 0.105 2.555 1.305 2.725 ;
        RECT 1.135 2.555 1.305 3.075 ;
        RECT 1.135 2.905 1.995 3.075 ;
        RECT 2.825 1.125 3.795 1.295 ;
        RECT 3.625 1.125 3.795 2.365 ;
        RECT 2.825 2.195 3.795 2.365 ;
        RECT 1.575 0.920 1.985 1.090 ;
        RECT 1.815 0.920 1.985 2.715 ;
        RECT 1.580 2.230 1.985 2.715 ;
        RECT 1.580 2.545 3.775 2.715 ;
        RECT 3.710 2.610 4.660 2.725 ;
        RECT 3.720 2.610 4.660 2.735 ;
        RECT 3.730 2.610 4.660 2.745 ;
        RECT 3.740 2.610 4.660 2.755 ;
        RECT 3.750 2.610 4.660 2.765 ;
        RECT 3.760 2.610 4.660 2.775 ;
        RECT 3.765 2.545 3.775 2.780 ;
        RECT 1.580 2.555 3.785 2.715 ;
        RECT 1.580 2.565 3.795 2.715 ;
        RECT 1.580 2.575 3.805 2.715 ;
        RECT 1.580 2.585 3.815 2.715 ;
        RECT 1.580 2.595 3.825 2.715 ;
        RECT 3.765 2.610 4.660 2.779 ;
        RECT 1.580 2.605 3.835 2.715 ;
        RECT 4.490 0.895 4.660 2.780 ;
        RECT 3.835 2.610 4.660 2.780 ;
        RECT 6.725 0.960 6.895 2.115 ;
        RECT 6.635 0.960 6.935 1.130 ;
        RECT 6.725 1.500 7.520 1.670 ;
        RECT 5.190 0.895 5.360 2.465 ;
        RECT 5.190 0.895 5.390 1.195 ;
        RECT 7.700 1.680 7.870 2.465 ;
        RECT 5.190 2.295 7.870 2.465 ;
        RECT 7.935 1.550 8.105 1.850 ;
        RECT 7.700 1.680 8.105 1.850 ;
        RECT 7.145 0.960 7.445 1.230 ;
        RECT 7.145 1.060 8.420 1.230 ;
        RECT 8.250 1.060 8.420 1.360 ;
        RECT 5.845 1.330 6.260 1.500 ;
        RECT 8.050 2.045 8.175 2.215 ;
        RECT 8.285 1.580 8.350 2.215 ;
        RECT 6.610 0.560 8.770 0.730 ;
        RECT 8.600 0.560 8.770 1.750 ;
        RECT 8.455 1.580 9.340 1.750 ;
        RECT 8.350 1.580 8.360 2.104 ;
        RECT 8.360 1.580 8.370 2.094 ;
        RECT 8.370 1.580 8.380 2.084 ;
        RECT 8.380 1.580 8.390 2.074 ;
        RECT 8.390 1.580 8.400 2.064 ;
        RECT 8.400 1.580 8.410 2.054 ;
        RECT 8.410 1.580 8.420 2.044 ;
        RECT 8.420 1.580 8.430 2.034 ;
        RECT 8.430 1.580 8.440 2.024 ;
        RECT 8.440 1.580 8.450 2.014 ;
        RECT 8.450 1.580 8.456 2.010 ;
        RECT 8.175 2.045 8.185 2.215 ;
        RECT 8.185 2.035 8.195 2.215 ;
        RECT 8.195 2.025 8.205 2.215 ;
        RECT 8.205 2.015 8.215 2.215 ;
        RECT 8.215 2.005 8.225 2.215 ;
        RECT 8.225 1.995 8.235 2.215 ;
        RECT 8.235 1.985 8.245 2.215 ;
        RECT 8.245 1.975 8.255 2.215 ;
        RECT 8.255 1.965 8.265 2.215 ;
        RECT 8.265 1.955 8.275 2.215 ;
        RECT 8.275 1.945 8.285 2.215 ;
        RECT 6.530 0.560 6.540 0.800 ;
        RECT 6.540 0.560 6.550 0.790 ;
        RECT 6.550 0.560 6.560 0.780 ;
        RECT 6.560 0.560 6.570 0.770 ;
        RECT 6.570 0.560 6.580 0.760 ;
        RECT 6.580 0.560 6.590 0.750 ;
        RECT 6.590 0.560 6.600 0.740 ;
        RECT 6.600 0.560 6.610 0.730 ;
        RECT 6.430 0.660 6.440 0.900 ;
        RECT 6.440 0.650 6.450 0.890 ;
        RECT 6.450 0.640 6.460 0.880 ;
        RECT 6.460 0.630 6.470 0.870 ;
        RECT 6.470 0.620 6.480 0.860 ;
        RECT 6.480 0.610 6.490 0.850 ;
        RECT 6.490 0.600 6.500 0.840 ;
        RECT 6.500 0.590 6.510 0.830 ;
        RECT 6.510 0.580 6.520 0.820 ;
        RECT 6.520 0.570 6.530 0.810 ;
        RECT 6.260 0.830 6.270 1.500 ;
        RECT 6.270 0.820 6.280 1.500 ;
        RECT 6.280 0.810 6.290 1.500 ;
        RECT 6.290 0.800 6.300 1.500 ;
        RECT 6.300 0.790 6.310 1.500 ;
        RECT 6.310 0.780 6.320 1.500 ;
        RECT 6.320 0.770 6.330 1.500 ;
        RECT 6.330 0.760 6.340 1.500 ;
        RECT 6.340 0.750 6.350 1.500 ;
        RECT 6.350 0.740 6.360 1.500 ;
        RECT 6.360 0.730 6.370 1.500 ;
        RECT 6.370 0.720 6.380 1.500 ;
        RECT 6.380 0.710 6.390 1.500 ;
        RECT 6.390 0.700 6.400 1.500 ;
        RECT 6.400 0.690 6.410 1.500 ;
        RECT 6.410 0.680 6.420 1.500 ;
        RECT 6.420 0.670 6.430 1.500 ;
        RECT 3.975 0.545 4.145 2.430 ;
        RECT 4.840 0.545 5.010 2.835 ;
        RECT 3.975 0.545 5.665 0.715 ;
        RECT 4.840 2.645 8.180 2.815 ;
        RECT 8.605 2.295 9.365 2.465 ;
        RECT 9.540 2.395 10.080 2.565 ;
        RECT 9.910 2.395 10.080 2.695 ;
        RECT 9.465 2.330 9.475 2.564 ;
        RECT 9.475 2.340 9.485 2.564 ;
        RECT 9.485 2.350 9.495 2.564 ;
        RECT 9.495 2.360 9.505 2.564 ;
        RECT 9.505 2.370 9.515 2.564 ;
        RECT 9.515 2.380 9.525 2.564 ;
        RECT 9.525 2.390 9.535 2.564 ;
        RECT 9.535 2.395 9.541 2.565 ;
        RECT 9.440 2.305 9.450 2.539 ;
        RECT 9.450 2.315 9.460 2.549 ;
        RECT 9.460 2.320 9.466 2.560 ;
        RECT 9.365 2.295 9.375 2.465 ;
        RECT 9.375 2.295 9.385 2.475 ;
        RECT 9.385 2.295 9.395 2.485 ;
        RECT 9.395 2.295 9.405 2.495 ;
        RECT 9.405 2.295 9.415 2.505 ;
        RECT 9.415 2.295 9.425 2.515 ;
        RECT 9.425 2.295 9.435 2.525 ;
        RECT 9.435 2.295 9.441 2.535 ;
        RECT 8.530 2.295 8.540 2.529 ;
        RECT 8.540 2.295 8.550 2.519 ;
        RECT 8.550 2.295 8.560 2.509 ;
        RECT 8.560 2.295 8.570 2.499 ;
        RECT 8.570 2.295 8.580 2.489 ;
        RECT 8.580 2.295 8.590 2.479 ;
        RECT 8.590 2.295 8.600 2.469 ;
        RECT 8.600 2.295 8.606 2.465 ;
        RECT 8.255 2.570 8.265 2.804 ;
        RECT 8.265 2.560 8.275 2.794 ;
        RECT 8.275 2.550 8.285 2.784 ;
        RECT 8.285 2.540 8.295 2.774 ;
        RECT 8.295 2.530 8.305 2.764 ;
        RECT 8.305 2.520 8.315 2.754 ;
        RECT 8.315 2.510 8.325 2.744 ;
        RECT 8.325 2.500 8.335 2.734 ;
        RECT 8.335 2.490 8.345 2.724 ;
        RECT 8.345 2.480 8.355 2.714 ;
        RECT 8.355 2.470 8.365 2.704 ;
        RECT 8.365 2.460 8.375 2.694 ;
        RECT 8.375 2.450 8.385 2.684 ;
        RECT 8.385 2.440 8.395 2.674 ;
        RECT 8.395 2.430 8.405 2.664 ;
        RECT 8.405 2.420 8.415 2.654 ;
        RECT 8.415 2.410 8.425 2.644 ;
        RECT 8.425 2.400 8.435 2.634 ;
        RECT 8.435 2.390 8.445 2.624 ;
        RECT 8.445 2.380 8.455 2.614 ;
        RECT 8.455 2.370 8.465 2.604 ;
        RECT 8.465 2.360 8.475 2.594 ;
        RECT 8.475 2.350 8.485 2.584 ;
        RECT 8.485 2.340 8.495 2.574 ;
        RECT 8.495 2.330 8.505 2.564 ;
        RECT 8.505 2.320 8.515 2.554 ;
        RECT 8.515 2.310 8.525 2.544 ;
        RECT 8.525 2.300 8.531 2.540 ;
        RECT 8.180 2.645 8.190 2.815 ;
        RECT 8.190 2.635 8.200 2.815 ;
        RECT 8.200 2.625 8.210 2.815 ;
        RECT 8.210 2.615 8.220 2.815 ;
        RECT 8.220 2.605 8.230 2.815 ;
        RECT 8.230 2.595 8.240 2.815 ;
        RECT 8.240 2.585 8.250 2.815 ;
        RECT 8.250 2.575 8.256 2.815 ;
        RECT 10.240 1.655 10.430 1.825 ;
        RECT 7.500 2.995 7.800 3.210 ;
        RECT 7.500 2.995 8.485 3.165 ;
        RECT 8.755 2.645 9.210 2.815 ;
        RECT 9.495 2.745 9.665 3.045 ;
        RECT 9.385 2.745 9.665 2.915 ;
        RECT 10.110 1.270 10.410 1.440 ;
        RECT 10.240 1.270 10.410 1.825 ;
        RECT 10.260 1.655 10.430 3.045 ;
        RECT 9.495 2.875 10.430 3.045 ;
        RECT 9.310 2.680 9.320 2.914 ;
        RECT 9.320 2.690 9.330 2.914 ;
        RECT 9.330 2.700 9.340 2.914 ;
        RECT 9.340 2.710 9.350 2.914 ;
        RECT 9.350 2.720 9.360 2.914 ;
        RECT 9.360 2.730 9.370 2.914 ;
        RECT 9.370 2.740 9.380 2.914 ;
        RECT 9.380 2.745 9.386 2.915 ;
        RECT 9.285 2.655 9.295 2.889 ;
        RECT 9.295 2.665 9.305 2.899 ;
        RECT 9.305 2.670 9.311 2.910 ;
        RECT 9.210 2.645 9.220 2.815 ;
        RECT 9.220 2.645 9.230 2.825 ;
        RECT 9.230 2.645 9.240 2.835 ;
        RECT 9.240 2.645 9.250 2.845 ;
        RECT 9.250 2.645 9.260 2.855 ;
        RECT 9.260 2.645 9.270 2.865 ;
        RECT 9.270 2.645 9.280 2.875 ;
        RECT 9.280 2.645 9.286 2.885 ;
        RECT 8.680 2.645 8.690 2.879 ;
        RECT 8.690 2.645 8.700 2.869 ;
        RECT 8.700 2.645 8.710 2.859 ;
        RECT 8.710 2.645 8.720 2.849 ;
        RECT 8.720 2.645 8.730 2.839 ;
        RECT 8.730 2.645 8.740 2.829 ;
        RECT 8.740 2.645 8.750 2.819 ;
        RECT 8.750 2.645 8.756 2.815 ;
        RECT 8.655 2.670 8.665 2.904 ;
        RECT 8.665 2.660 8.675 2.894 ;
        RECT 8.675 2.650 8.681 2.890 ;
        RECT 8.485 2.840 8.495 3.164 ;
        RECT 8.495 2.830 8.505 3.164 ;
        RECT 8.505 2.820 8.515 3.164 ;
        RECT 8.515 2.810 8.525 3.164 ;
        RECT 8.525 2.800 8.535 3.164 ;
        RECT 8.535 2.790 8.545 3.164 ;
        RECT 8.545 2.780 8.555 3.164 ;
        RECT 8.555 2.770 8.565 3.164 ;
        RECT 8.565 2.760 8.575 3.164 ;
        RECT 8.575 2.750 8.585 3.164 ;
        RECT 8.585 2.740 8.595 3.164 ;
        RECT 8.595 2.730 8.605 3.164 ;
        RECT 8.605 2.720 8.615 3.164 ;
        RECT 8.615 2.710 8.625 3.164 ;
        RECT 8.625 2.700 8.635 3.164 ;
        RECT 8.635 2.690 8.645 3.164 ;
        RECT 8.645 2.680 8.655 3.164 ;
        RECT 11.295 0.640 11.465 1.280 ;
        RECT 11.165 1.110 11.465 1.280 ;
        RECT 11.295 0.640 12.575 0.810 ;
        RECT 11.120 1.460 11.290 1.760 ;
        RECT 11.745 1.110 12.045 1.630 ;
        RECT 11.120 1.460 12.045 1.630 ;
        RECT 11.875 1.110 12.045 2.345 ;
        RECT 12.895 1.475 13.065 2.345 ;
        RECT 11.875 2.175 13.065 2.345 ;
        RECT 12.895 1.475 13.330 1.775 ;
        RECT 9.705 0.900 9.875 2.215 ;
        RECT 9.705 2.045 10.035 2.215 ;
        RECT 9.705 0.900 10.490 1.070 ;
        RECT 10.725 1.060 10.865 2.110 ;
        RECT 10.725 1.940 11.550 2.110 ;
        RECT 11.380 1.940 11.550 2.750 ;
        RECT 11.975 2.580 12.275 2.855 ;
        RECT 13.390 2.440 13.560 2.750 ;
        RECT 11.380 2.580 13.560 2.750 ;
        RECT 13.390 2.440 14.160 2.610 ;
        RECT 13.990 1.520 14.160 2.610 ;
        RECT 13.990 1.520 14.230 1.820 ;
        RECT 10.695 1.040 10.705 2.110 ;
        RECT 10.705 1.050 10.715 2.110 ;
        RECT 10.715 1.060 10.725 2.110 ;
        RECT 10.650 0.995 10.660 1.229 ;
        RECT 10.660 1.005 10.670 1.229 ;
        RECT 10.670 1.015 10.680 1.229 ;
        RECT 10.680 1.025 10.690 1.229 ;
        RECT 10.690 1.030 10.696 1.230 ;
        RECT 10.565 0.910 10.575 1.144 ;
        RECT 10.575 0.920 10.585 1.154 ;
        RECT 10.585 0.930 10.595 1.164 ;
        RECT 10.595 0.940 10.605 1.174 ;
        RECT 10.605 0.950 10.615 1.184 ;
        RECT 10.615 0.960 10.625 1.194 ;
        RECT 10.625 0.970 10.635 1.204 ;
        RECT 10.635 0.980 10.645 1.214 ;
        RECT 10.645 0.985 10.651 1.225 ;
        RECT 10.490 0.900 10.500 1.070 ;
        RECT 10.500 0.900 10.510 1.080 ;
        RECT 10.510 0.900 10.520 1.090 ;
        RECT 10.520 0.900 10.530 1.100 ;
        RECT 10.530 0.900 10.540 1.110 ;
        RECT 10.540 0.900 10.550 1.120 ;
        RECT 10.550 0.900 10.560 1.130 ;
        RECT 10.560 0.900 10.566 1.140 ;
  END 
END FFSDSRHDLXHT

MACRO FFSDSRHD2XHT
  CLASS  CORE ;
  FOREIGN FFSDSRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.400 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 15.325 1.300 15.795 1.470 ;
        RECT 15.325 0.785 15.625 1.470 ;
        RECT 15.325 2.045 15.625 2.895 ;
        RECT 15.625 1.300 15.795 2.360 ;
        RECT 15.325 2.045 15.795 2.360 ;
        RECT 15.325 2.150 15.970 2.360 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.285 0.785 14.585 1.295 ;
        RECT 14.285 1.125 14.785 1.295 ;
        RECT 14.615 1.125 14.785 2.385 ;
        RECT 14.285 2.130 14.785 2.385 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.870 1.240 1.605 1.540 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.760 1.425 6.430 1.955 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.520 1.735 0.690 2.100 ;
        RECT 0.815 1.930 1.290 2.365 ;
        RECT 1.400 1.735 1.570 2.100 ;
        RECT 0.520 1.930 1.570 2.100 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.995 ;
        RECT 2.435 -0.300 2.735 0.745 ;
        RECT 3.405 -0.300 3.705 0.715 ;
        RECT 6.000 -0.300 6.300 0.990 ;
        RECT 9.025 -0.300 9.195 1.020 ;
        RECT 11.035 -0.300 11.335 0.815 ;
        RECT 13.290 -0.300 13.930 1.055 ;
        RECT 14.805 -0.300 15.105 0.715 ;
        RECT 15.845 -0.300 16.145 1.055 ;
        RECT 0.000 -0.300 16.400 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.970 1.475 3.320 2.015 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.290 1.500 2.775 2.015 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 13.350 1.325 13.520 1.775 ;
        RECT 13.350 1.325 13.965 1.545 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.995 0.895 3.990 ;
        RECT 2.515 2.895 3.495 3.990 ;
        RECT 6.165 2.995 7.145 3.990 ;
        RECT 8.945 2.995 9.245 3.990 ;
        RECT 11.020 2.385 11.190 3.990 ;
        RECT 12.795 3.015 13.095 3.990 ;
        RECT 13.765 2.975 14.065 3.990 ;
        RECT 14.805 2.975 15.105 3.990 ;
        RECT 15.845 2.635 16.145 3.990 ;
        RECT 0.000 3.390 16.400 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.825 0.275 2.735 ;
        RECT 0.105 2.290 0.340 2.735 ;
        RECT 0.105 0.825 0.405 0.995 ;
        RECT 0.105 2.565 1.340 2.735 ;
        RECT 1.170 2.565 1.340 3.210 ;
        RECT 1.170 3.040 1.995 3.210 ;
        RECT 2.825 1.125 3.675 1.295 ;
        RECT 3.505 1.125 3.675 2.365 ;
        RECT 2.825 2.195 3.675 2.365 ;
        RECT 3.505 1.525 3.795 1.825 ;
        RECT 1.515 0.790 1.985 0.960 ;
        RECT 1.700 2.365 1.985 2.715 ;
        RECT 1.815 0.790 1.985 2.715 ;
        RECT 1.580 2.370 1.985 2.715 ;
        RECT 1.580 2.545 4.600 2.715 ;
        RECT 4.430 0.935 4.600 2.785 ;
        RECT 6.670 0.895 6.840 2.050 ;
        RECT 6.670 1.495 6.970 2.050 ;
        RECT 6.670 1.495 7.570 1.665 ;
        RECT 5.130 0.895 5.300 2.465 ;
        RECT 7.765 1.675 7.935 2.465 ;
        RECT 5.130 2.295 7.935 2.465 ;
        RECT 7.765 1.675 8.220 1.845 ;
        RECT 7.160 0.960 7.460 1.220 ;
        RECT 8.325 0.920 8.495 1.220 ;
        RECT 7.160 1.040 8.495 1.220 ;
        RECT 6.815 0.480 7.115 0.710 ;
        RECT 8.115 2.045 8.340 2.215 ;
        RECT 6.815 0.540 8.845 0.710 ;
        RECT 8.675 0.540 8.845 1.705 ;
        RECT 8.620 1.535 9.455 1.705 ;
        RECT 8.450 1.535 8.460 2.169 ;
        RECT 8.460 1.535 8.470 2.159 ;
        RECT 8.470 1.535 8.480 2.149 ;
        RECT 8.480 1.535 8.490 2.139 ;
        RECT 8.490 1.535 8.500 2.129 ;
        RECT 8.500 1.535 8.510 2.119 ;
        RECT 8.510 1.535 8.520 2.109 ;
        RECT 8.520 1.535 8.530 2.099 ;
        RECT 8.530 1.535 8.540 2.089 ;
        RECT 8.540 1.535 8.550 2.079 ;
        RECT 8.550 1.535 8.560 2.069 ;
        RECT 8.560 1.535 8.570 2.059 ;
        RECT 8.570 1.535 8.580 2.049 ;
        RECT 8.580 1.535 8.590 2.039 ;
        RECT 8.590 1.535 8.600 2.029 ;
        RECT 8.600 1.535 8.610 2.019 ;
        RECT 8.610 1.535 8.620 2.009 ;
        RECT 8.415 1.970 8.425 2.204 ;
        RECT 8.425 1.960 8.435 2.194 ;
        RECT 8.435 1.950 8.445 2.184 ;
        RECT 8.445 1.940 8.451 2.180 ;
        RECT 8.340 2.045 8.350 2.215 ;
        RECT 8.350 2.035 8.360 2.215 ;
        RECT 8.360 2.025 8.370 2.215 ;
        RECT 8.370 2.015 8.380 2.215 ;
        RECT 8.380 2.005 8.390 2.215 ;
        RECT 8.390 1.995 8.400 2.215 ;
        RECT 8.400 1.985 8.410 2.215 ;
        RECT 8.410 1.975 8.416 2.215 ;
        RECT 3.975 0.530 4.145 2.340 ;
        RECT 3.855 1.125 4.155 1.295 ;
        RECT 4.780 0.530 4.950 2.815 ;
        RECT 3.975 0.530 5.545 0.700 ;
        RECT 4.780 2.645 8.245 2.815 ;
        RECT 8.670 2.295 9.485 2.465 ;
        RECT 10.280 1.610 10.450 2.630 ;
        RECT 9.725 2.460 10.450 2.630 ;
        RECT 9.650 2.395 9.660 2.629 ;
        RECT 9.660 2.405 9.670 2.629 ;
        RECT 9.670 2.415 9.680 2.629 ;
        RECT 9.680 2.425 9.690 2.629 ;
        RECT 9.690 2.435 9.700 2.629 ;
        RECT 9.700 2.445 9.710 2.629 ;
        RECT 9.710 2.455 9.720 2.629 ;
        RECT 9.720 2.460 9.726 2.630 ;
        RECT 9.560 2.305 9.570 2.539 ;
        RECT 9.570 2.315 9.580 2.549 ;
        RECT 9.580 2.325 9.590 2.559 ;
        RECT 9.590 2.335 9.600 2.569 ;
        RECT 9.600 2.345 9.610 2.579 ;
        RECT 9.610 2.355 9.620 2.589 ;
        RECT 9.620 2.365 9.630 2.599 ;
        RECT 9.630 2.375 9.640 2.609 ;
        RECT 9.640 2.385 9.650 2.619 ;
        RECT 9.485 2.295 9.495 2.465 ;
        RECT 9.495 2.295 9.505 2.475 ;
        RECT 9.505 2.295 9.515 2.485 ;
        RECT 9.515 2.295 9.525 2.495 ;
        RECT 9.525 2.295 9.535 2.505 ;
        RECT 9.535 2.295 9.545 2.515 ;
        RECT 9.545 2.295 9.555 2.525 ;
        RECT 9.555 2.295 9.561 2.535 ;
        RECT 8.595 2.295 8.605 2.529 ;
        RECT 8.605 2.295 8.615 2.519 ;
        RECT 8.615 2.295 8.625 2.509 ;
        RECT 8.625 2.295 8.635 2.499 ;
        RECT 8.635 2.295 8.645 2.489 ;
        RECT 8.645 2.295 8.655 2.479 ;
        RECT 8.655 2.295 8.665 2.469 ;
        RECT 8.665 2.295 8.671 2.465 ;
        RECT 8.320 2.570 8.330 2.804 ;
        RECT 8.330 2.560 8.340 2.794 ;
        RECT 8.340 2.550 8.350 2.784 ;
        RECT 8.350 2.540 8.360 2.774 ;
        RECT 8.360 2.530 8.370 2.764 ;
        RECT 8.370 2.520 8.380 2.754 ;
        RECT 8.380 2.510 8.390 2.744 ;
        RECT 8.390 2.500 8.400 2.734 ;
        RECT 8.400 2.490 8.410 2.724 ;
        RECT 8.410 2.480 8.420 2.714 ;
        RECT 8.420 2.470 8.430 2.704 ;
        RECT 8.430 2.460 8.440 2.694 ;
        RECT 8.440 2.450 8.450 2.684 ;
        RECT 8.450 2.440 8.460 2.674 ;
        RECT 8.460 2.430 8.470 2.664 ;
        RECT 8.470 2.420 8.480 2.654 ;
        RECT 8.480 2.410 8.490 2.644 ;
        RECT 8.490 2.400 8.500 2.634 ;
        RECT 8.500 2.390 8.510 2.624 ;
        RECT 8.510 2.380 8.520 2.614 ;
        RECT 8.520 2.370 8.530 2.604 ;
        RECT 8.530 2.360 8.540 2.594 ;
        RECT 8.540 2.350 8.550 2.584 ;
        RECT 8.550 2.340 8.560 2.574 ;
        RECT 8.560 2.330 8.570 2.564 ;
        RECT 8.570 2.320 8.580 2.554 ;
        RECT 8.580 2.310 8.590 2.544 ;
        RECT 8.590 2.300 8.596 2.540 ;
        RECT 8.245 2.645 8.255 2.815 ;
        RECT 8.255 2.635 8.265 2.815 ;
        RECT 8.265 2.625 8.275 2.815 ;
        RECT 8.275 2.615 8.285 2.815 ;
        RECT 8.285 2.605 8.295 2.815 ;
        RECT 8.295 2.595 8.305 2.815 ;
        RECT 8.305 2.585 8.315 2.815 ;
        RECT 8.315 2.575 8.321 2.815 ;
        RECT 8.255 3.040 8.595 3.210 ;
        RECT 8.845 2.645 9.330 2.815 ;
        RECT 10.325 1.195 10.535 1.365 ;
        RECT 9.675 2.915 10.630 3.085 ;
        RECT 10.630 1.225 10.640 3.085 ;
        RECT 10.640 1.235 10.650 3.085 ;
        RECT 10.650 1.245 10.660 3.085 ;
        RECT 10.660 1.255 10.670 3.085 ;
        RECT 10.670 1.265 10.680 3.085 ;
        RECT 10.680 1.275 10.690 3.085 ;
        RECT 10.690 1.285 10.700 3.085 ;
        RECT 10.700 1.295 10.710 3.085 ;
        RECT 10.710 1.305 10.720 3.085 ;
        RECT 10.720 1.315 10.730 3.085 ;
        RECT 10.730 1.325 10.740 3.085 ;
        RECT 10.740 1.335 10.750 3.085 ;
        RECT 10.750 1.345 10.760 3.085 ;
        RECT 10.760 1.355 10.770 3.085 ;
        RECT 10.770 1.365 10.780 3.085 ;
        RECT 10.780 1.375 10.790 3.085 ;
        RECT 10.790 1.385 10.800 3.085 ;
        RECT 10.625 1.215 10.631 1.455 ;
        RECT 10.535 1.195 10.545 1.365 ;
        RECT 10.545 1.195 10.555 1.375 ;
        RECT 10.555 1.195 10.565 1.385 ;
        RECT 10.565 1.195 10.575 1.395 ;
        RECT 10.575 1.195 10.585 1.405 ;
        RECT 10.585 1.195 10.595 1.415 ;
        RECT 10.595 1.195 10.605 1.425 ;
        RECT 10.605 1.195 10.615 1.435 ;
        RECT 10.615 1.195 10.625 1.445 ;
        RECT 9.600 2.850 9.610 3.084 ;
        RECT 9.610 2.860 9.620 3.084 ;
        RECT 9.620 2.870 9.630 3.084 ;
        RECT 9.630 2.880 9.640 3.084 ;
        RECT 9.640 2.890 9.650 3.084 ;
        RECT 9.650 2.900 9.660 3.084 ;
        RECT 9.660 2.910 9.670 3.084 ;
        RECT 9.670 2.915 9.676 3.085 ;
        RECT 9.405 2.655 9.415 2.889 ;
        RECT 9.415 2.665 9.425 2.899 ;
        RECT 9.425 2.675 9.435 2.909 ;
        RECT 9.435 2.685 9.445 2.919 ;
        RECT 9.445 2.695 9.455 2.929 ;
        RECT 9.455 2.705 9.465 2.939 ;
        RECT 9.465 2.715 9.475 2.949 ;
        RECT 9.475 2.725 9.485 2.959 ;
        RECT 9.485 2.735 9.495 2.969 ;
        RECT 9.495 2.745 9.505 2.979 ;
        RECT 9.505 2.755 9.515 2.989 ;
        RECT 9.515 2.765 9.525 2.999 ;
        RECT 9.525 2.775 9.535 3.009 ;
        RECT 9.535 2.785 9.545 3.019 ;
        RECT 9.545 2.795 9.555 3.029 ;
        RECT 9.555 2.805 9.565 3.039 ;
        RECT 9.565 2.815 9.575 3.049 ;
        RECT 9.575 2.825 9.585 3.059 ;
        RECT 9.585 2.835 9.595 3.069 ;
        RECT 9.595 2.840 9.601 3.080 ;
        RECT 9.330 2.645 9.340 2.815 ;
        RECT 9.340 2.645 9.350 2.825 ;
        RECT 9.350 2.645 9.360 2.835 ;
        RECT 9.360 2.645 9.370 2.845 ;
        RECT 9.370 2.645 9.380 2.855 ;
        RECT 9.380 2.645 9.390 2.865 ;
        RECT 9.390 2.645 9.400 2.875 ;
        RECT 9.400 2.645 9.406 2.885 ;
        RECT 8.770 2.645 8.780 2.879 ;
        RECT 8.780 2.645 8.790 2.869 ;
        RECT 8.790 2.645 8.800 2.859 ;
        RECT 8.800 2.645 8.810 2.849 ;
        RECT 8.810 2.645 8.820 2.839 ;
        RECT 8.820 2.645 8.830 2.829 ;
        RECT 8.830 2.645 8.840 2.819 ;
        RECT 8.840 2.645 8.846 2.815 ;
        RECT 8.765 2.650 8.771 2.890 ;
        RECT 8.595 2.820 8.605 3.210 ;
        RECT 8.605 2.810 8.615 3.210 ;
        RECT 8.615 2.800 8.625 3.210 ;
        RECT 8.625 2.790 8.635 3.210 ;
        RECT 8.635 2.780 8.645 3.210 ;
        RECT 8.645 2.770 8.655 3.210 ;
        RECT 8.655 2.760 8.665 3.210 ;
        RECT 8.665 2.750 8.675 3.210 ;
        RECT 8.675 2.740 8.685 3.210 ;
        RECT 8.685 2.730 8.695 3.210 ;
        RECT 8.695 2.720 8.705 3.210 ;
        RECT 8.705 2.710 8.715 3.210 ;
        RECT 8.715 2.700 8.725 3.210 ;
        RECT 8.725 2.690 8.735 3.210 ;
        RECT 8.735 2.680 8.745 3.210 ;
        RECT 8.745 2.670 8.755 3.210 ;
        RECT 8.755 2.660 8.765 3.210 ;
        RECT 11.365 1.650 12.820 1.820 ;
        RECT 12.650 1.650 12.820 2.135 ;
        RECT 11.850 0.725 12.020 0.945 ;
        RECT 11.550 0.725 12.020 0.895 ;
        RECT 11.850 0.775 12.950 0.945 ;
        RECT 12.650 0.775 12.950 0.955 ;
        RECT 11.330 1.105 11.500 1.470 ;
        RECT 12.100 1.125 12.400 1.470 ;
        RECT 12.460 2.340 14.095 2.440 ;
        RECT 12.470 2.330 12.486 2.560 ;
        RECT 12.450 2.350 14.095 2.440 ;
        RECT 12.480 2.320 12.486 2.560 ;
        RECT 12.440 2.360 14.095 2.440 ;
        RECT 11.875 2.390 12.486 2.560 ;
        RECT 11.875 2.390 12.495 2.549 ;
        RECT 11.875 2.390 12.505 2.539 ;
        RECT 11.875 2.390 12.515 2.529 ;
        RECT 11.875 2.390 12.525 2.519 ;
        RECT 11.875 2.390 12.535 2.509 ;
        RECT 11.875 2.390 12.545 2.499 ;
        RECT 11.875 2.390 12.555 2.489 ;
        RECT 11.330 1.300 13.170 1.470 ;
        RECT 12.485 2.315 13.170 2.485 ;
        RECT 12.430 2.370 14.095 2.440 ;
        RECT 13.000 1.300 13.170 2.485 ;
        RECT 13.000 2.270 14.095 2.440 ;
        RECT 12.420 2.380 14.095 2.440 ;
        RECT 13.925 1.780 14.095 2.440 ;
        RECT 14.200 1.540 14.370 1.950 ;
        RECT 13.925 1.780 14.370 1.950 ;
        RECT 9.930 0.785 10.100 2.280 ;
        RECT 9.930 0.785 10.670 0.955 ;
        RECT 10.955 0.995 11.150 1.165 ;
        RECT 10.980 0.995 11.150 2.190 ;
        RECT 11.525 2.020 11.695 2.910 ;
        RECT 10.980 2.020 12.315 2.190 ;
        RECT 11.525 2.740 12.565 2.910 ;
        RECT 12.715 2.665 13.510 2.835 ;
        RECT 13.550 2.625 13.585 2.835 ;
        RECT 14.965 1.650 15.135 2.795 ;
        RECT 13.625 2.625 15.135 2.795 ;
        RECT 14.965 1.650 15.445 1.820 ;
        RECT 13.585 2.625 13.595 2.825 ;
        RECT 13.595 2.625 13.605 2.815 ;
        RECT 13.605 2.625 13.615 2.805 ;
        RECT 13.615 2.625 13.625 2.795 ;
        RECT 13.510 2.665 13.520 2.835 ;
        RECT 13.520 2.655 13.530 2.835 ;
        RECT 13.530 2.645 13.540 2.835 ;
        RECT 13.540 2.635 13.550 2.835 ;
        RECT 12.640 2.665 12.650 2.899 ;
        RECT 12.650 2.665 12.660 2.889 ;
        RECT 12.660 2.665 12.670 2.879 ;
        RECT 12.670 2.665 12.680 2.869 ;
        RECT 12.680 2.665 12.690 2.859 ;
        RECT 12.690 2.665 12.700 2.849 ;
        RECT 12.700 2.665 12.710 2.839 ;
        RECT 12.710 2.665 12.716 2.835 ;
        RECT 12.565 2.740 12.575 2.910 ;
        RECT 12.575 2.730 12.585 2.910 ;
        RECT 12.585 2.720 12.595 2.910 ;
        RECT 12.595 2.710 12.605 2.910 ;
        RECT 12.605 2.700 12.615 2.910 ;
        RECT 12.615 2.690 12.625 2.910 ;
        RECT 12.625 2.680 12.635 2.910 ;
        RECT 12.635 2.670 12.641 2.910 ;
        RECT 10.880 0.930 10.890 1.164 ;
        RECT 10.890 0.940 10.900 1.164 ;
        RECT 10.900 0.950 10.910 1.164 ;
        RECT 10.910 0.960 10.920 1.164 ;
        RECT 10.920 0.970 10.930 1.164 ;
        RECT 10.930 0.980 10.940 1.164 ;
        RECT 10.940 0.990 10.950 1.164 ;
        RECT 10.950 0.995 10.956 1.165 ;
        RECT 10.745 0.795 10.755 1.029 ;
        RECT 10.755 0.805 10.765 1.039 ;
        RECT 10.765 0.815 10.775 1.049 ;
        RECT 10.775 0.825 10.785 1.059 ;
        RECT 10.785 0.835 10.795 1.069 ;
        RECT 10.795 0.845 10.805 1.079 ;
        RECT 10.805 0.855 10.815 1.089 ;
        RECT 10.815 0.865 10.825 1.099 ;
        RECT 10.825 0.875 10.835 1.109 ;
        RECT 10.835 0.885 10.845 1.119 ;
        RECT 10.845 0.895 10.855 1.129 ;
        RECT 10.855 0.905 10.865 1.139 ;
        RECT 10.865 0.915 10.875 1.149 ;
        RECT 10.875 0.920 10.881 1.160 ;
        RECT 10.670 0.785 10.680 0.955 ;
        RECT 10.680 0.785 10.690 0.965 ;
        RECT 10.690 0.785 10.700 0.975 ;
        RECT 10.700 0.785 10.710 0.985 ;
        RECT 10.710 0.785 10.720 0.995 ;
        RECT 10.720 0.785 10.730 1.005 ;
        RECT 10.730 0.785 10.740 1.015 ;
        RECT 10.740 0.785 10.746 1.025 ;
  END 
END FFSDSRHD2XHT

MACRO FFSDSRHD1XHT
  CLASS  CORE ;
  FOREIGN FFSDSRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.760 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.405 0.720 14.575 2.960 ;
        RECT 14.355 1.980 14.575 2.960 ;
        RECT 14.355 2.490 14.660 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.220 1.190 13.655 1.360 ;
        RECT 13.485 0.720 13.535 2.215 ;
        RECT 13.220 0.720 13.535 1.360 ;
        RECT 13.485 1.190 13.655 2.215 ;
        RECT 13.250 2.045 13.655 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 1.290 1.605 1.540 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.155 1.410 6.490 2.045 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.520 1.735 0.690 2.100 ;
        RECT 0.815 1.930 1.230 2.360 ;
        RECT 1.400 1.735 1.570 2.100 ;
        RECT 0.520 1.930 1.570 2.100 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.995 ;
        RECT 2.435 -0.300 2.735 0.785 ;
        RECT 3.400 -0.300 3.700 0.945 ;
        RECT 6.075 -0.300 6.375 1.130 ;
        RECT 8.870 -0.300 9.040 1.220 ;
        RECT 10.750 -0.300 11.050 0.795 ;
        RECT 12.835 -0.300 13.005 1.345 ;
        RECT 13.885 -0.300 14.055 1.120 ;
        RECT 0.000 -0.300 14.760 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.970 1.550 3.325 2.015 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.290 1.610 2.775 2.015 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 12.400 1.540 12.720 2.015 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.905 0.895 3.990 ;
        RECT 2.540 2.895 3.520 3.990 ;
        RECT 6.250 2.995 7.230 3.990 ;
        RECT 8.780 2.995 9.080 3.990 ;
        RECT 10.805 2.415 11.105 3.990 ;
        RECT 12.710 2.895 13.010 3.990 ;
        RECT 13.770 2.975 14.070 3.990 ;
        RECT 0.000 3.390 14.760 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.170 0.340 2.470 ;
        RECT 0.105 0.825 0.275 2.470 ;
        RECT 0.170 2.170 0.340 2.725 ;
        RECT 0.105 0.825 0.405 0.995 ;
        RECT 0.170 2.555 1.305 2.725 ;
        RECT 1.135 2.555 1.305 3.210 ;
        RECT 1.135 3.040 1.995 3.210 ;
        RECT 2.830 1.125 3.855 1.295 ;
        RECT 3.685 1.125 3.855 2.365 ;
        RECT 2.910 2.195 3.855 2.365 ;
        RECT 1.580 0.725 1.750 1.055 ;
        RECT 1.580 0.885 1.985 1.055 ;
        RECT 1.815 0.885 1.985 2.715 ;
        RECT 1.580 2.370 1.985 2.715 ;
        RECT 1.580 2.545 3.760 2.715 ;
        RECT 4.550 0.895 4.720 2.830 ;
        RECT 3.950 2.660 4.720 2.830 ;
        RECT 3.875 2.595 3.885 2.829 ;
        RECT 3.885 2.605 3.895 2.829 ;
        RECT 3.895 2.615 3.905 2.829 ;
        RECT 3.905 2.625 3.915 2.829 ;
        RECT 3.915 2.635 3.925 2.829 ;
        RECT 3.925 2.645 3.935 2.829 ;
        RECT 3.935 2.655 3.945 2.829 ;
        RECT 3.945 2.660 3.951 2.830 ;
        RECT 3.835 2.555 3.845 2.789 ;
        RECT 3.845 2.565 3.855 2.799 ;
        RECT 3.855 2.575 3.865 2.809 ;
        RECT 3.865 2.585 3.875 2.819 ;
        RECT 3.760 2.545 3.770 2.715 ;
        RECT 3.770 2.545 3.780 2.725 ;
        RECT 3.780 2.545 3.790 2.735 ;
        RECT 3.790 2.545 3.800 2.745 ;
        RECT 3.800 2.545 3.810 2.755 ;
        RECT 3.810 2.545 3.820 2.765 ;
        RECT 3.820 2.545 3.830 2.775 ;
        RECT 3.830 2.545 3.836 2.785 ;
        RECT 6.690 0.960 6.860 2.115 ;
        RECT 6.595 0.960 6.895 1.130 ;
        RECT 6.690 1.500 7.465 1.670 ;
        RECT 5.250 0.895 5.420 2.465 ;
        RECT 7.645 1.680 7.815 2.465 ;
        RECT 5.250 2.295 7.815 2.465 ;
        RECT 7.880 1.550 8.050 1.850 ;
        RECT 7.645 1.680 8.050 1.850 ;
        RECT 7.105 0.960 7.405 1.230 ;
        RECT 7.105 1.060 8.340 1.230 ;
        RECT 8.170 1.060 8.340 1.360 ;
        RECT 6.735 0.480 7.035 0.695 ;
        RECT 7.995 2.045 8.120 2.215 ;
        RECT 8.230 1.580 8.295 2.215 ;
        RECT 6.735 0.525 8.690 0.695 ;
        RECT 8.520 0.525 8.690 1.750 ;
        RECT 8.400 1.580 9.285 1.750 ;
        RECT 8.295 1.580 8.305 2.104 ;
        RECT 8.305 1.580 8.315 2.094 ;
        RECT 8.315 1.580 8.325 2.084 ;
        RECT 8.325 1.580 8.335 2.074 ;
        RECT 8.335 1.580 8.345 2.064 ;
        RECT 8.345 1.580 8.355 2.054 ;
        RECT 8.355 1.580 8.365 2.044 ;
        RECT 8.365 1.580 8.375 2.034 ;
        RECT 8.375 1.580 8.385 2.024 ;
        RECT 8.385 1.580 8.395 2.014 ;
        RECT 8.395 1.580 8.401 2.010 ;
        RECT 8.120 2.045 8.130 2.215 ;
        RECT 8.130 2.035 8.140 2.215 ;
        RECT 8.140 2.025 8.150 2.215 ;
        RECT 8.150 2.015 8.160 2.215 ;
        RECT 8.160 2.005 8.170 2.215 ;
        RECT 8.170 1.995 8.180 2.215 ;
        RECT 8.180 1.985 8.190 2.215 ;
        RECT 8.190 1.975 8.200 2.215 ;
        RECT 8.200 1.965 8.210 2.215 ;
        RECT 8.210 1.955 8.220 2.215 ;
        RECT 8.220 1.945 8.230 2.215 ;
        RECT 4.035 0.545 4.205 2.430 ;
        RECT 4.900 0.545 5.070 2.835 ;
        RECT 4.035 0.545 5.665 0.715 ;
        RECT 4.900 2.645 8.125 2.815 ;
        RECT 8.550 2.295 9.310 2.465 ;
        RECT 9.485 2.395 10.210 2.565 ;
        RECT 10.040 2.395 10.210 2.770 ;
        RECT 9.410 2.330 9.420 2.564 ;
        RECT 9.420 2.340 9.430 2.564 ;
        RECT 9.430 2.350 9.440 2.564 ;
        RECT 9.440 2.360 9.450 2.564 ;
        RECT 9.450 2.370 9.460 2.564 ;
        RECT 9.460 2.380 9.470 2.564 ;
        RECT 9.470 2.390 9.480 2.564 ;
        RECT 9.480 2.395 9.486 2.565 ;
        RECT 9.385 2.305 9.395 2.539 ;
        RECT 9.395 2.315 9.405 2.549 ;
        RECT 9.405 2.320 9.411 2.560 ;
        RECT 9.310 2.295 9.320 2.465 ;
        RECT 9.320 2.295 9.330 2.475 ;
        RECT 9.330 2.295 9.340 2.485 ;
        RECT 9.340 2.295 9.350 2.495 ;
        RECT 9.350 2.295 9.360 2.505 ;
        RECT 9.360 2.295 9.370 2.515 ;
        RECT 9.370 2.295 9.380 2.525 ;
        RECT 9.380 2.295 9.386 2.535 ;
        RECT 8.475 2.295 8.485 2.529 ;
        RECT 8.485 2.295 8.495 2.519 ;
        RECT 8.495 2.295 8.505 2.509 ;
        RECT 8.505 2.295 8.515 2.499 ;
        RECT 8.515 2.295 8.525 2.489 ;
        RECT 8.525 2.295 8.535 2.479 ;
        RECT 8.535 2.295 8.545 2.469 ;
        RECT 8.545 2.295 8.551 2.465 ;
        RECT 8.200 2.570 8.210 2.804 ;
        RECT 8.210 2.560 8.220 2.794 ;
        RECT 8.220 2.550 8.230 2.784 ;
        RECT 8.230 2.540 8.240 2.774 ;
        RECT 8.240 2.530 8.250 2.764 ;
        RECT 8.250 2.520 8.260 2.754 ;
        RECT 8.260 2.510 8.270 2.744 ;
        RECT 8.270 2.500 8.280 2.734 ;
        RECT 8.280 2.490 8.290 2.724 ;
        RECT 8.290 2.480 8.300 2.714 ;
        RECT 8.300 2.470 8.310 2.704 ;
        RECT 8.310 2.460 8.320 2.694 ;
        RECT 8.320 2.450 8.330 2.684 ;
        RECT 8.330 2.440 8.340 2.674 ;
        RECT 8.340 2.430 8.350 2.664 ;
        RECT 8.350 2.420 8.360 2.654 ;
        RECT 8.360 2.410 8.370 2.644 ;
        RECT 8.370 2.400 8.380 2.634 ;
        RECT 8.380 2.390 8.390 2.624 ;
        RECT 8.390 2.380 8.400 2.614 ;
        RECT 8.400 2.370 8.410 2.604 ;
        RECT 8.410 2.360 8.420 2.594 ;
        RECT 8.420 2.350 8.430 2.584 ;
        RECT 8.430 2.340 8.440 2.574 ;
        RECT 8.440 2.330 8.450 2.564 ;
        RECT 8.450 2.320 8.460 2.554 ;
        RECT 8.460 2.310 8.470 2.544 ;
        RECT 8.470 2.300 8.476 2.540 ;
        RECT 8.125 2.645 8.135 2.815 ;
        RECT 8.135 2.635 8.145 2.815 ;
        RECT 8.145 2.625 8.155 2.815 ;
        RECT 8.155 2.615 8.165 2.815 ;
        RECT 8.165 2.605 8.175 2.815 ;
        RECT 8.175 2.595 8.185 2.815 ;
        RECT 8.185 2.585 8.195 2.815 ;
        RECT 8.195 2.575 8.201 2.815 ;
        RECT 8.065 3.040 8.430 3.210 ;
        RECT 8.700 2.645 9.155 2.815 ;
        RECT 9.330 2.745 9.770 2.915 ;
        RECT 9.600 2.745 9.770 3.120 ;
        RECT 10.060 1.270 10.360 1.440 ;
        RECT 10.190 1.270 10.360 1.825 ;
        RECT 10.190 1.655 10.560 1.825 ;
        RECT 10.390 1.655 10.560 3.120 ;
        RECT 9.600 2.950 10.560 3.120 ;
        RECT 9.255 2.680 9.265 2.914 ;
        RECT 9.265 2.690 9.275 2.914 ;
        RECT 9.275 2.700 9.285 2.914 ;
        RECT 9.285 2.710 9.295 2.914 ;
        RECT 9.295 2.720 9.305 2.914 ;
        RECT 9.305 2.730 9.315 2.914 ;
        RECT 9.315 2.740 9.325 2.914 ;
        RECT 9.325 2.745 9.331 2.915 ;
        RECT 9.230 2.655 9.240 2.889 ;
        RECT 9.240 2.665 9.250 2.899 ;
        RECT 9.250 2.670 9.256 2.910 ;
        RECT 9.155 2.645 9.165 2.815 ;
        RECT 9.165 2.645 9.175 2.825 ;
        RECT 9.175 2.645 9.185 2.835 ;
        RECT 9.185 2.645 9.195 2.845 ;
        RECT 9.195 2.645 9.205 2.855 ;
        RECT 9.205 2.645 9.215 2.865 ;
        RECT 9.215 2.645 9.225 2.875 ;
        RECT 9.225 2.645 9.231 2.885 ;
        RECT 8.625 2.645 8.635 2.879 ;
        RECT 8.635 2.645 8.645 2.869 ;
        RECT 8.645 2.645 8.655 2.859 ;
        RECT 8.655 2.645 8.665 2.849 ;
        RECT 8.665 2.645 8.675 2.839 ;
        RECT 8.675 2.645 8.685 2.829 ;
        RECT 8.685 2.645 8.695 2.819 ;
        RECT 8.695 2.645 8.701 2.815 ;
        RECT 8.600 2.670 8.610 2.904 ;
        RECT 8.610 2.660 8.620 2.894 ;
        RECT 8.620 2.650 8.626 2.890 ;
        RECT 8.430 2.840 8.440 3.210 ;
        RECT 8.440 2.830 8.450 3.210 ;
        RECT 8.450 2.820 8.460 3.210 ;
        RECT 8.460 2.810 8.470 3.210 ;
        RECT 8.470 2.800 8.480 3.210 ;
        RECT 8.480 2.790 8.490 3.210 ;
        RECT 8.490 2.780 8.500 3.210 ;
        RECT 8.500 2.770 8.510 3.210 ;
        RECT 8.510 2.760 8.520 3.210 ;
        RECT 8.520 2.750 8.530 3.210 ;
        RECT 8.530 2.740 8.540 3.210 ;
        RECT 8.540 2.730 8.550 3.210 ;
        RECT 8.550 2.720 8.560 3.210 ;
        RECT 8.560 2.710 8.570 3.210 ;
        RECT 8.570 2.700 8.580 3.210 ;
        RECT 8.580 2.690 8.590 3.210 ;
        RECT 8.590 2.680 8.600 3.210 ;
        RECT 11.310 0.760 11.480 1.280 ;
        RECT 11.180 1.110 11.480 1.280 ;
        RECT 11.310 0.760 12.390 0.930 ;
        RECT 12.220 0.760 12.390 1.280 ;
        RECT 12.220 1.110 12.520 1.280 ;
        RECT 11.090 1.460 11.260 1.760 ;
        RECT 11.700 1.110 12.000 1.630 ;
        RECT 11.090 1.460 12.000 1.630 ;
        RECT 11.830 1.110 12.000 2.365 ;
        RECT 12.900 1.540 13.070 2.365 ;
        RECT 11.830 2.195 13.070 2.365 ;
        RECT 12.900 1.540 13.305 1.840 ;
        RECT 9.650 0.900 9.820 2.215 ;
        RECT 9.650 2.045 9.950 2.215 ;
        RECT 9.650 0.900 10.435 1.070 ;
        RECT 10.670 1.060 10.910 1.230 ;
        RECT 10.740 1.060 10.910 2.110 ;
        RECT 10.740 1.940 11.495 2.110 ;
        RECT 11.325 1.940 11.495 2.715 ;
        RECT 11.920 2.545 12.220 2.965 ;
        RECT 13.980 1.505 14.150 2.715 ;
        RECT 11.325 2.545 14.150 2.715 ;
        RECT 13.980 1.505 14.225 1.805 ;
        RECT 10.595 0.995 10.605 1.229 ;
        RECT 10.605 1.005 10.615 1.229 ;
        RECT 10.615 1.015 10.625 1.229 ;
        RECT 10.625 1.025 10.635 1.229 ;
        RECT 10.635 1.035 10.645 1.229 ;
        RECT 10.645 1.045 10.655 1.229 ;
        RECT 10.655 1.055 10.665 1.229 ;
        RECT 10.665 1.060 10.671 1.230 ;
        RECT 10.510 0.910 10.520 1.144 ;
        RECT 10.520 0.920 10.530 1.154 ;
        RECT 10.530 0.930 10.540 1.164 ;
        RECT 10.540 0.940 10.550 1.174 ;
        RECT 10.550 0.950 10.560 1.184 ;
        RECT 10.560 0.960 10.570 1.194 ;
        RECT 10.570 0.970 10.580 1.204 ;
        RECT 10.580 0.980 10.590 1.214 ;
        RECT 10.590 0.985 10.596 1.225 ;
        RECT 10.435 0.900 10.445 1.070 ;
        RECT 10.445 0.900 10.455 1.080 ;
        RECT 10.455 0.900 10.465 1.090 ;
        RECT 10.465 0.900 10.475 1.100 ;
        RECT 10.475 0.900 10.485 1.110 ;
        RECT 10.485 0.900 10.495 1.120 ;
        RECT 10.495 0.900 10.505 1.130 ;
        RECT 10.505 0.900 10.511 1.140 ;
  END 
END FFSDSRHD1XHT

MACRO FFSDSHQHDMXHT
  CLASS  CORE ;
  FOREIGN FFSDSHQHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.710 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 12.370 0.980 12.620 2.455 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.160 1.135 1.775 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.575 0.380 2.020 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.870 ;
        RECT 2.545 -0.300 2.845 0.595 ;
        RECT 3.525 -0.300 3.825 0.595 ;
        RECT 4.375 -0.300 4.675 0.595 ;
        RECT 7.370 -0.300 7.670 0.595 ;
        RECT 8.900 -0.300 9.200 0.595 ;
        RECT 10.935 -0.300 11.105 0.805 ;
        RECT 11.820 -0.300 11.990 0.780 ;
        RECT 0.000 -0.300 12.710 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 4.495 1.605 5.010 2.020 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.345 1.530 2.785 2.020 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 10.755 2.485 10.995 2.915 ;
        RECT 8.185 2.745 11.445 2.915 ;
        RECT 11.145 2.745 11.445 2.920 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.655 0.955 3.990 ;
        RECT 2.555 2.470 2.730 3.990 ;
        RECT 3.555 2.780 3.855 3.990 ;
        RECT 4.375 2.780 4.675 3.990 ;
        RECT 7.385 2.930 7.685 3.990 ;
        RECT 8.745 3.095 9.045 3.990 ;
        RECT 10.770 3.095 11.070 3.990 ;
        RECT 11.850 2.910 12.020 3.990 ;
        RECT 0.000 3.390 12.710 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 2.220 0.340 2.520 ;
        RECT 0.105 1.075 0.730 1.245 ;
        RECT 0.560 1.075 0.730 2.390 ;
        RECT 0.170 2.220 0.730 2.390 ;
        RECT 1.355 1.510 1.525 2.125 ;
        RECT 0.560 1.955 1.525 2.125 ;
        RECT 1.355 1.510 1.630 1.810 ;
        RECT 3.390 1.605 3.560 1.910 ;
        RECT 3.390 1.605 4.285 1.780 ;
        RECT 3.985 1.125 4.285 2.215 ;
        RECT 4.925 1.125 5.650 1.295 ;
        RECT 5.480 1.125 5.650 2.215 ;
        RECT 5.295 2.045 5.650 2.215 ;
        RECT 1.640 1.070 1.980 1.260 ;
        RECT 1.640 0.960 1.810 1.260 ;
        RECT 1.575 2.330 1.875 2.840 ;
        RECT 1.810 1.070 1.980 2.585 ;
        RECT 1.575 2.330 1.980 2.585 ;
        RECT 2.485 0.775 2.655 1.240 ;
        RECT 1.640 1.070 2.655 1.240 ;
        RECT 2.485 0.775 6.050 0.945 ;
        RECT 5.880 0.775 6.050 2.320 ;
        RECT 6.600 1.060 6.770 2.400 ;
        RECT 7.610 1.675 7.780 2.210 ;
        RECT 6.600 2.040 7.780 2.210 ;
        RECT 7.610 1.675 7.985 1.845 ;
        RECT 7.260 1.220 7.430 1.820 ;
        RECT 8.345 1.125 8.645 1.390 ;
        RECT 7.260 1.220 8.965 1.390 ;
        RECT 8.795 1.220 8.965 2.215 ;
        RECT 7.960 2.045 8.965 2.215 ;
        RECT 8.795 1.515 9.085 1.815 ;
        RECT 3.005 1.125 3.185 2.600 ;
        RECT 3.005 1.125 3.305 1.295 ;
        RECT 3.005 2.115 3.305 2.600 ;
        RECT 5.115 2.430 5.415 2.700 ;
        RECT 3.005 2.430 5.415 2.600 ;
        RECT 6.250 0.650 6.420 2.700 ;
        RECT 5.115 2.530 6.420 2.700 ;
        RECT 6.980 0.650 7.150 0.945 ;
        RECT 6.250 0.650 7.150 0.830 ;
        RECT 6.980 0.775 9.480 0.945 ;
        RECT 9.310 0.775 9.480 1.610 ;
        RECT 9.310 1.310 9.845 1.610 ;
        RECT 7.545 2.395 7.715 2.750 ;
        RECT 6.715 2.580 7.715 2.750 ;
        RECT 9.270 1.925 9.440 2.565 ;
        RECT 7.545 2.395 9.440 2.565 ;
        RECT 10.030 0.985 10.200 2.095 ;
        RECT 9.270 1.925 10.200 2.095 ;
        RECT 10.030 0.985 10.380 1.285 ;
        RECT 10.380 1.480 10.550 2.530 ;
        RECT 9.820 2.360 10.550 2.530 ;
        RECT 9.855 0.570 10.730 0.740 ;
        RECT 10.560 0.570 10.730 1.705 ;
        RECT 10.380 1.480 10.730 1.705 ;
        RECT 10.380 1.535 11.765 1.705 ;
        RECT 11.595 1.470 11.765 1.770 ;
        RECT 10.730 1.885 10.900 2.185 ;
        RECT 10.935 1.055 11.105 1.355 ;
        RECT 10.730 2.015 11.495 2.185 ;
        RECT 11.325 2.015 11.495 2.500 ;
        RECT 10.935 1.110 12.190 1.280 ;
        RECT 12.000 1.110 12.190 2.500 ;
        RECT 11.325 2.330 12.190 2.500 ;
  END 
END FFSDSHQHDMXHT

MACRO FFSDSHQHD3XHT
  CLASS  CORE ;
  FOREIGN FFSDSHQHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.400 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 15.020 0.480 15.190 1.120 ;
        RECT 15.020 2.405 15.190 3.045 ;
        RECT 15.020 0.950 16.305 1.120 ;
        RECT 15.940 0.950 16.305 2.705 ;
        RECT 15.020 2.405 16.305 2.705 ;
        RECT 15.995 0.480 16.305 3.045 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.205 1.165 1.770 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.545 0.380 2.020 ;
        RECT 0.150 0.755 0.450 0.945 ;
        RECT 1.215 0.485 1.385 0.945 ;
        RECT 0.150 0.775 1.385 0.945 ;
        RECT 1.215 0.485 2.155 0.655 ;
        RECT 0.265 2.580 0.450 2.840 ;
        RECT 0.150 2.670 0.450 2.840 ;
        RECT 0.265 2.580 1.340 2.750 ;
        RECT 0.150 2.670 1.340 2.750 ;
        RECT 1.170 2.580 1.340 3.190 ;
        RECT 1.170 3.020 2.310 3.190 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.595 ;
        RECT 2.550 -0.300 2.850 0.595 ;
        RECT 3.475 -0.300 3.775 0.595 ;
        RECT 4.435 -0.300 4.735 0.595 ;
        RECT 5.535 -0.300 5.855 0.595 ;
        RECT 7.585 -0.300 7.885 0.595 ;
        RECT 9.445 -0.300 9.745 0.595 ;
        RECT 10.990 -0.300 11.290 0.655 ;
        RECT 13.275 -0.300 13.445 0.800 ;
        RECT 14.500 -0.300 14.670 0.780 ;
        RECT 15.475 -0.300 15.775 0.715 ;
        RECT 0.000 -0.300 16.400 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 4.590 1.605 5.085 2.020 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.145 1.530 2.505 2.020 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 9.260 2.665 14.095 2.795 ;
        RECT 9.260 2.320 9.430 2.795 ;
        RECT 10.975 2.625 11.145 2.835 ;
        RECT 9.260 2.625 11.145 2.795 ;
        RECT 13.570 2.555 14.095 2.835 ;
        RECT 10.975 2.665 14.095 2.835 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.975 0.955 3.990 ;
        RECT 2.555 2.860 2.730 3.990 ;
        RECT 3.670 2.830 3.840 3.990 ;
        RECT 4.455 2.875 4.755 3.990 ;
        RECT 7.425 2.975 7.725 3.990 ;
        RECT 8.560 2.910 8.730 3.990 ;
        RECT 10.530 2.975 10.830 3.990 ;
        RECT 13.405 3.015 13.705 3.990 ;
        RECT 14.500 2.905 14.670 3.990 ;
        RECT 15.540 2.910 15.710 3.990 ;
        RECT 0.000 3.390 16.400 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 0.730 1.295 ;
        RECT 0.560 1.125 0.730 2.400 ;
        RECT 0.105 2.230 0.730 2.400 ;
        RECT 1.345 1.590 1.515 2.120 ;
        RECT 0.560 1.950 1.515 2.120 ;
        RECT 1.345 1.590 1.965 1.760 ;
        RECT 1.795 1.525 1.965 1.825 ;
        RECT 3.430 1.605 3.600 1.905 ;
        RECT 3.430 1.605 4.325 1.780 ;
        RECT 4.025 1.125 4.325 2.215 ;
        RECT 4.985 1.125 5.750 1.295 ;
        RECT 5.580 1.125 5.750 2.370 ;
        RECT 5.375 2.200 5.750 2.370 ;
        RECT 1.575 2.330 1.875 2.840 ;
        RECT 1.575 1.120 2.855 1.300 ;
        RECT 2.685 0.775 2.855 2.500 ;
        RECT 1.575 2.330 2.855 2.500 ;
        RECT 2.685 0.775 6.160 0.945 ;
        RECT 5.990 0.775 6.160 2.660 ;
        RECT 6.690 1.060 6.860 2.400 ;
        RECT 6.690 2.040 7.560 2.210 ;
        RECT 7.960 1.600 8.115 1.900 ;
        RECT 7.815 1.600 7.825 2.034 ;
        RECT 7.825 1.600 7.835 2.024 ;
        RECT 7.835 1.600 7.845 2.014 ;
        RECT 7.845 1.600 7.855 2.004 ;
        RECT 7.855 1.600 7.865 1.994 ;
        RECT 7.865 1.600 7.875 1.984 ;
        RECT 7.875 1.600 7.885 1.974 ;
        RECT 7.885 1.600 7.895 1.964 ;
        RECT 7.895 1.600 7.905 1.954 ;
        RECT 7.905 1.600 7.915 1.944 ;
        RECT 7.915 1.600 7.925 1.934 ;
        RECT 7.925 1.600 7.935 1.924 ;
        RECT 7.935 1.600 7.945 1.914 ;
        RECT 7.945 1.600 7.955 1.904 ;
        RECT 7.955 1.600 7.961 1.900 ;
        RECT 7.650 1.950 7.660 2.200 ;
        RECT 7.660 1.940 7.670 2.190 ;
        RECT 7.670 1.930 7.680 2.180 ;
        RECT 7.680 1.920 7.690 2.170 ;
        RECT 7.690 1.910 7.700 2.160 ;
        RECT 7.700 1.900 7.710 2.150 ;
        RECT 7.710 1.890 7.720 2.140 ;
        RECT 7.720 1.880 7.730 2.130 ;
        RECT 7.730 1.870 7.740 2.120 ;
        RECT 7.740 1.860 7.750 2.110 ;
        RECT 7.750 1.850 7.760 2.100 ;
        RECT 7.760 1.840 7.770 2.090 ;
        RECT 7.770 1.830 7.780 2.080 ;
        RECT 7.780 1.820 7.790 2.070 ;
        RECT 7.790 1.810 7.800 2.060 ;
        RECT 7.800 1.800 7.810 2.050 ;
        RECT 7.810 1.790 7.816 2.044 ;
        RECT 7.560 2.040 7.570 2.210 ;
        RECT 7.570 2.030 7.580 2.210 ;
        RECT 7.580 2.020 7.590 2.210 ;
        RECT 7.590 2.010 7.600 2.210 ;
        RECT 7.600 2.000 7.610 2.210 ;
        RECT 7.610 1.990 7.620 2.210 ;
        RECT 7.620 1.980 7.630 2.210 ;
        RECT 7.630 1.970 7.640 2.210 ;
        RECT 7.640 1.960 7.650 2.210 ;
        RECT 7.350 1.125 7.520 1.730 ;
        RECT 7.350 1.125 8.825 1.295 ;
        RECT 8.300 1.125 8.470 2.380 ;
        RECT 8.040 2.080 8.470 2.380 ;
        RECT 8.300 1.125 8.825 1.475 ;
        RECT 8.300 1.305 9.275 1.475 ;
        RECT 9.055 1.305 9.275 1.705 ;
        RECT 9.055 1.535 11.080 1.705 ;
        RECT 3.045 1.125 3.225 2.615 ;
        RECT 3.045 1.125 3.345 1.295 ;
        RECT 3.045 2.105 3.345 2.615 ;
        RECT 3.045 2.430 5.135 2.600 ;
        RECT 4.965 2.430 5.135 3.145 ;
        RECT 4.965 2.885 5.495 3.145 ;
        RECT 6.340 0.550 6.510 3.145 ;
        RECT 4.965 2.975 6.510 3.145 ;
        RECT 6.340 0.550 7.200 0.730 ;
        RECT 7.030 0.550 7.200 0.945 ;
        RECT 7.030 0.775 9.935 0.945 ;
        RECT 9.765 0.775 9.935 1.355 ;
        RECT 9.765 1.185 11.915 1.355 ;
        RECT 11.745 1.185 11.915 1.685 ;
        RECT 7.055 2.560 7.225 3.140 ;
        RECT 6.800 2.970 7.225 3.140 ;
        RECT 7.055 2.560 9.080 2.730 ;
        RECT 8.910 1.925 9.080 3.190 ;
        RECT 8.910 3.020 9.515 3.190 ;
        RECT 11.485 1.965 12.425 2.105 ;
        RECT 11.495 1.965 12.425 2.115 ;
        RECT 11.505 1.965 12.425 2.125 ;
        RECT 8.910 1.925 11.585 2.095 ;
        RECT 8.910 1.935 11.595 2.095 ;
        RECT 8.910 1.945 11.605 2.095 ;
        RECT 8.910 1.955 11.615 2.095 ;
        RECT 12.255 0.885 12.425 2.135 ;
        RECT 11.515 1.965 12.425 2.135 ;
        RECT 11.480 3.015 12.450 3.185 ;
        RECT 10.135 0.705 10.305 1.005 ;
        RECT 11.270 2.315 12.790 2.455 ;
        RECT 11.280 2.315 12.790 2.465 ;
        RECT 11.290 2.315 12.790 2.475 ;
        RECT 9.610 2.275 11.340 2.445 ;
        RECT 9.610 2.285 11.350 2.445 ;
        RECT 9.610 2.295 11.360 2.445 ;
        RECT 9.610 2.305 11.370 2.445 ;
        RECT 11.840 0.530 12.010 1.005 ;
        RECT 10.135 0.835 12.010 1.005 ;
        RECT 11.840 0.530 12.790 0.700 ;
        RECT 12.620 0.530 12.790 2.485 ;
        RECT 11.300 2.315 12.790 2.485 ;
        RECT 12.620 1.000 13.490 1.170 ;
        RECT 13.320 1.000 13.490 1.820 ;
        RECT 13.320 1.650 15.305 1.820 ;
        RECT 12.970 1.470 13.140 2.345 ;
        RECT 13.670 1.060 13.840 1.360 ;
        RECT 13.975 2.025 14.275 2.345 ;
        RECT 12.970 2.170 14.275 2.345 ;
        RECT 13.670 1.125 14.695 1.295 ;
        RECT 14.525 1.125 14.695 1.470 ;
        RECT 14.525 1.300 15.710 1.470 ;
        RECT 13.975 2.025 15.710 2.200 ;
        RECT 15.540 1.300 15.710 2.200 ;
  END 
END FFSDSHQHD3XHT

MACRO FFSDSHQHD1XHT
  CLASS  CORE ;
  FOREIGN FFSDSHQHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.710 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 12.370 0.720 12.620 2.965 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.240 1.165 1.765 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.575 0.380 2.020 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.045 ;
        RECT 2.545 -0.300 2.845 0.595 ;
        RECT 3.525 -0.300 3.825 0.595 ;
        RECT 4.475 -0.300 4.775 0.595 ;
        RECT 7.410 -0.300 7.710 0.595 ;
        RECT 8.900 -0.300 9.200 0.595 ;
        RECT 10.895 -0.300 11.065 0.805 ;
        RECT 11.850 -0.300 12.020 0.780 ;
        RECT 0.000 -0.300 12.710 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 4.495 1.540 5.010 2.020 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.345 1.530 2.785 2.020 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 8.300 2.745 8.485 3.010 ;
        RECT 8.185 2.840 8.485 3.010 ;
        RECT 10.755 2.495 10.995 2.915 ;
        RECT 8.300 2.745 11.445 2.915 ;
        RECT 8.185 2.840 11.445 2.915 ;
        RECT 11.145 2.745 11.445 2.920 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.655 0.955 3.990 ;
        RECT 2.555 2.470 2.730 3.990 ;
        RECT 3.555 2.745 3.855 3.990 ;
        RECT 4.375 2.745 4.675 3.990 ;
        RECT 7.385 2.885 7.685 3.990 ;
        RECT 8.770 3.095 9.070 3.990 ;
        RECT 10.770 3.095 11.070 3.990 ;
        RECT 11.850 2.910 12.020 3.990 ;
        RECT 0.000 3.390 12.710 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.010 0.340 1.395 ;
        RECT 0.170 2.220 0.340 2.520 ;
        RECT 0.170 1.225 0.730 1.395 ;
        RECT 0.560 1.225 0.730 2.390 ;
        RECT 0.170 2.220 0.730 2.390 ;
        RECT 1.355 1.510 1.525 2.115 ;
        RECT 0.560 1.945 1.525 2.115 ;
        RECT 1.355 1.510 1.630 1.810 ;
        RECT 3.390 1.605 3.560 1.910 ;
        RECT 3.390 1.605 4.285 1.780 ;
        RECT 3.985 1.125 4.285 2.215 ;
        RECT 5.025 1.125 5.650 1.295 ;
        RECT 5.480 1.125 5.650 2.215 ;
        RECT 5.295 2.045 5.650 2.215 ;
        RECT 1.640 0.960 1.980 1.260 ;
        RECT 1.575 2.330 1.875 2.840 ;
        RECT 1.810 0.960 1.980 2.585 ;
        RECT 1.575 2.330 1.980 2.585 ;
        RECT 2.545 0.775 2.715 1.130 ;
        RECT 1.640 0.960 2.715 1.130 ;
        RECT 2.545 0.775 6.040 0.945 ;
        RECT 5.870 0.775 6.040 2.320 ;
        RECT 6.570 1.060 6.740 2.355 ;
        RECT 7.610 1.675 7.780 2.210 ;
        RECT 6.570 2.040 7.780 2.210 ;
        RECT 7.610 1.675 7.990 1.845 ;
        RECT 7.260 1.220 7.430 1.820 ;
        RECT 8.345 1.125 8.645 1.390 ;
        RECT 7.260 1.220 8.965 1.390 ;
        RECT 8.795 1.220 8.965 2.215 ;
        RECT 7.960 2.045 8.965 2.215 ;
        RECT 8.795 1.515 9.085 1.815 ;
        RECT 3.005 1.125 3.185 2.565 ;
        RECT 3.005 2.255 3.240 2.565 ;
        RECT 3.005 1.125 3.305 1.295 ;
        RECT 5.115 2.395 5.415 2.675 ;
        RECT 3.005 2.395 5.415 2.565 ;
        RECT 6.220 0.690 6.390 2.675 ;
        RECT 5.115 2.505 6.390 2.675 ;
        RECT 6.950 0.690 7.120 0.945 ;
        RECT 6.220 0.690 7.120 0.870 ;
        RECT 6.950 0.775 9.480 0.945 ;
        RECT 9.310 0.775 9.480 1.610 ;
        RECT 9.310 1.310 9.825 1.610 ;
        RECT 7.545 2.395 7.715 2.705 ;
        RECT 6.685 2.535 7.715 2.705 ;
        RECT 7.545 2.395 9.440 2.565 ;
        RECT 9.270 1.925 9.440 2.565 ;
        RECT 10.005 0.985 10.175 2.095 ;
        RECT 9.270 1.925 10.175 2.095 ;
        RECT 10.005 0.985 10.335 1.285 ;
        RECT 9.855 0.570 10.685 0.740 ;
        RECT 10.380 1.480 10.550 2.530 ;
        RECT 9.820 2.360 10.550 2.530 ;
        RECT 10.515 0.570 10.685 1.695 ;
        RECT 10.380 1.480 10.685 1.695 ;
        RECT 10.380 1.525 11.830 1.695 ;
        RECT 10.730 1.885 10.900 2.185 ;
        RECT 10.730 1.930 11.495 2.100 ;
        RECT 11.325 1.930 11.495 2.500 ;
        RECT 10.870 1.125 12.180 1.295 ;
        RECT 12.010 1.125 12.180 2.500 ;
        RECT 11.325 2.330 12.180 2.500 ;
  END 
END FFSDSHQHD1XHT

MACRO FFSDSHDMXHT
  CLASS  CORE ;
  FOREIGN FFSDSHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.890 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.550 1.060 11.790 1.360 ;
        RECT 11.580 1.060 11.790 2.435 ;
        RECT 11.550 1.980 11.790 2.435 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.445 1.125 10.970 1.295 ;
        RECT 10.760 1.125 10.970 2.240 ;
        RECT 10.445 2.070 10.970 2.240 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.425 -0.300 2.725 0.595 ;
        RECT 3.305 -0.300 3.605 0.595 ;
        RECT 5.925 -0.300 6.225 0.745 ;
        RECT 7.165 -0.300 7.335 0.850 ;
        RECT 9.150 -0.300 9.320 0.640 ;
        RECT 10.995 -0.300 11.295 0.595 ;
        RECT 0.000 -0.300 11.890 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.740 1.525 3.230 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.530 0.520 7.700 1.910 ;
        RECT 6.885 1.610 7.700 1.910 ;
        RECT 7.530 0.520 8.905 0.690 ;
        RECT 8.735 0.520 8.905 1.145 ;
        RECT 9.595 0.540 9.765 1.145 ;
        RECT 8.735 0.920 9.765 1.145 ;
        RECT 9.595 0.540 10.055 0.710 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.580 2.740 3.220 3.990 ;
        RECT 5.855 3.160 6.155 3.990 ;
        RECT 7.100 3.160 7.400 3.990 ;
        RECT 9.105 2.770 9.405 3.990 ;
        RECT 9.810 2.880 9.980 3.990 ;
        RECT 10.995 2.935 11.295 3.990 ;
        RECT 0.000 3.390 11.890 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.525 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.070 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.965 0.775 2.135 1.035 ;
        RECT 1.530 0.865 2.135 1.035 ;
        RECT 1.965 0.775 4.510 0.945 ;
        RECT 4.340 0.775 4.510 2.280 ;
        RECT 4.340 1.960 4.520 2.280 ;
        RECT 4.340 1.970 4.530 2.280 ;
        RECT 4.340 1.980 4.540 2.280 ;
        RECT 5.040 1.255 5.245 1.425 ;
        RECT 5.040 0.900 5.210 1.425 ;
        RECT 5.075 1.255 5.245 2.280 ;
        RECT 5.075 1.595 6.355 1.765 ;
        RECT 6.535 1.060 6.705 2.215 ;
        RECT 6.405 2.045 6.705 2.215 ;
        RECT 6.535 1.060 7.350 1.360 ;
        RECT 2.725 1.125 3.585 1.295 ;
        RECT 2.785 2.190 3.585 2.360 ;
        RECT 3.415 1.125 3.585 2.980 ;
        RECT 3.415 1.525 3.710 1.825 ;
        RECT 3.415 2.810 8.045 2.980 ;
        RECT 3.765 1.125 4.085 1.295 ;
        RECT 3.915 1.125 4.085 2.630 ;
        RECT 4.690 0.535 4.860 1.795 ;
        RECT 4.700 1.725 4.890 1.805 ;
        RECT 4.710 1.725 4.890 1.815 ;
        RECT 3.825 2.460 4.860 2.630 ;
        RECT 4.690 1.705 4.870 1.795 ;
        RECT 4.690 1.715 4.880 1.795 ;
        RECT 4.720 1.725 4.890 2.629 ;
        RECT 4.690 0.535 5.485 0.705 ;
        RECT 7.880 1.645 8.050 2.630 ;
        RECT 7.910 1.245 8.080 1.815 ;
        RECT 7.880 1.645 8.080 1.815 ;
        RECT 4.890 2.460 8.720 2.630 ;
        RECT 8.550 2.460 8.720 2.760 ;
        RECT 8.905 1.325 10.170 1.495 ;
        RECT 10.000 0.890 10.170 2.215 ;
        RECT 9.655 2.045 10.170 2.215 ;
        RECT 10.000 1.540 10.580 1.840 ;
        RECT 8.185 0.870 8.515 1.040 ;
        RECT 8.345 0.870 8.515 2.215 ;
        RECT 8.345 1.675 8.530 2.215 ;
        RECT 8.230 2.045 8.530 2.215 ;
        RECT 9.010 1.675 9.180 2.590 ;
        RECT 8.345 1.675 9.685 1.845 ;
        RECT 11.200 1.610 11.370 2.590 ;
        RECT 9.010 2.420 11.370 2.590 ;
        RECT 11.200 1.610 11.380 1.910 ;
  END 
END FFSDSHDMXHT

MACRO FFSDSHDLXHT
  CLASS  CORE ;
  FOREIGN FFSDSHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.890 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.550 1.060 11.790 1.360 ;
        RECT 11.580 1.060 11.790 2.430 ;
        RECT 11.550 1.980 11.790 2.430 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.485 1.125 10.970 1.295 ;
        RECT 10.760 1.125 10.970 2.240 ;
        RECT 10.445 2.070 10.970 2.240 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.525 2.980 ;
        RECT 0.100 2.810 1.525 2.980 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.435 -0.300 2.735 0.595 ;
        RECT 3.325 -0.300 3.625 0.595 ;
        RECT 5.945 -0.300 6.245 0.745 ;
        RECT 7.165 -0.300 7.335 0.850 ;
        RECT 9.150 -0.300 9.320 0.640 ;
        RECT 10.995 -0.300 11.295 0.595 ;
        RECT 0.000 -0.300 11.890 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.760 1.525 3.250 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.560 0.520 7.730 1.910 ;
        RECT 6.885 1.610 7.730 1.910 ;
        RECT 7.560 0.520 8.905 0.690 ;
        RECT 8.735 0.520 8.905 1.145 ;
        RECT 9.595 0.540 9.765 1.145 ;
        RECT 8.735 0.920 9.765 1.145 ;
        RECT 9.595 0.540 10.005 0.710 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.565 2.715 3.215 3.990 ;
        RECT 5.855 3.160 6.155 3.990 ;
        RECT 7.100 3.160 7.400 3.990 ;
        RECT 9.075 2.770 9.375 3.990 ;
        RECT 9.720 2.810 9.890 3.990 ;
        RECT 10.995 2.770 11.295 3.990 ;
        RECT 0.000 3.390 11.890 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.525 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 2.955 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.530 0.865 1.720 1.185 ;
        RECT 1.985 0.775 2.155 1.035 ;
        RECT 1.530 0.865 2.155 1.035 ;
        RECT 1.985 0.775 4.530 0.945 ;
        RECT 4.360 0.775 4.530 2.280 ;
        RECT 5.060 0.900 5.230 2.280 ;
        RECT 5.060 1.675 6.355 1.845 ;
        RECT 6.535 1.060 6.705 2.215 ;
        RECT 6.435 2.045 6.735 2.215 ;
        RECT 6.535 1.060 7.380 1.360 ;
        RECT 2.745 1.125 3.605 1.295 ;
        RECT 2.775 2.190 3.605 2.360 ;
        RECT 3.435 1.125 3.605 2.980 ;
        RECT 3.435 1.525 3.730 1.825 ;
        RECT 3.435 2.810 8.045 2.980 ;
        RECT 3.785 1.125 4.115 1.295 ;
        RECT 3.935 1.125 4.115 2.630 ;
        RECT 3.815 2.455 4.115 2.630 ;
        RECT 4.710 0.535 4.880 2.630 ;
        RECT 4.710 0.535 5.505 0.705 ;
        RECT 7.910 1.205 8.080 2.630 ;
        RECT 3.815 2.460 8.755 2.630 ;
        RECT 10.000 1.325 10.170 2.215 ;
        RECT 9.655 2.045 10.170 2.215 ;
        RECT 10.030 0.890 10.200 1.775 ;
        RECT 8.905 1.325 10.200 1.495 ;
        RECT 10.000 1.475 10.580 1.775 ;
        RECT 8.305 0.870 8.475 2.280 ;
        RECT 8.295 1.980 8.475 2.280 ;
        RECT 8.185 0.870 8.485 1.040 ;
        RECT 9.010 1.675 9.180 2.590 ;
        RECT 8.305 1.675 9.685 1.845 ;
        RECT 11.200 1.610 11.370 2.590 ;
        RECT 9.010 2.420 11.370 2.590 ;
        RECT 11.200 1.610 11.380 1.910 ;
  END 
END FFSDSHDLXHT

MACRO FFSDSHD2XHT
  CLASS  CORE ;
  FOREIGN FFSDSHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.530 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 12.670 0.720 12.840 2.960 ;
        RECT 12.670 1.645 13.020 2.015 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.580 0.720 11.800 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.595 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.265 -0.300 2.565 0.595 ;
        RECT 3.325 -0.300 3.625 0.595 ;
        RECT 5.885 -0.300 6.185 0.905 ;
        RECT 7.375 -0.300 7.675 0.715 ;
        RECT 9.540 -0.300 9.840 0.740 ;
        RECT 11.045 -0.300 11.345 1.055 ;
        RECT 12.085 -0.300 12.385 1.055 ;
        RECT 13.125 -0.300 13.425 1.055 ;
        RECT 0.000 -0.300 13.530 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.730 1.525 3.220 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.265 0.960 7.435 1.565 ;
        RECT 7.160 1.265 7.435 1.565 ;
        RECT 7.855 0.605 8.025 1.130 ;
        RECT 7.265 0.960 8.025 1.130 ;
        RECT 7.855 0.605 9.185 0.775 ;
        RECT 9.015 0.605 9.185 1.145 ;
        RECT 9.875 0.920 10.420 1.145 ;
        RECT 10.250 0.515 10.420 1.145 ;
        RECT 9.015 0.975 10.420 1.145 ;
        RECT 10.250 0.515 10.580 0.685 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.585 2.830 3.225 3.990 ;
        RECT 5.855 3.095 6.155 3.990 ;
        RECT 7.005 3.095 7.645 3.990 ;
        RECT 9.425 2.790 9.725 3.990 ;
        RECT 10.535 2.790 10.835 3.990 ;
        RECT 11.045 2.975 11.345 3.990 ;
        RECT 12.085 2.975 12.385 3.990 ;
        RECT 13.125 2.295 13.425 3.990 ;
        RECT 0.000 3.390 13.530 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.575 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.150 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.950 0.775 2.120 1.035 ;
        RECT 1.530 0.865 2.120 1.035 ;
        RECT 1.950 0.775 4.500 0.945 ;
        RECT 4.330 0.775 4.500 2.280 ;
        RECT 5.030 0.910 5.200 2.280 ;
        RECT 6.105 1.675 6.405 1.865 ;
        RECT 5.030 1.695 6.405 1.865 ;
        RECT 5.625 1.245 5.925 1.515 ;
        RECT 5.625 1.245 6.980 1.415 ;
        RECT 6.810 0.670 6.980 2.215 ;
        RECT 6.405 2.045 6.980 2.215 ;
        RECT 6.810 0.670 7.030 0.970 ;
        RECT 7.655 1.610 7.825 1.915 ;
        RECT 6.810 1.745 7.825 1.915 ;
        RECT 2.775 1.125 3.575 1.295 ;
        RECT 2.775 2.190 3.575 2.360 ;
        RECT 3.405 1.125 3.575 3.055 ;
        RECT 3.405 1.525 3.700 1.825 ;
        RECT 3.405 2.885 5.505 3.055 ;
        RECT 5.765 2.745 8.470 2.915 ;
        RECT 8.290 2.745 8.470 3.185 ;
        RECT 8.290 3.015 8.910 3.185 ;
        RECT 5.645 2.745 5.655 3.025 ;
        RECT 5.655 2.745 5.665 3.015 ;
        RECT 5.665 2.745 5.675 3.005 ;
        RECT 5.675 2.745 5.685 2.995 ;
        RECT 5.685 2.745 5.695 2.985 ;
        RECT 5.695 2.745 5.705 2.975 ;
        RECT 5.705 2.745 5.715 2.965 ;
        RECT 5.715 2.745 5.725 2.955 ;
        RECT 5.725 2.745 5.735 2.945 ;
        RECT 5.735 2.745 5.745 2.935 ;
        RECT 5.745 2.745 5.755 2.925 ;
        RECT 5.755 2.745 5.765 2.915 ;
        RECT 5.625 2.765 5.635 3.045 ;
        RECT 5.635 2.755 5.645 3.035 ;
        RECT 5.505 2.885 5.515 3.055 ;
        RECT 5.515 2.875 5.525 3.055 ;
        RECT 5.525 2.865 5.535 3.055 ;
        RECT 5.535 2.855 5.545 3.055 ;
        RECT 5.545 2.845 5.555 3.055 ;
        RECT 5.555 2.835 5.565 3.055 ;
        RECT 5.565 2.825 5.575 3.055 ;
        RECT 5.575 2.815 5.585 3.055 ;
        RECT 5.585 2.805 5.595 3.055 ;
        RECT 5.595 2.795 5.605 3.055 ;
        RECT 5.605 2.785 5.615 3.055 ;
        RECT 5.615 2.775 5.625 3.055 ;
        RECT 3.755 1.125 4.075 1.295 ;
        RECT 3.905 1.125 4.075 2.635 ;
        RECT 3.820 1.980 4.075 2.635 ;
        RECT 4.680 0.535 4.850 2.700 ;
        RECT 4.595 2.465 4.895 2.700 ;
        RECT 5.355 2.425 5.435 2.635 ;
        RECT 5.345 2.435 9.000 2.565 ;
        RECT 5.365 2.415 5.435 2.635 ;
        RECT 5.335 2.445 9.000 2.565 ;
        RECT 5.375 2.405 5.435 2.635 ;
        RECT 5.325 2.455 9.000 2.565 ;
        RECT 3.820 2.465 5.435 2.635 ;
        RECT 4.680 0.535 5.445 0.705 ;
        RECT 3.820 2.465 5.445 2.625 ;
        RECT 3.820 2.465 5.455 2.615 ;
        RECT 3.820 2.465 5.465 2.605 ;
        RECT 3.820 2.465 5.475 2.595 ;
        RECT 3.820 2.465 5.485 2.585 ;
        RECT 3.820 2.465 5.495 2.575 ;
        RECT 8.135 1.290 8.305 2.565 ;
        RECT 5.385 2.395 9.000 2.565 ;
        RECT 8.830 2.395 9.000 2.770 ;
        RECT 9.235 1.325 10.770 1.495 ;
        RECT 10.600 1.060 10.770 2.215 ;
        RECT 9.985 2.045 10.770 2.215 ;
        RECT 10.600 1.675 11.400 1.845 ;
        RECT 8.580 0.955 8.795 2.215 ;
        RECT 8.535 0.955 8.835 1.125 ;
        RECT 8.560 2.045 8.860 2.215 ;
        RECT 9.635 1.675 9.805 2.610 ;
        RECT 8.580 1.675 10.050 1.845 ;
        RECT 11.030 2.440 11.275 2.630 ;
        RECT 9.635 2.440 11.275 2.610 ;
        RECT 12.320 1.610 12.490 2.630 ;
        RECT 11.030 2.460 12.490 2.630 ;
  END 
END FFSDSHD2XHT

MACRO FFSDSHD1XHT
  CLASS  CORE ;
  FOREIGN FFSDSHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.890 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.550 0.720 11.790 1.360 ;
        RECT 11.580 0.720 11.790 2.960 ;
        RECT 11.550 1.980 11.790 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.510 0.720 10.680 1.360 ;
        RECT 10.510 1.190 10.970 1.360 ;
        RECT 10.760 1.190 10.970 2.240 ;
        RECT 10.445 2.070 10.970 2.240 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.385 -0.300 2.685 0.595 ;
        RECT 3.335 -0.300 3.635 0.595 ;
        RECT 6.760 -0.300 7.335 0.780 ;
        RECT 9.150 -0.300 9.320 0.590 ;
        RECT 10.965 -0.300 11.265 0.715 ;
        RECT 0.000 -0.300 11.890 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.740 1.525 3.230 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.435 1.800 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.530 0.605 7.700 1.910 ;
        RECT 6.885 1.610 7.700 1.910 ;
        RECT 7.530 0.605 8.905 0.775 ;
        RECT 8.735 0.605 8.905 1.145 ;
        RECT 9.595 0.520 9.765 1.145 ;
        RECT 8.735 0.920 9.765 1.145 ;
        RECT 9.595 0.520 10.055 0.690 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.585 2.740 3.225 3.990 ;
        RECT 5.855 3.160 6.155 3.990 ;
        RECT 7.100 3.160 7.400 3.990 ;
        RECT 9.105 3.035 10.105 3.990 ;
        RECT 10.965 2.975 11.265 3.990 ;
        RECT 0.000 3.390 11.890 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.575 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.150 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.955 0.775 2.125 1.035 ;
        RECT 1.530 0.865 2.125 1.035 ;
        RECT 1.955 0.775 4.510 0.945 ;
        RECT 4.340 0.775 4.510 2.280 ;
        RECT 5.040 0.900 5.210 2.280 ;
        RECT 5.040 1.605 6.355 1.775 ;
        RECT 6.535 1.060 6.705 2.215 ;
        RECT 6.405 2.045 6.705 2.215 ;
        RECT 6.535 1.060 7.350 1.360 ;
        RECT 2.785 1.125 3.585 1.295 ;
        RECT 2.785 2.190 3.585 2.360 ;
        RECT 3.415 1.125 3.585 2.980 ;
        RECT 3.415 1.525 3.710 1.825 ;
        RECT 3.415 2.810 8.205 2.980 ;
        RECT 3.765 1.125 4.085 1.295 ;
        RECT 3.830 1.980 4.085 2.280 ;
        RECT 3.915 1.125 4.085 2.630 ;
        RECT 4.690 0.535 4.860 2.630 ;
        RECT 4.690 0.535 5.485 0.705 ;
        RECT 7.880 1.645 8.050 2.630 ;
        RECT 7.910 1.245 8.080 1.815 ;
        RECT 7.880 1.645 8.080 1.815 ;
        RECT 3.915 2.460 8.720 2.630 ;
        RECT 8.550 2.460 8.720 2.770 ;
        RECT 8.905 1.325 10.240 1.495 ;
        RECT 10.000 0.890 10.170 1.495 ;
        RECT 10.070 1.325 10.240 2.215 ;
        RECT 9.655 2.045 10.240 2.215 ;
        RECT 10.070 1.540 10.580 1.840 ;
        RECT 8.215 0.955 8.515 1.125 ;
        RECT 8.345 0.955 8.515 2.215 ;
        RECT 8.345 1.675 8.530 2.215 ;
        RECT 8.230 2.045 8.530 2.215 ;
        RECT 9.010 1.675 9.180 2.590 ;
        RECT 8.345 1.675 9.685 1.845 ;
        RECT 11.200 1.610 11.370 2.590 ;
        RECT 9.010 2.420 11.370 2.590 ;
        RECT 11.200 1.610 11.380 1.910 ;
  END 
END FFSDSHD1XHT

MACRO FFSDRHQHDMXHT
  CLASS  CORE ;
  FOREIGN FFSDRHQHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.940 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.545 1.060 13.845 2.455 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.270 1.280 1.775 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 11.075 0.920 11.510 1.350 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.615 0.380 2.115 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.085 ;
        RECT 2.545 -0.300 2.845 0.595 ;
        RECT 3.555 -0.300 3.855 0.595 ;
        RECT 4.495 -0.300 4.795 0.595 ;
        RECT 7.500 -0.300 7.800 0.595 ;
        RECT 8.990 -0.300 9.290 0.990 ;
        RECT 10.960 -0.300 11.260 0.740 ;
        RECT 12.060 -0.300 12.360 0.535 ;
        RECT 12.995 -0.300 13.165 0.780 ;
        RECT 0.000 -0.300 13.940 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 4.495 1.605 5.010 2.020 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.235 1.530 2.785 2.020 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.655 0.955 3.990 ;
        RECT 2.555 2.470 2.730 3.990 ;
        RECT 3.555 2.745 3.855 3.990 ;
        RECT 4.375 2.745 4.675 3.990 ;
        RECT 7.515 2.885 7.815 3.990 ;
        RECT 8.995 3.095 9.295 3.990 ;
        RECT 10.880 3.095 11.180 3.990 ;
        RECT 12.995 2.650 13.165 3.990 ;
        RECT 0.000 3.390 13.940 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.010 0.340 1.435 ;
        RECT 0.170 1.265 0.730 1.435 ;
        RECT 0.560 1.265 0.730 2.465 ;
        RECT 0.105 2.295 0.730 2.465 ;
        RECT 1.460 1.510 1.630 2.125 ;
        RECT 0.560 1.955 1.630 2.125 ;
        RECT 3.390 1.600 3.560 1.905 ;
        RECT 3.390 1.600 4.285 1.780 ;
        RECT 3.985 1.125 4.285 2.215 ;
        RECT 5.045 1.125 5.705 1.295 ;
        RECT 5.535 1.125 5.705 2.215 ;
        RECT 5.295 2.045 5.705 2.215 ;
        RECT 1.640 1.070 1.980 1.260 ;
        RECT 1.640 0.960 1.810 1.260 ;
        RECT 1.640 2.330 1.810 2.970 ;
        RECT 1.810 1.070 1.980 2.560 ;
        RECT 1.640 2.330 1.980 2.560 ;
        RECT 2.485 0.775 2.655 1.240 ;
        RECT 1.640 1.070 2.655 1.240 ;
        RECT 2.485 0.775 6.180 0.945 ;
        RECT 6.010 0.775 6.180 2.320 ;
        RECT 6.710 1.060 6.880 2.355 ;
        RECT 7.785 1.585 7.955 2.210 ;
        RECT 6.710 2.040 7.955 2.210 ;
        RECT 7.785 1.585 8.085 1.755 ;
        RECT 7.370 1.220 7.540 1.820 ;
        RECT 8.070 1.125 8.435 1.390 ;
        RECT 7.370 1.220 8.435 1.390 ;
        RECT 8.265 1.125 8.435 2.215 ;
        RECT 8.265 2.045 8.815 2.215 ;
        RECT 8.265 1.525 9.180 1.825 ;
        RECT 3.005 1.125 3.185 2.565 ;
        RECT 3.005 2.100 3.240 2.565 ;
        RECT 3.005 1.125 3.305 1.295 ;
        RECT 5.115 2.395 5.415 2.670 ;
        RECT 3.005 2.395 5.415 2.565 ;
        RECT 6.360 0.650 6.530 2.670 ;
        RECT 5.115 2.500 6.530 2.670 ;
        RECT 7.110 0.650 7.280 0.945 ;
        RECT 6.360 0.650 7.280 0.830 ;
        RECT 7.110 0.775 8.785 0.945 ;
        RECT 8.615 0.775 8.785 1.345 ;
        RECT 8.615 1.175 9.925 1.345 ;
        RECT 9.755 1.175 9.925 1.610 ;
        RECT 7.675 2.395 7.845 2.705 ;
        RECT 6.825 2.535 7.845 2.705 ;
        RECT 7.675 2.395 9.535 2.565 ;
        RECT 9.365 1.925 9.535 2.565 ;
        RECT 10.125 0.920 10.295 2.095 ;
        RECT 9.365 1.925 10.295 2.095 ;
        RECT 10.125 0.920 10.430 1.220 ;
        RECT 8.650 2.745 8.820 3.045 ;
        RECT 8.310 2.875 8.820 3.045 ;
        RECT 8.650 2.745 11.765 2.915 ;
        RECT 11.430 2.480 11.730 2.915 ;
        RECT 11.430 2.535 11.765 2.915 ;
        RECT 11.430 2.535 12.535 2.705 ;
        RECT 11.490 0.570 11.860 0.740 ;
        RECT 11.690 0.570 11.860 0.925 ;
        RECT 11.690 0.755 12.620 0.925 ;
        RECT 9.950 0.570 10.780 0.740 ;
        RECT 10.475 1.550 10.645 2.565 ;
        RECT 9.915 2.395 10.645 2.565 ;
        RECT 10.610 0.570 10.780 1.720 ;
        RECT 10.475 1.550 12.950 1.720 ;
        RECT 10.825 1.925 11.075 2.225 ;
        RECT 12.495 1.125 13.335 1.295 ;
        RECT 13.145 1.125 13.335 2.225 ;
        RECT 10.825 2.055 13.335 2.225 ;
  END 
END FFSDRHQHDMXHT

MACRO FFSDRHQHD3XHT
  CLASS  CORE ;
  FOREIGN FFSDRHQHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.220 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 15.840 0.480 16.010 1.130 ;
        RECT 15.840 2.405 16.010 3.045 ;
        RECT 15.840 0.960 17.125 1.130 ;
        RECT 16.760 0.960 17.125 2.705 ;
        RECT 15.840 2.405 17.125 2.705 ;
        RECT 16.815 0.720 17.125 2.895 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.240 1.165 1.775 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 13.885 1.465 14.315 1.965 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.545 0.380 2.020 ;
        RECT 0.250 0.755 0.550 0.945 ;
        RECT 1.165 0.485 1.335 0.945 ;
        RECT 0.250 0.775 1.335 0.945 ;
        RECT 1.165 0.485 2.155 0.655 ;
        RECT 0.285 2.580 0.470 2.840 ;
        RECT 0.170 2.670 0.470 2.840 ;
        RECT 0.285 2.580 1.340 2.750 ;
        RECT 0.170 2.670 1.340 2.750 ;
        RECT 1.170 2.580 1.340 3.180 ;
        RECT 1.170 3.010 2.245 3.180 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.595 ;
        RECT 2.550 -0.300 2.850 0.595 ;
        RECT 3.475 -0.300 3.775 0.595 ;
        RECT 4.415 -0.300 4.715 0.485 ;
        RECT 5.515 -0.300 5.815 0.595 ;
        RECT 7.545 -0.300 7.845 0.595 ;
        RECT 8.750 -0.300 9.390 0.595 ;
        RECT 11.075 -0.300 11.375 0.595 ;
        RECT 13.400 -0.300 13.570 0.800 ;
        RECT 14.365 -0.300 14.665 0.510 ;
        RECT 15.320 -0.300 15.490 0.780 ;
        RECT 16.360 -0.300 16.530 0.780 ;
        RECT 0.000 -0.300 17.220 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 4.550 1.605 5.305 2.020 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.145 1.530 2.505 2.020 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.975 0.955 3.990 ;
        RECT 2.555 2.830 2.730 3.990 ;
        RECT 3.670 2.830 3.840 3.990 ;
        RECT 4.435 2.875 4.735 3.990 ;
        RECT 7.475 2.880 7.775 3.990 ;
        RECT 9.395 3.075 9.565 3.990 ;
        RECT 11.135 2.975 11.435 3.990 ;
        RECT 13.290 2.885 13.590 3.990 ;
        RECT 15.320 2.910 15.490 3.990 ;
        RECT 16.360 2.910 16.530 3.990 ;
        RECT 0.000 3.390 17.220 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 0.730 1.295 ;
        RECT 0.560 1.125 0.730 2.400 ;
        RECT 0.105 2.230 0.730 2.400 ;
        RECT 1.355 1.460 1.525 2.125 ;
        RECT 0.560 1.955 1.525 2.125 ;
        RECT 1.355 1.460 1.965 1.760 ;
        RECT 3.430 1.605 3.600 1.905 ;
        RECT 3.430 1.605 4.325 1.780 ;
        RECT 4.025 1.125 4.325 2.215 ;
        RECT 4.965 1.125 5.760 1.295 ;
        RECT 5.590 1.125 5.760 2.370 ;
        RECT 5.355 2.200 5.760 2.370 ;
        RECT 1.575 2.305 1.875 2.815 ;
        RECT 1.575 0.930 2.855 1.110 ;
        RECT 2.685 0.775 2.855 2.475 ;
        RECT 1.575 2.305 2.855 2.475 ;
        RECT 2.685 0.775 6.140 0.945 ;
        RECT 5.970 0.775 6.140 2.415 ;
        RECT 6.670 1.060 6.840 2.400 ;
        RECT 7.750 1.515 7.920 2.210 ;
        RECT 6.670 2.040 7.920 2.210 ;
        RECT 7.750 1.515 8.050 1.685 ;
        RECT 7.335 1.125 7.505 1.820 ;
        RECT 7.335 1.125 8.720 1.295 ;
        RECT 8.550 1.125 8.720 2.215 ;
        RECT 8.410 2.045 8.720 2.215 ;
        RECT 9.865 1.305 10.035 1.645 ;
        RECT 8.550 1.305 10.035 1.475 ;
        RECT 9.865 1.475 11.400 1.645 ;
        RECT 3.045 1.125 3.225 2.680 ;
        RECT 3.045 2.040 3.280 2.680 ;
        RECT 3.045 1.125 3.345 1.295 ;
        RECT 3.045 2.430 5.125 2.600 ;
        RECT 4.955 2.430 5.125 3.145 ;
        RECT 4.955 2.885 5.475 3.145 ;
        RECT 6.320 0.550 6.490 3.145 ;
        RECT 4.955 2.975 6.490 3.145 ;
        RECT 6.320 0.550 7.180 0.730 ;
        RECT 7.010 0.550 7.180 0.945 ;
        RECT 9.690 0.565 9.860 1.085 ;
        RECT 7.010 0.775 9.860 0.945 ;
        RECT 9.635 0.915 10.470 1.085 ;
        RECT 10.300 0.915 10.470 1.295 ;
        RECT 10.300 1.125 12.075 1.295 ;
        RECT 11.905 1.125 12.075 1.520 ;
        RECT 11.905 1.350 12.510 1.520 ;
        RECT 12.340 1.350 12.510 1.650 ;
        RECT 7.020 2.530 7.190 2.810 ;
        RECT 6.835 2.640 7.190 2.810 ;
        RECT 7.020 2.530 9.505 2.700 ;
        RECT 9.890 2.885 10.245 3.055 ;
        RECT 9.945 2.885 10.245 3.140 ;
        RECT 11.795 1.735 12.095 2.000 ;
        RECT 12.690 0.870 12.860 2.000 ;
        RECT 9.675 1.830 12.860 2.000 ;
        RECT 9.810 2.815 9.820 3.055 ;
        RECT 9.820 2.825 9.830 3.055 ;
        RECT 9.830 2.835 9.840 3.055 ;
        RECT 9.840 2.845 9.850 3.055 ;
        RECT 9.850 2.855 9.860 3.055 ;
        RECT 9.860 2.865 9.870 3.055 ;
        RECT 9.870 2.875 9.880 3.055 ;
        RECT 9.880 2.885 9.890 3.055 ;
        RECT 9.675 2.680 9.685 2.920 ;
        RECT 9.685 2.690 9.695 2.930 ;
        RECT 9.695 2.700 9.705 2.940 ;
        RECT 9.705 2.710 9.715 2.950 ;
        RECT 9.715 2.720 9.725 2.960 ;
        RECT 9.725 2.730 9.735 2.970 ;
        RECT 9.735 2.740 9.745 2.980 ;
        RECT 9.745 2.750 9.755 2.990 ;
        RECT 9.755 2.760 9.765 3.000 ;
        RECT 9.765 2.770 9.775 3.010 ;
        RECT 9.775 2.780 9.785 3.020 ;
        RECT 9.785 2.790 9.795 3.030 ;
        RECT 9.795 2.800 9.805 3.040 ;
        RECT 9.805 2.805 9.811 3.049 ;
        RECT 9.505 1.830 9.515 2.750 ;
        RECT 9.515 1.830 9.525 2.760 ;
        RECT 9.525 1.830 9.535 2.770 ;
        RECT 9.535 1.830 9.545 2.780 ;
        RECT 9.545 1.830 9.555 2.790 ;
        RECT 9.555 1.830 9.565 2.800 ;
        RECT 9.565 1.830 9.575 2.810 ;
        RECT 9.575 1.830 9.585 2.820 ;
        RECT 9.585 1.830 9.595 2.830 ;
        RECT 9.595 1.830 9.605 2.840 ;
        RECT 9.605 1.830 9.615 2.850 ;
        RECT 9.615 1.830 9.625 2.860 ;
        RECT 9.625 1.830 9.635 2.870 ;
        RECT 9.635 1.830 9.645 2.880 ;
        RECT 9.645 1.830 9.655 2.890 ;
        RECT 9.655 1.830 9.665 2.900 ;
        RECT 9.665 1.830 9.675 2.910 ;
        RECT 9.990 2.205 10.025 2.700 ;
        RECT 10.080 2.530 11.795 2.700 ;
        RECT 11.625 2.530 11.795 3.100 ;
        RECT 12.605 2.535 12.775 3.100 ;
        RECT 11.625 2.930 12.775 3.100 ;
        RECT 12.605 2.535 14.905 2.705 ;
        RECT 10.025 2.485 10.035 2.699 ;
        RECT 10.035 2.495 10.045 2.699 ;
        RECT 10.045 2.505 10.055 2.699 ;
        RECT 10.055 2.515 10.065 2.699 ;
        RECT 10.065 2.525 10.075 2.699 ;
        RECT 10.075 2.530 10.081 2.700 ;
        RECT 9.855 2.205 9.865 2.565 ;
        RECT 9.865 2.205 9.875 2.575 ;
        RECT 9.875 2.205 9.885 2.585 ;
        RECT 9.885 2.205 9.895 2.595 ;
        RECT 9.895 2.205 9.905 2.605 ;
        RECT 9.905 2.205 9.915 2.615 ;
        RECT 9.915 2.205 9.925 2.625 ;
        RECT 9.925 2.205 9.935 2.635 ;
        RECT 9.935 2.205 9.945 2.645 ;
        RECT 9.945 2.205 9.955 2.655 ;
        RECT 9.955 2.205 9.965 2.665 ;
        RECT 9.965 2.205 9.975 2.675 ;
        RECT 9.975 2.205 9.985 2.685 ;
        RECT 9.985 2.205 9.991 2.695 ;
        RECT 13.855 0.710 14.915 0.880 ;
        RECT 10.045 0.545 10.880 0.715 ;
        RECT 10.710 0.545 10.880 0.945 ;
        RECT 10.710 0.775 12.440 0.945 ;
        RECT 12.075 2.180 12.375 2.695 ;
        RECT 12.270 0.480 12.440 1.120 ;
        RECT 12.270 0.480 13.210 0.650 ;
        RECT 13.040 0.480 13.210 2.350 ;
        RECT 10.225 2.180 13.210 2.350 ;
        RECT 13.040 1.095 14.680 1.265 ;
        RECT 14.510 1.095 14.680 1.830 ;
        RECT 14.510 1.660 16.130 1.830 ;
        RECT 13.410 1.445 13.580 2.350 ;
        RECT 14.860 1.060 15.030 1.360 ;
        RECT 14.905 2.025 15.075 2.350 ;
        RECT 13.410 2.155 15.075 2.350 ;
        RECT 14.860 1.125 15.515 1.295 ;
        RECT 15.345 1.125 15.515 1.480 ;
        RECT 15.345 1.310 16.530 1.480 ;
        RECT 14.905 2.025 16.530 2.200 ;
        RECT 16.360 1.310 16.530 2.200 ;
  END 
END FFSDRHQHD3XHT

MACRO FFSDRHQHD2XHT
  CLASS  CORE ;
  FOREIGN FFSDRHQHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.990 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 15.075 0.720 15.245 2.960 ;
        RECT 15.075 1.660 15.480 2.035 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.090 1.135 1.775 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 12.545 0.915 13.080 1.340 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.545 0.380 2.020 ;
        RECT 0.300 2.580 0.485 2.840 ;
        RECT 0.185 2.670 0.485 2.840 ;
        RECT 0.300 2.580 1.340 2.750 ;
        RECT 0.185 2.670 1.340 2.750 ;
        RECT 1.170 2.580 1.340 3.180 ;
        RECT 1.170 3.010 2.245 3.180 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.900 ;
        RECT 2.545 -0.300 2.845 0.595 ;
        RECT 3.455 -0.300 3.755 0.595 ;
        RECT 4.515 -0.300 4.815 0.595 ;
        RECT 7.605 -0.300 7.905 0.585 ;
        RECT 8.870 -0.300 9.170 0.585 ;
        RECT 10.580 -0.300 10.880 0.665 ;
        RECT 12.545 -0.300 12.845 0.725 ;
        RECT 13.620 -0.300 13.920 0.545 ;
        RECT 14.555 -0.300 14.725 0.780 ;
        RECT 15.595 -0.300 15.765 1.120 ;
        RECT 0.000 -0.300 15.990 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 4.525 1.560 5.040 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.145 1.550 2.500 2.010 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.945 0.955 3.990 ;
        RECT 2.555 2.850 2.730 3.990 ;
        RECT 3.585 2.760 3.885 3.990 ;
        RECT 4.395 2.760 4.705 3.990 ;
        RECT 7.375 2.830 7.680 3.990 ;
        RECT 9.220 3.170 9.540 3.990 ;
        RECT 10.580 3.085 10.885 3.990 ;
        RECT 12.445 3.085 12.745 3.990 ;
        RECT 14.555 2.910 14.725 3.990 ;
        RECT 15.595 2.220 15.765 3.990 ;
        RECT 0.000 3.390 15.990 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.085 0.730 1.255 ;
        RECT 0.560 1.085 0.730 2.400 ;
        RECT 0.105 2.230 0.730 2.400 ;
        RECT 1.795 1.460 1.965 2.125 ;
        RECT 0.560 1.955 1.965 2.125 ;
        RECT 3.410 1.595 3.580 1.895 ;
        RECT 3.410 1.595 4.305 1.770 ;
        RECT 4.005 1.125 4.305 2.215 ;
        RECT 5.065 1.125 5.695 1.295 ;
        RECT 5.525 1.125 5.695 2.215 ;
        RECT 5.315 2.045 5.695 2.215 ;
        RECT 1.575 2.305 1.875 2.815 ;
        RECT 2.425 0.775 2.435 1.005 ;
        RECT 1.575 0.825 2.435 1.005 ;
        RECT 1.575 2.305 2.510 2.475 ;
        RECT 2.605 0.775 6.060 0.945 ;
        RECT 5.890 0.775 6.060 2.405 ;
        RECT 2.685 1.235 2.695 2.375 ;
        RECT 2.695 1.245 2.705 2.365 ;
        RECT 2.705 1.255 2.715 2.355 ;
        RECT 2.715 1.265 2.725 2.345 ;
        RECT 2.725 1.275 2.735 2.335 ;
        RECT 2.735 1.285 2.745 2.325 ;
        RECT 2.745 1.295 2.755 2.315 ;
        RECT 2.755 1.305 2.765 2.305 ;
        RECT 2.765 1.315 2.775 2.295 ;
        RECT 2.775 1.325 2.785 2.285 ;
        RECT 2.785 1.335 2.795 2.275 ;
        RECT 2.795 1.345 2.805 2.265 ;
        RECT 2.805 1.355 2.815 2.255 ;
        RECT 2.815 1.365 2.825 2.245 ;
        RECT 2.825 1.375 2.835 2.235 ;
        RECT 2.835 1.385 2.845 2.225 ;
        RECT 2.845 1.395 2.855 2.215 ;
        RECT 2.605 1.155 2.615 1.395 ;
        RECT 2.615 1.165 2.625 1.405 ;
        RECT 2.625 1.175 2.635 1.415 ;
        RECT 2.635 1.185 2.645 1.425 ;
        RECT 2.645 1.195 2.655 1.435 ;
        RECT 2.655 1.205 2.665 1.445 ;
        RECT 2.665 1.215 2.675 1.455 ;
        RECT 2.675 1.225 2.685 1.465 ;
        RECT 2.595 2.220 2.605 2.464 ;
        RECT 2.605 2.210 2.615 2.454 ;
        RECT 2.615 2.200 2.625 2.444 ;
        RECT 2.625 2.190 2.635 2.434 ;
        RECT 2.635 2.180 2.645 2.424 ;
        RECT 2.645 2.170 2.655 2.414 ;
        RECT 2.655 2.160 2.665 2.404 ;
        RECT 2.665 2.150 2.675 2.394 ;
        RECT 2.675 2.140 2.685 2.384 ;
        RECT 2.435 0.775 2.445 1.225 ;
        RECT 2.445 0.775 2.455 1.235 ;
        RECT 2.455 0.775 2.465 1.245 ;
        RECT 2.465 0.775 2.475 1.255 ;
        RECT 2.475 0.775 2.485 1.265 ;
        RECT 2.485 0.775 2.495 1.275 ;
        RECT 2.495 0.775 2.505 1.285 ;
        RECT 2.505 0.775 2.515 1.295 ;
        RECT 2.515 0.775 2.525 1.305 ;
        RECT 2.525 0.775 2.535 1.315 ;
        RECT 2.535 0.775 2.545 1.325 ;
        RECT 2.545 0.775 2.555 1.335 ;
        RECT 2.555 0.775 2.565 1.345 ;
        RECT 2.565 0.775 2.575 1.355 ;
        RECT 2.575 0.775 2.585 1.365 ;
        RECT 2.585 0.775 2.595 1.375 ;
        RECT 2.595 0.775 2.605 1.385 ;
        RECT 2.510 2.305 2.520 2.475 ;
        RECT 2.520 2.295 2.530 2.475 ;
        RECT 2.530 2.285 2.540 2.475 ;
        RECT 2.540 2.275 2.550 2.475 ;
        RECT 2.550 2.265 2.560 2.475 ;
        RECT 2.560 2.255 2.570 2.475 ;
        RECT 2.570 2.245 2.580 2.475 ;
        RECT 2.580 2.235 2.590 2.475 ;
        RECT 2.590 2.225 2.596 2.475 ;
        RECT 6.590 1.050 6.760 2.355 ;
        RECT 7.695 1.485 7.865 2.200 ;
        RECT 6.590 2.030 7.865 2.200 ;
        RECT 7.695 1.485 7.995 1.655 ;
        RECT 7.280 1.115 7.450 1.810 ;
        RECT 8.365 1.115 8.535 2.290 ;
        RECT 7.280 1.115 8.600 1.285 ;
        RECT 8.300 2.120 8.600 2.290 ;
        RECT 8.365 1.560 10.855 1.730 ;
        RECT 3.060 1.125 3.230 2.880 ;
        RECT 3.025 1.125 3.325 1.295 ;
        RECT 3.025 2.305 3.325 2.880 ;
        RECT 3.025 2.395 5.435 2.565 ;
        RECT 5.135 2.395 5.435 2.860 ;
        RECT 6.240 0.540 6.410 2.860 ;
        RECT 5.135 2.690 6.410 2.860 ;
        RECT 6.240 0.540 7.255 0.720 ;
        RECT 7.085 0.540 7.255 0.935 ;
        RECT 7.085 0.765 8.685 0.935 ;
        RECT 8.970 0.950 9.040 1.365 ;
        RECT 8.970 1.195 11.505 1.365 ;
        RECT 11.335 1.195 11.505 1.685 ;
        RECT 8.870 0.860 8.880 1.364 ;
        RECT 8.880 0.870 8.890 1.364 ;
        RECT 8.890 0.880 8.900 1.364 ;
        RECT 8.900 0.890 8.910 1.364 ;
        RECT 8.910 0.900 8.920 1.364 ;
        RECT 8.920 0.910 8.930 1.364 ;
        RECT 8.930 0.920 8.940 1.364 ;
        RECT 8.940 0.930 8.950 1.364 ;
        RECT 8.950 0.940 8.960 1.364 ;
        RECT 8.960 0.950 8.970 1.364 ;
        RECT 8.785 0.775 8.795 1.035 ;
        RECT 8.795 0.785 8.805 1.045 ;
        RECT 8.805 0.795 8.815 1.055 ;
        RECT 8.815 0.805 8.825 1.065 ;
        RECT 8.825 0.815 8.835 1.075 ;
        RECT 8.835 0.825 8.845 1.085 ;
        RECT 8.845 0.835 8.855 1.095 ;
        RECT 8.855 0.845 8.865 1.105 ;
        RECT 8.865 0.850 8.871 1.114 ;
        RECT 8.685 0.765 8.695 0.935 ;
        RECT 8.695 0.765 8.705 0.945 ;
        RECT 8.705 0.765 8.715 0.955 ;
        RECT 8.715 0.765 8.725 0.965 ;
        RECT 8.725 0.765 8.735 0.975 ;
        RECT 8.735 0.765 8.745 0.985 ;
        RECT 8.745 0.765 8.755 0.995 ;
        RECT 8.755 0.765 8.765 1.005 ;
        RECT 8.765 0.765 8.775 1.015 ;
        RECT 8.775 0.765 8.785 1.025 ;
        RECT 6.940 2.470 7.110 2.780 ;
        RECT 6.730 2.610 7.110 2.780 ;
        RECT 6.940 2.470 8.950 2.640 ;
        RECT 8.780 1.930 8.950 2.640 ;
        RECT 11.685 1.065 11.855 2.100 ;
        RECT 8.780 1.930 11.855 2.100 ;
        RECT 11.685 1.065 12.015 1.365 ;
        RECT 8.360 2.820 8.530 3.120 ;
        RECT 9.120 2.735 9.290 2.990 ;
        RECT 8.360 2.820 9.290 2.990 ;
        RECT 9.120 2.735 13.175 2.905 ;
        RECT 13.000 2.570 13.175 2.905 ;
        RECT 13.000 2.570 14.085 2.740 ;
        RECT 13.065 0.555 13.440 0.725 ;
        RECT 13.270 0.555 13.440 0.915 ;
        RECT 13.270 0.745 14.150 0.915 ;
        RECT 11.335 0.715 11.505 1.015 ;
        RECT 9.595 0.845 11.505 1.015 ;
        RECT 11.335 0.715 12.365 0.885 ;
        RECT 12.055 1.545 12.225 2.520 ;
        RECT 9.655 2.350 12.225 2.520 ;
        RECT 12.195 0.715 12.365 1.715 ;
        RECT 12.055 1.545 14.475 1.715 ;
        RECT 12.405 1.915 12.575 2.215 ;
        RECT 13.510 2.045 13.810 2.285 ;
        RECT 14.030 1.125 14.845 1.295 ;
        RECT 14.655 1.125 14.845 2.215 ;
        RECT 12.405 2.045 14.845 2.215 ;
  END 
END FFSDRHQHD2XHT

MACRO FFSDRHQHD1XHT
  CLASS  CORE ;
  FOREIGN FFSDRHQHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.940 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.545 0.720 13.845 2.965 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.225 1.165 1.775 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 11.100 0.920 11.515 1.350 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.575 0.380 2.020 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.045 ;
        RECT 2.545 -0.300 2.845 0.595 ;
        RECT 3.525 -0.300 3.825 0.595 ;
        RECT 4.495 -0.300 4.795 0.595 ;
        RECT 7.585 -0.300 7.885 0.470 ;
        RECT 8.960 -0.300 9.260 0.470 ;
        RECT 10.960 -0.300 11.260 0.740 ;
        RECT 12.055 -0.300 12.355 0.515 ;
        RECT 13.025 -0.300 13.195 0.780 ;
        RECT 0.000 -0.300 13.940 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 4.495 1.535 5.010 2.020 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.235 1.530 2.785 2.020 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.655 0.955 3.990 ;
        RECT 2.555 2.470 2.730 3.990 ;
        RECT 3.555 2.745 3.855 3.990 ;
        RECT 4.375 2.745 4.675 3.990 ;
        RECT 7.515 2.745 7.815 3.990 ;
        RECT 8.995 3.095 9.295 3.990 ;
        RECT 10.880 3.095 11.180 3.990 ;
        RECT 13.025 2.910 13.195 3.990 ;
        RECT 0.000 3.390 13.940 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.010 0.340 1.395 ;
        RECT 0.170 2.220 0.340 2.520 ;
        RECT 0.170 1.225 0.730 1.395 ;
        RECT 0.560 1.225 0.730 2.390 ;
        RECT 0.170 2.220 0.730 2.390 ;
        RECT 1.355 1.510 1.525 2.125 ;
        RECT 0.560 1.955 1.525 2.125 ;
        RECT 1.355 1.510 1.630 1.810 ;
        RECT 3.390 1.600 3.560 1.905 ;
        RECT 3.390 1.600 4.285 1.780 ;
        RECT 3.985 1.125 4.285 2.215 ;
        RECT 5.045 1.125 5.800 1.295 ;
        RECT 5.630 1.125 5.800 2.215 ;
        RECT 5.295 2.045 5.800 2.215 ;
        RECT 1.640 1.070 1.980 1.260 ;
        RECT 1.640 0.960 1.810 1.260 ;
        RECT 1.640 2.330 1.810 2.970 ;
        RECT 1.810 1.070 1.980 2.560 ;
        RECT 1.640 2.330 1.980 2.560 ;
        RECT 2.485 0.775 2.655 1.240 ;
        RECT 1.640 1.070 2.655 1.240 ;
        RECT 2.485 0.775 6.170 0.945 ;
        RECT 6.000 0.775 6.170 2.320 ;
        RECT 6.710 1.000 6.880 2.355 ;
        RECT 7.795 1.585 7.965 2.205 ;
        RECT 6.710 2.035 7.965 2.205 ;
        RECT 7.795 1.585 8.135 1.755 ;
        RECT 7.420 1.160 7.590 1.820 ;
        RECT 8.175 1.065 8.475 1.330 ;
        RECT 7.420 1.160 8.910 1.330 ;
        RECT 8.740 1.160 8.910 2.205 ;
        RECT 8.515 2.035 8.910 2.205 ;
        RECT 8.740 1.515 9.180 1.815 ;
        RECT 3.005 1.125 3.185 2.565 ;
        RECT 3.005 2.135 3.240 2.565 ;
        RECT 3.005 1.125 3.305 1.295 ;
        RECT 5.115 2.395 5.415 2.700 ;
        RECT 3.005 2.395 5.415 2.565 ;
        RECT 6.360 0.650 6.530 2.700 ;
        RECT 5.115 2.530 6.530 2.700 ;
        RECT 6.360 0.650 9.575 0.820 ;
        RECT 9.405 0.650 9.575 1.610 ;
        RECT 9.405 1.310 9.920 1.610 ;
        RECT 7.065 2.385 7.235 2.705 ;
        RECT 6.825 2.535 7.235 2.705 ;
        RECT 7.065 2.385 9.535 2.555 ;
        RECT 9.365 1.925 9.535 2.555 ;
        RECT 10.120 0.985 10.290 2.095 ;
        RECT 9.365 1.925 10.290 2.095 ;
        RECT 10.120 0.985 10.430 1.285 ;
        RECT 8.630 2.740 8.800 3.205 ;
        RECT 8.310 3.035 8.800 3.205 ;
        RECT 11.430 2.480 11.610 2.910 ;
        RECT 8.630 2.740 11.610 2.910 ;
        RECT 11.430 2.480 11.730 2.765 ;
        RECT 11.430 2.595 12.460 2.765 ;
        RECT 11.490 0.570 11.875 0.740 ;
        RECT 11.705 0.570 11.875 0.925 ;
        RECT 11.705 0.755 12.620 0.925 ;
        RECT 9.950 0.570 10.780 0.740 ;
        RECT 10.475 1.550 10.645 2.530 ;
        RECT 9.915 2.360 10.645 2.530 ;
        RECT 10.610 0.570 10.780 1.720 ;
        RECT 10.475 1.550 12.950 1.720 ;
        RECT 10.825 1.925 11.075 2.225 ;
        RECT 12.495 1.125 13.320 1.295 ;
        RECT 13.130 1.125 13.320 2.225 ;
        RECT 10.825 2.055 13.320 2.225 ;
  END 
END FFSDRHQHD1XHT

MACRO FFSDRHDMXHT
  CLASS  CORE ;
  FOREIGN FFSDRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.120 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 12.780 1.060 13.020 1.360 ;
        RECT 12.810 1.060 13.020 2.280 ;
        RECT 12.780 1.980 13.020 2.280 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.580 0.860 11.910 1.470 ;
        RECT 11.580 1.300 12.250 1.470 ;
        RECT 12.080 1.300 12.250 2.215 ;
        RECT 11.675 2.045 12.250 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 8.030 1.515 8.510 2.010 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.595 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.435 -0.300 2.735 0.595 ;
        RECT 3.245 -0.300 3.545 0.595 ;
        RECT 5.945 -0.300 6.245 1.145 ;
        RECT 7.055 -0.300 7.355 0.595 ;
        RECT 8.125 -0.300 8.295 0.810 ;
        RECT 10.065 -0.300 10.365 0.525 ;
        RECT 11.195 -0.300 11.495 0.530 ;
        RECT 12.225 -0.300 12.525 0.595 ;
        RECT 0.000 -0.300 13.120 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.740 1.525 3.230 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.545 2.740 3.185 3.990 ;
        RECT 6.005 3.195 6.305 3.990 ;
        RECT 8.165 3.195 8.465 3.990 ;
        RECT 10.165 2.810 10.465 3.990 ;
        RECT 12.225 2.925 12.525 3.990 ;
        RECT 0.000 3.390 13.120 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.525 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.055 ;
        RECT 1.530 0.885 1.700 2.280 ;
        RECT 1.945 0.775 2.115 1.055 ;
        RECT 1.530 0.885 2.115 1.055 ;
        RECT 1.945 0.775 4.510 0.945 ;
        RECT 4.340 0.775 4.510 2.280 ;
        RECT 4.340 1.960 4.520 2.280 ;
        RECT 4.340 1.970 4.530 2.280 ;
        RECT 4.340 1.980 4.540 2.280 ;
        RECT 5.070 0.910 5.210 2.280 ;
        RECT 6.235 1.675 6.535 1.865 ;
        RECT 5.440 1.695 6.535 1.865 ;
        RECT 5.240 1.505 5.250 1.865 ;
        RECT 5.250 1.515 5.260 1.865 ;
        RECT 5.260 1.525 5.270 1.865 ;
        RECT 5.270 1.535 5.280 1.865 ;
        RECT 5.280 1.545 5.290 1.865 ;
        RECT 5.290 1.555 5.300 1.865 ;
        RECT 5.300 1.565 5.310 1.865 ;
        RECT 5.310 1.575 5.320 1.865 ;
        RECT 5.320 1.585 5.330 1.865 ;
        RECT 5.330 1.595 5.340 1.865 ;
        RECT 5.340 1.605 5.350 1.865 ;
        RECT 5.350 1.615 5.360 1.865 ;
        RECT 5.360 1.625 5.370 1.865 ;
        RECT 5.370 1.635 5.380 1.865 ;
        RECT 5.380 1.645 5.390 1.865 ;
        RECT 5.390 1.655 5.400 1.865 ;
        RECT 5.400 1.665 5.410 1.865 ;
        RECT 5.410 1.675 5.420 1.865 ;
        RECT 5.420 1.685 5.430 1.865 ;
        RECT 5.430 1.695 5.440 1.865 ;
        RECT 5.210 1.475 5.220 2.279 ;
        RECT 5.220 1.485 5.230 2.279 ;
        RECT 5.230 1.495 5.240 2.279 ;
        RECT 5.040 0.910 5.050 1.574 ;
        RECT 5.050 0.910 5.060 1.584 ;
        RECT 5.060 0.910 5.070 1.594 ;
        RECT 5.685 1.325 5.985 1.515 ;
        RECT 6.650 0.775 6.885 1.495 ;
        RECT 5.685 1.325 6.885 1.495 ;
        RECT 6.715 0.775 6.885 2.215 ;
        RECT 6.715 2.045 7.255 2.215 ;
        RECT 7.540 0.480 7.710 0.945 ;
        RECT 6.650 0.775 7.710 0.945 ;
        RECT 2.725 1.125 3.585 1.295 ;
        RECT 2.785 2.190 3.585 2.360 ;
        RECT 3.415 1.125 3.585 2.985 ;
        RECT 3.415 1.525 3.710 1.825 ;
        RECT 8.460 2.745 8.630 2.985 ;
        RECT 3.415 2.815 8.630 2.985 ;
        RECT 8.460 2.745 9.205 2.915 ;
        RECT 3.765 1.125 4.085 1.295 ;
        RECT 3.860 1.980 4.085 2.280 ;
        RECT 3.915 1.125 4.085 2.635 ;
        RECT 4.700 1.745 4.890 1.825 ;
        RECT 4.710 1.745 4.890 1.835 ;
        RECT 4.690 0.535 4.860 1.815 ;
        RECT 4.690 1.725 4.870 1.815 ;
        RECT 4.690 1.735 4.880 1.815 ;
        RECT 4.720 1.745 4.890 2.635 ;
        RECT 4.690 0.535 5.485 0.705 ;
        RECT 8.105 2.395 8.275 2.635 ;
        RECT 3.915 2.465 8.275 2.635 ;
        RECT 8.825 1.330 8.995 2.565 ;
        RECT 8.825 1.330 9.125 1.500 ;
        RECT 8.105 2.395 9.720 2.565 ;
        RECT 9.550 2.395 9.720 2.695 ;
        RECT 7.065 1.615 7.810 1.785 ;
        RECT 7.640 1.125 7.810 2.280 ;
        RECT 8.475 0.605 8.645 1.295 ;
        RECT 7.615 1.125 8.645 1.295 ;
        RECT 9.690 0.605 9.860 0.945 ;
        RECT 8.475 0.605 9.860 0.775 ;
        RECT 9.690 0.775 11.335 0.945 ;
        RECT 11.165 0.775 11.335 1.515 ;
        RECT 10.615 1.125 10.985 1.495 ;
        RECT 9.855 1.325 10.985 1.495 ;
        RECT 10.815 1.125 10.985 1.865 ;
        RECT 11.150 1.695 11.320 2.280 ;
        RECT 11.600 1.675 11.900 1.865 ;
        RECT 10.815 1.695 11.900 1.865 ;
        RECT 9.115 0.955 9.475 1.125 ;
        RECT 9.305 0.955 9.475 2.215 ;
        RECT 9.220 2.045 9.520 2.215 ;
        RECT 9.305 1.675 10.635 1.845 ;
        RECT 10.465 1.675 10.635 2.630 ;
        RECT 12.430 1.610 12.600 2.630 ;
        RECT 10.465 2.460 12.600 2.630 ;
  END 
END FFSDRHDMXHT

MACRO FFSDRHDLXHT
  CLASS  CORE ;
  FOREIGN FFSDRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.120 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 12.780 1.060 13.020 2.455 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.580 0.860 11.910 1.470 ;
        RECT 11.580 1.300 12.250 1.470 ;
        RECT 12.080 1.300 12.250 2.215 ;
        RECT 11.675 2.045 12.250 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 8.030 1.535 8.510 2.010 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.595 2.980 ;
        RECT 0.100 2.810 1.350 2.980 ;
        RECT 1.180 2.810 1.350 3.135 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.435 -0.300 2.735 0.595 ;
        RECT 3.395 -0.300 3.695 0.595 ;
        RECT 6.035 -0.300 6.335 1.145 ;
        RECT 7.055 -0.300 7.355 0.595 ;
        RECT 8.125 -0.300 8.295 0.810 ;
        RECT 10.065 -0.300 10.365 0.525 ;
        RECT 11.195 -0.300 11.495 0.530 ;
        RECT 12.225 -0.300 12.525 0.745 ;
        RECT 0.000 -0.300 13.120 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.800 1.525 3.290 1.950 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.935 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.645 2.650 3.285 3.990 ;
        RECT 6.035 3.165 6.335 3.990 ;
        RECT 8.165 3.165 8.465 3.990 ;
        RECT 10.165 2.810 10.465 3.990 ;
        RECT 12.225 2.810 12.525 3.990 ;
        RECT 0.000 3.390 13.120 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.535 1.350 2.630 ;
        RECT 1.180 0.535 1.525 0.705 ;
        RECT 1.180 2.460 1.880 2.630 ;
        RECT 1.710 2.460 1.880 2.825 ;
        RECT 1.530 0.885 1.700 2.280 ;
        RECT 1.530 0.885 1.720 1.185 ;
        RECT 1.980 0.775 2.150 1.055 ;
        RECT 1.530 0.885 2.150 1.055 ;
        RECT 1.980 0.775 4.600 0.945 ;
        RECT 4.430 0.775 4.600 2.280 ;
        RECT 5.130 0.900 5.300 2.280 ;
        RECT 6.235 1.675 6.535 1.865 ;
        RECT 5.130 1.695 6.535 1.865 ;
        RECT 5.755 1.325 6.055 1.515 ;
        RECT 6.650 0.775 6.885 1.495 ;
        RECT 5.755 1.325 6.885 1.495 ;
        RECT 6.715 0.775 6.885 2.215 ;
        RECT 6.715 2.045 7.255 2.215 ;
        RECT 7.540 0.480 7.710 0.945 ;
        RECT 6.650 0.775 7.710 0.945 ;
        RECT 2.815 1.125 3.645 1.295 ;
        RECT 2.815 2.130 3.645 2.300 ;
        RECT 3.475 1.125 3.645 2.985 ;
        RECT 3.475 1.525 3.800 1.825 ;
        RECT 8.460 2.745 8.630 2.985 ;
        RECT 3.475 2.815 8.630 2.985 ;
        RECT 8.460 2.745 9.045 2.915 ;
        RECT 3.855 1.125 4.175 1.295 ;
        RECT 4.005 1.125 4.175 2.635 ;
        RECT 4.780 0.535 4.950 2.635 ;
        RECT 4.780 0.535 5.575 0.705 ;
        RECT 8.105 2.395 8.275 2.635 ;
        RECT 3.885 2.465 8.275 2.635 ;
        RECT 8.825 1.330 8.995 2.565 ;
        RECT 8.825 1.330 9.125 1.500 ;
        RECT 8.105 2.395 9.720 2.565 ;
        RECT 9.550 2.395 9.720 2.695 ;
        RECT 7.065 1.595 7.810 1.765 ;
        RECT 7.640 1.125 7.810 2.280 ;
        RECT 8.475 0.605 8.645 1.295 ;
        RECT 7.615 1.125 8.645 1.295 ;
        RECT 9.690 0.605 9.860 0.945 ;
        RECT 8.475 0.605 9.860 0.775 ;
        RECT 9.690 0.775 11.335 0.945 ;
        RECT 11.165 0.775 11.335 1.515 ;
        RECT 9.855 1.325 10.985 1.495 ;
        RECT 10.615 1.125 10.915 1.495 ;
        RECT 10.815 1.325 10.985 1.865 ;
        RECT 11.150 1.695 11.320 2.280 ;
        RECT 11.600 1.675 11.900 1.865 ;
        RECT 10.815 1.695 11.900 1.865 ;
        RECT 9.115 0.955 9.475 1.125 ;
        RECT 9.305 0.955 9.475 2.215 ;
        RECT 9.220 2.045 9.520 2.215 ;
        RECT 9.305 1.675 10.635 1.845 ;
        RECT 10.465 1.675 10.635 2.630 ;
        RECT 12.430 1.610 12.600 2.630 ;
        RECT 10.465 2.460 12.600 2.630 ;
  END 
END FFSDRHDLXHT

MACRO FFSDRHD2XHT
  CLASS  CORE ;
  FOREIGN FFSDRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.940 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.080 0.720 13.250 2.960 ;
        RECT 13.080 1.645 13.430 2.015 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.990 0.720 12.210 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.940 1.530 8.530 1.830 ;
        RECT 8.140 1.530 8.530 2.130 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.595 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.265 -0.300 2.565 0.595 ;
        RECT 3.325 -0.300 3.625 0.595 ;
        RECT 5.895 -0.300 6.195 1.055 ;
        RECT 6.965 -0.300 7.265 0.595 ;
        RECT 8.070 -0.300 8.370 0.715 ;
        RECT 9.970 -0.300 10.270 0.595 ;
        RECT 11.455 -0.300 11.755 1.055 ;
        RECT 12.495 -0.300 12.795 1.055 ;
        RECT 13.535 -0.300 13.835 1.055 ;
        RECT 0.000 -0.300 13.940 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.730 1.525 3.220 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.925 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.565 2.830 3.205 3.990 ;
        RECT 5.910 3.140 6.210 3.990 ;
        RECT 8.070 3.095 8.370 3.990 ;
        RECT 10.070 2.810 10.370 3.990 ;
        RECT 11.455 2.975 11.755 3.990 ;
        RECT 12.495 2.975 12.795 3.990 ;
        RECT 13.535 2.295 13.835 3.990 ;
        RECT 0.000 3.390 13.940 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.555 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.150 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.965 0.775 2.135 1.035 ;
        RECT 1.530 0.865 2.135 1.035 ;
        RECT 1.965 0.775 4.500 0.945 ;
        RECT 4.330 0.775 4.500 2.280 ;
        RECT 5.030 0.910 5.200 2.280 ;
        RECT 6.105 1.675 6.405 1.865 ;
        RECT 5.030 1.695 6.405 1.865 ;
        RECT 5.625 1.325 5.925 1.515 ;
        RECT 5.625 1.325 6.755 1.495 ;
        RECT 6.480 0.775 6.650 1.495 ;
        RECT 6.585 1.325 6.755 2.215 ;
        RECT 6.585 2.045 7.235 2.215 ;
        RECT 7.445 0.480 7.615 0.945 ;
        RECT 6.480 0.775 7.615 0.945 ;
        RECT 2.775 1.125 3.575 1.295 ;
        RECT 2.775 2.190 3.575 2.360 ;
        RECT 3.405 1.125 3.575 3.035 ;
        RECT 3.405 1.525 3.700 1.825 ;
        RECT 5.575 2.815 5.645 3.035 ;
        RECT 5.565 2.825 8.940 2.915 ;
        RECT 5.585 2.805 5.645 3.035 ;
        RECT 5.555 2.835 8.940 2.915 ;
        RECT 5.595 2.795 5.645 3.035 ;
        RECT 5.545 2.845 8.940 2.915 ;
        RECT 3.405 2.865 5.645 3.035 ;
        RECT 3.405 2.865 5.655 3.024 ;
        RECT 3.405 2.865 5.665 3.014 ;
        RECT 3.405 2.865 5.675 3.004 ;
        RECT 3.405 2.865 5.685 2.994 ;
        RECT 3.405 2.865 5.695 2.984 ;
        RECT 3.405 2.865 5.705 2.974 ;
        RECT 3.405 2.865 5.715 2.964 ;
        RECT 5.600 2.790 7.920 2.960 ;
        RECT 5.535 2.855 8.940 2.915 ;
        RECT 7.750 2.745 7.920 2.960 ;
        RECT 7.750 2.745 8.940 2.915 ;
        RECT 8.770 2.745 8.940 3.210 ;
        RECT 8.770 3.040 9.600 3.210 ;
        RECT 3.755 1.125 4.075 1.295 ;
        RECT 3.880 1.125 4.075 2.635 ;
        RECT 3.820 1.980 4.075 2.635 ;
        RECT 4.680 0.535 4.850 2.685 ;
        RECT 4.595 2.465 4.895 2.685 ;
        RECT 5.335 2.445 9.625 2.565 ;
        RECT 3.820 2.465 5.435 2.635 ;
        RECT 4.680 0.535 5.445 0.705 ;
        RECT 3.820 2.465 5.445 2.624 ;
        RECT 3.820 2.465 5.455 2.614 ;
        RECT 5.340 2.440 7.565 2.610 ;
        RECT 5.325 2.455 9.625 2.565 ;
        RECT 7.395 2.395 7.565 2.610 ;
        RECT 8.730 1.355 8.900 2.565 ;
        RECT 8.730 1.355 9.030 1.525 ;
        RECT 7.395 2.395 9.625 2.565 ;
        RECT 9.455 2.395 9.625 2.795 ;
        RECT 6.935 1.590 7.760 1.760 ;
        RECT 7.590 1.125 7.760 2.215 ;
        RECT 7.520 2.045 7.820 2.215 ;
        RECT 8.020 0.960 8.190 1.295 ;
        RECT 7.520 1.125 8.190 1.295 ;
        RECT 8.020 0.960 8.775 1.130 ;
        RECT 8.605 0.635 8.775 1.130 ;
        RECT 9.605 0.635 9.775 0.945 ;
        RECT 8.605 0.635 9.775 0.805 ;
        RECT 9.605 0.775 11.240 0.945 ;
        RECT 11.070 0.775 11.240 1.490 ;
        RECT 10.520 1.125 10.890 1.495 ;
        RECT 9.710 1.325 10.890 1.495 ;
        RECT 10.720 1.125 10.890 1.845 ;
        RECT 11.055 1.675 11.225 2.280 ;
        RECT 10.720 1.675 11.810 1.845 ;
        RECT 9.020 0.985 9.425 1.155 ;
        RECT 9.255 0.985 9.425 2.215 ;
        RECT 9.125 2.045 9.425 2.215 ;
        RECT 9.255 1.675 10.540 1.845 ;
        RECT 10.370 1.675 10.540 2.630 ;
        RECT 12.730 1.610 12.900 2.630 ;
        RECT 10.370 2.460 12.900 2.630 ;
  END 
END FFSDRHD2XHT

MACRO FFSDRHD1XHT
  CLASS  CORE ;
  FOREIGN FFSDRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.120 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 12.780 0.720 13.020 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.580 0.720 11.910 1.470 ;
        RECT 11.580 1.300 12.250 1.470 ;
        RECT 12.080 1.300 12.250 2.215 ;
        RECT 11.675 2.045 12.250 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 8.030 1.510 8.510 2.010 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.595 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.385 -0.300 2.685 0.595 ;
        RECT 3.335 -0.300 3.635 0.595 ;
        RECT 5.945 -0.300 6.245 1.145 ;
        RECT 7.055 -0.300 7.355 0.545 ;
        RECT 8.125 -0.300 8.295 0.810 ;
        RECT 10.065 -0.300 10.365 0.525 ;
        RECT 11.165 -0.300 11.465 0.480 ;
        RECT 12.195 -0.300 12.495 1.055 ;
        RECT 0.000 -0.300 13.120 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.740 1.525 3.230 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.590 2.740 3.230 3.990 ;
        RECT 5.995 3.195 6.295 3.990 ;
        RECT 8.165 3.195 8.465 3.990 ;
        RECT 10.230 2.810 10.400 3.990 ;
        RECT 12.195 2.975 12.495 3.990 ;
        RECT 0.000 3.390 13.120 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.575 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.150 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.995 0.775 2.165 1.035 ;
        RECT 1.530 0.865 2.165 1.035 ;
        RECT 1.995 0.775 4.510 0.945 ;
        RECT 4.340 0.775 4.510 2.280 ;
        RECT 5.040 0.900 5.210 2.280 ;
        RECT 6.235 1.675 6.535 1.865 ;
        RECT 5.040 1.695 6.535 1.865 ;
        RECT 5.685 1.325 5.985 1.515 ;
        RECT 6.650 0.775 6.885 1.495 ;
        RECT 5.685 1.325 6.885 1.495 ;
        RECT 6.715 0.775 6.885 2.215 ;
        RECT 6.715 2.045 7.255 2.215 ;
        RECT 7.540 0.480 7.710 0.945 ;
        RECT 6.650 0.775 7.710 0.945 ;
        RECT 2.785 1.125 3.585 1.295 ;
        RECT 2.785 2.190 3.585 2.360 ;
        RECT 3.415 1.125 3.585 2.985 ;
        RECT 3.415 1.525 3.710 1.825 ;
        RECT 8.460 2.745 8.630 2.985 ;
        RECT 3.415 2.815 8.630 2.985 ;
        RECT 8.460 2.745 9.205 2.915 ;
        RECT 3.830 1.980 4.085 2.280 ;
        RECT 3.765 1.125 4.085 1.295 ;
        RECT 3.890 1.125 4.085 2.635 ;
        RECT 3.850 1.980 4.085 2.635 ;
        RECT 4.690 0.535 4.860 2.635 ;
        RECT 4.690 0.535 5.485 0.705 ;
        RECT 8.105 2.395 8.275 2.635 ;
        RECT 3.850 2.465 8.275 2.635 ;
        RECT 8.825 1.330 8.995 2.565 ;
        RECT 8.825 1.330 9.125 1.500 ;
        RECT 8.105 2.395 9.720 2.565 ;
        RECT 9.550 2.395 9.720 2.795 ;
        RECT 7.065 1.585 7.810 1.755 ;
        RECT 7.640 1.125 7.810 2.280 ;
        RECT 8.475 0.605 8.645 1.295 ;
        RECT 7.615 1.125 8.645 1.295 ;
        RECT 9.690 0.605 9.860 0.945 ;
        RECT 8.475 0.605 9.860 0.775 ;
        RECT 9.690 0.775 11.335 0.945 ;
        RECT 11.165 0.775 11.335 1.515 ;
        RECT 10.615 1.125 10.985 1.495 ;
        RECT 9.805 1.325 10.985 1.495 ;
        RECT 10.815 1.125 10.985 1.865 ;
        RECT 11.150 1.695 11.320 2.280 ;
        RECT 11.600 1.675 11.900 1.865 ;
        RECT 10.815 1.695 11.900 1.865 ;
        RECT 9.115 0.955 9.475 1.125 ;
        RECT 9.305 0.955 9.475 2.215 ;
        RECT 9.220 2.045 9.520 2.215 ;
        RECT 9.305 1.675 10.635 1.845 ;
        RECT 10.465 1.675 10.635 2.630 ;
        RECT 12.430 1.610 12.600 2.630 ;
        RECT 10.465 2.460 12.600 2.630 ;
  END 
END FFSDRHD1XHT

MACRO FFSDQSRHDMXHT
  CLASS  CORE ;
  FOREIGN FFSDQSRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.530 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.190 1.045 13.430 2.280 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.835 1.290 1.605 1.540 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.760 1.540 6.385 1.955 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.520 1.735 0.690 2.100 ;
        RECT 0.815 1.930 1.230 2.360 ;
        RECT 1.400 1.735 1.570 2.100 ;
        RECT 0.520 1.930 1.570 2.100 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.995 ;
        RECT 2.525 -0.300 3.505 0.785 ;
        RECT 5.970 -0.300 6.270 1.130 ;
        RECT 8.765 -0.300 8.935 0.890 ;
        RECT 10.645 -0.300 10.945 0.795 ;
        RECT 12.575 -0.300 12.875 0.715 ;
        RECT 0.000 -0.300 13.530 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.965 1.550 3.305 2.015 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.290 1.610 2.775 2.015 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 12.175 1.540 12.640 2.015 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.905 0.895 3.990 ;
        RECT 2.540 2.895 3.520 3.990 ;
        RECT 6.145 2.995 7.125 3.990 ;
        RECT 8.675 2.995 8.975 3.990 ;
        RECT 10.700 2.315 11.000 3.990 ;
        RECT 12.545 2.975 12.845 3.990 ;
        RECT 0.000 3.390 13.530 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.170 0.340 2.470 ;
        RECT 0.105 0.825 0.275 2.470 ;
        RECT 0.170 2.170 0.340 2.725 ;
        RECT 0.105 0.825 0.405 0.995 ;
        RECT 0.170 2.555 1.305 2.725 ;
        RECT 1.135 2.555 1.305 3.125 ;
        RECT 1.135 2.955 1.995 3.125 ;
        RECT 2.740 1.125 3.690 1.295 ;
        RECT 3.530 1.525 3.750 1.619 ;
        RECT 3.540 1.525 3.750 1.629 ;
        RECT 3.550 1.525 3.750 1.639 ;
        RECT 3.560 1.525 3.750 1.649 ;
        RECT 3.570 1.525 3.750 1.659 ;
        RECT 3.520 1.125 3.690 1.609 ;
        RECT 3.520 1.475 3.700 1.609 ;
        RECT 3.520 1.485 3.710 1.609 ;
        RECT 3.520 1.495 3.720 1.609 ;
        RECT 3.520 1.505 3.730 1.609 ;
        RECT 3.520 1.515 3.740 1.609 ;
        RECT 3.580 1.525 3.750 2.365 ;
        RECT 2.825 2.195 3.750 2.365 ;
        RECT 1.575 0.695 1.985 0.865 ;
        RECT 1.815 0.695 1.985 2.715 ;
        RECT 1.580 2.370 1.985 2.715 ;
        RECT 1.580 2.545 3.655 2.715 ;
        RECT 4.445 0.895 4.555 2.830 ;
        RECT 3.845 2.660 4.555 2.830 ;
        RECT 4.555 1.945 4.565 2.829 ;
        RECT 4.565 1.955 4.575 2.829 ;
        RECT 4.575 1.965 4.585 2.829 ;
        RECT 4.585 1.975 4.595 2.829 ;
        RECT 4.595 1.985 4.605 2.829 ;
        RECT 4.605 1.995 4.615 2.829 ;
        RECT 4.385 0.895 4.395 2.105 ;
        RECT 4.395 0.895 4.405 2.115 ;
        RECT 4.405 0.895 4.415 2.125 ;
        RECT 4.415 0.895 4.425 2.135 ;
        RECT 4.425 0.895 4.435 2.145 ;
        RECT 4.435 0.895 4.445 2.155 ;
        RECT 3.770 2.595 3.780 2.829 ;
        RECT 3.780 2.605 3.790 2.829 ;
        RECT 3.790 2.615 3.800 2.829 ;
        RECT 3.800 2.625 3.810 2.829 ;
        RECT 3.810 2.635 3.820 2.829 ;
        RECT 3.820 2.645 3.830 2.829 ;
        RECT 3.830 2.655 3.840 2.829 ;
        RECT 3.840 2.660 3.846 2.830 ;
        RECT 3.730 2.555 3.740 2.789 ;
        RECT 3.740 2.565 3.750 2.799 ;
        RECT 3.750 2.575 3.760 2.809 ;
        RECT 3.760 2.585 3.770 2.819 ;
        RECT 3.655 2.545 3.665 2.715 ;
        RECT 3.665 2.545 3.675 2.725 ;
        RECT 3.675 2.545 3.685 2.735 ;
        RECT 3.685 2.545 3.695 2.745 ;
        RECT 3.695 2.545 3.705 2.755 ;
        RECT 3.705 2.545 3.715 2.765 ;
        RECT 3.715 2.545 3.725 2.775 ;
        RECT 3.725 2.545 3.731 2.785 ;
        RECT 6.585 0.960 6.755 2.115 ;
        RECT 6.490 0.960 6.790 1.130 ;
        RECT 6.585 1.500 7.360 1.670 ;
        RECT 5.095 1.335 5.315 1.425 ;
        RECT 5.105 1.335 5.315 1.435 ;
        RECT 5.115 1.335 5.315 1.445 ;
        RECT 5.125 1.335 5.315 1.455 ;
        RECT 5.135 1.335 5.315 1.465 ;
        RECT 5.085 0.895 5.255 1.415 ;
        RECT 5.085 1.285 5.265 1.415 ;
        RECT 5.085 1.295 5.275 1.415 ;
        RECT 5.085 1.305 5.285 1.415 ;
        RECT 5.085 1.315 5.295 1.415 ;
        RECT 5.085 1.325 5.305 1.415 ;
        RECT 5.145 1.335 5.315 2.465 ;
        RECT 7.540 1.680 7.710 2.465 ;
        RECT 5.145 2.295 7.710 2.465 ;
        RECT 7.775 1.550 7.945 1.850 ;
        RECT 7.540 1.680 7.945 1.850 ;
        RECT 7.000 0.960 7.300 1.230 ;
        RECT 7.000 1.060 8.235 1.230 ;
        RECT 8.065 1.060 8.235 1.360 ;
        RECT 6.630 0.480 6.930 0.730 ;
        RECT 7.890 2.045 8.015 2.215 ;
        RECT 8.125 1.580 8.190 2.215 ;
        RECT 6.630 0.560 8.585 0.730 ;
        RECT 8.415 0.560 8.585 1.750 ;
        RECT 8.295 1.580 9.180 1.750 ;
        RECT 8.190 1.580 8.200 2.104 ;
        RECT 8.200 1.580 8.210 2.094 ;
        RECT 8.210 1.580 8.220 2.084 ;
        RECT 8.220 1.580 8.230 2.074 ;
        RECT 8.230 1.580 8.240 2.064 ;
        RECT 8.240 1.580 8.250 2.054 ;
        RECT 8.250 1.580 8.260 2.044 ;
        RECT 8.260 1.580 8.270 2.034 ;
        RECT 8.270 1.580 8.280 2.024 ;
        RECT 8.280 1.580 8.290 2.014 ;
        RECT 8.290 1.580 8.296 2.010 ;
        RECT 8.015 2.045 8.025 2.215 ;
        RECT 8.025 2.035 8.035 2.215 ;
        RECT 8.035 2.025 8.045 2.215 ;
        RECT 8.045 2.015 8.055 2.215 ;
        RECT 8.055 2.005 8.065 2.215 ;
        RECT 8.065 1.995 8.075 2.215 ;
        RECT 8.075 1.985 8.085 2.215 ;
        RECT 8.085 1.975 8.095 2.215 ;
        RECT 8.095 1.965 8.105 2.215 ;
        RECT 8.105 1.955 8.115 2.215 ;
        RECT 8.115 1.945 8.125 2.215 ;
        RECT 3.930 0.520 4.100 2.430 ;
        RECT 3.930 0.520 4.735 0.690 ;
        RECT 4.795 0.520 4.905 2.835 ;
        RECT 4.795 0.520 5.530 0.690 ;
        RECT 4.965 2.645 8.020 2.815 ;
        RECT 8.445 2.295 9.205 2.465 ;
        RECT 9.380 2.395 10.105 2.565 ;
        RECT 9.935 2.395 10.105 2.695 ;
        RECT 9.305 2.330 9.315 2.564 ;
        RECT 9.315 2.340 9.325 2.564 ;
        RECT 9.325 2.350 9.335 2.564 ;
        RECT 9.335 2.360 9.345 2.564 ;
        RECT 9.345 2.370 9.355 2.564 ;
        RECT 9.355 2.380 9.365 2.564 ;
        RECT 9.365 2.390 9.375 2.564 ;
        RECT 9.375 2.395 9.381 2.565 ;
        RECT 9.280 2.305 9.290 2.539 ;
        RECT 9.290 2.315 9.300 2.549 ;
        RECT 9.300 2.320 9.306 2.560 ;
        RECT 9.205 2.295 9.215 2.465 ;
        RECT 9.215 2.295 9.225 2.475 ;
        RECT 9.225 2.295 9.235 2.485 ;
        RECT 9.235 2.295 9.245 2.495 ;
        RECT 9.245 2.295 9.255 2.505 ;
        RECT 9.255 2.295 9.265 2.515 ;
        RECT 9.265 2.295 9.275 2.525 ;
        RECT 9.275 2.295 9.281 2.535 ;
        RECT 8.370 2.295 8.380 2.529 ;
        RECT 8.380 2.295 8.390 2.519 ;
        RECT 8.390 2.295 8.400 2.509 ;
        RECT 8.400 2.295 8.410 2.499 ;
        RECT 8.410 2.295 8.420 2.489 ;
        RECT 8.420 2.295 8.430 2.479 ;
        RECT 8.430 2.295 8.440 2.469 ;
        RECT 8.440 2.295 8.446 2.465 ;
        RECT 8.095 2.570 8.105 2.804 ;
        RECT 8.105 2.560 8.115 2.794 ;
        RECT 8.115 2.550 8.125 2.784 ;
        RECT 8.125 2.540 8.135 2.774 ;
        RECT 8.135 2.530 8.145 2.764 ;
        RECT 8.145 2.520 8.155 2.754 ;
        RECT 8.155 2.510 8.165 2.744 ;
        RECT 8.165 2.500 8.175 2.734 ;
        RECT 8.175 2.490 8.185 2.724 ;
        RECT 8.185 2.480 8.195 2.714 ;
        RECT 8.195 2.470 8.205 2.704 ;
        RECT 8.205 2.460 8.215 2.694 ;
        RECT 8.215 2.450 8.225 2.684 ;
        RECT 8.225 2.440 8.235 2.674 ;
        RECT 8.235 2.430 8.245 2.664 ;
        RECT 8.245 2.420 8.255 2.654 ;
        RECT 8.255 2.410 8.265 2.644 ;
        RECT 8.265 2.400 8.275 2.634 ;
        RECT 8.275 2.390 8.285 2.624 ;
        RECT 8.285 2.380 8.295 2.614 ;
        RECT 8.295 2.370 8.305 2.604 ;
        RECT 8.305 2.360 8.315 2.594 ;
        RECT 8.315 2.350 8.325 2.584 ;
        RECT 8.325 2.340 8.335 2.574 ;
        RECT 8.335 2.330 8.345 2.564 ;
        RECT 8.345 2.320 8.355 2.554 ;
        RECT 8.355 2.310 8.365 2.544 ;
        RECT 8.365 2.300 8.371 2.540 ;
        RECT 8.020 2.645 8.030 2.815 ;
        RECT 8.030 2.635 8.040 2.815 ;
        RECT 8.040 2.625 8.050 2.815 ;
        RECT 8.050 2.615 8.060 2.815 ;
        RECT 8.060 2.605 8.070 2.815 ;
        RECT 8.070 2.595 8.080 2.815 ;
        RECT 8.080 2.585 8.090 2.815 ;
        RECT 8.090 2.575 8.096 2.815 ;
        RECT 4.905 1.560 4.915 2.834 ;
        RECT 4.915 1.570 4.925 2.834 ;
        RECT 4.925 1.580 4.935 2.834 ;
        RECT 4.935 1.590 4.945 2.834 ;
        RECT 4.945 1.600 4.955 2.834 ;
        RECT 4.955 1.610 4.965 2.834 ;
        RECT 4.735 0.520 4.745 1.660 ;
        RECT 4.745 0.520 4.755 1.670 ;
        RECT 4.755 0.520 4.765 1.680 ;
        RECT 4.765 0.520 4.775 1.690 ;
        RECT 4.775 0.520 4.785 1.700 ;
        RECT 4.785 0.520 4.795 1.710 ;
        RECT 3.875 0.520 3.885 1.360 ;
        RECT 3.885 0.520 3.895 1.370 ;
        RECT 3.895 0.520 3.905 1.380 ;
        RECT 3.905 0.520 3.915 1.390 ;
        RECT 3.915 0.520 3.925 1.400 ;
        RECT 3.925 0.520 3.931 1.410 ;
        RECT 7.340 2.995 7.640 3.210 ;
        RECT 7.340 2.995 8.325 3.165 ;
        RECT 8.595 2.645 9.050 2.815 ;
        RECT 9.495 2.745 9.665 3.045 ;
        RECT 9.225 2.745 9.665 2.915 ;
        RECT 9.955 1.270 10.255 1.440 ;
        RECT 10.085 1.270 10.255 1.825 ;
        RECT 10.085 1.655 10.455 1.825 ;
        RECT 10.285 1.655 10.455 3.045 ;
        RECT 9.495 2.875 10.455 3.045 ;
        RECT 9.150 2.680 9.160 2.914 ;
        RECT 9.160 2.690 9.170 2.914 ;
        RECT 9.170 2.700 9.180 2.914 ;
        RECT 9.180 2.710 9.190 2.914 ;
        RECT 9.190 2.720 9.200 2.914 ;
        RECT 9.200 2.730 9.210 2.914 ;
        RECT 9.210 2.740 9.220 2.914 ;
        RECT 9.220 2.745 9.226 2.915 ;
        RECT 9.125 2.655 9.135 2.889 ;
        RECT 9.135 2.665 9.145 2.899 ;
        RECT 9.145 2.670 9.151 2.910 ;
        RECT 9.050 2.645 9.060 2.815 ;
        RECT 9.060 2.645 9.070 2.825 ;
        RECT 9.070 2.645 9.080 2.835 ;
        RECT 9.080 2.645 9.090 2.845 ;
        RECT 9.090 2.645 9.100 2.855 ;
        RECT 9.100 2.645 9.110 2.865 ;
        RECT 9.110 2.645 9.120 2.875 ;
        RECT 9.120 2.645 9.126 2.885 ;
        RECT 8.520 2.645 8.530 2.879 ;
        RECT 8.530 2.645 8.540 2.869 ;
        RECT 8.540 2.645 8.550 2.859 ;
        RECT 8.550 2.645 8.560 2.849 ;
        RECT 8.560 2.645 8.570 2.839 ;
        RECT 8.570 2.645 8.580 2.829 ;
        RECT 8.580 2.645 8.590 2.819 ;
        RECT 8.590 2.645 8.596 2.815 ;
        RECT 8.495 2.670 8.505 2.904 ;
        RECT 8.505 2.660 8.515 2.894 ;
        RECT 8.515 2.650 8.521 2.890 ;
        RECT 8.325 2.840 8.335 3.164 ;
        RECT 8.335 2.830 8.345 3.164 ;
        RECT 8.345 2.820 8.355 3.164 ;
        RECT 8.355 2.810 8.365 3.164 ;
        RECT 8.365 2.800 8.375 3.164 ;
        RECT 8.375 2.790 8.385 3.164 ;
        RECT 8.385 2.780 8.395 3.164 ;
        RECT 8.395 2.770 8.405 3.164 ;
        RECT 8.405 2.760 8.415 3.164 ;
        RECT 8.415 2.750 8.425 3.164 ;
        RECT 8.425 2.740 8.435 3.164 ;
        RECT 8.435 2.730 8.445 3.164 ;
        RECT 8.445 2.720 8.455 3.164 ;
        RECT 8.455 2.710 8.465 3.164 ;
        RECT 8.465 2.700 8.475 3.164 ;
        RECT 8.475 2.690 8.485 3.164 ;
        RECT 8.485 2.680 8.495 3.164 ;
        RECT 10.985 1.460 11.155 1.760 ;
        RECT 11.595 1.110 11.895 1.630 ;
        RECT 10.985 1.460 11.895 1.630 ;
        RECT 11.725 1.110 11.895 2.365 ;
        RECT 11.725 2.195 12.295 2.365 ;
        RECT 11.205 0.760 11.375 1.280 ;
        RECT 11.075 1.110 11.375 1.280 ;
        RECT 11.205 0.760 12.285 0.930 ;
        RECT 12.115 0.760 12.285 1.280 ;
        RECT 12.115 1.110 12.415 1.280 ;
        RECT 9.545 0.900 9.715 2.215 ;
        RECT 9.545 2.045 9.850 2.215 ;
        RECT 9.545 0.900 10.330 1.070 ;
        RECT 10.565 1.060 10.805 1.230 ;
        RECT 10.635 1.060 10.805 2.110 ;
        RECT 10.635 1.940 11.390 2.110 ;
        RECT 11.220 1.940 11.390 2.795 ;
        RECT 11.815 2.625 12.115 2.855 ;
        RECT 12.840 1.610 13.010 2.795 ;
        RECT 11.220 2.625 13.010 2.795 ;
        RECT 10.490 0.995 10.500 1.229 ;
        RECT 10.500 1.005 10.510 1.229 ;
        RECT 10.510 1.015 10.520 1.229 ;
        RECT 10.520 1.025 10.530 1.229 ;
        RECT 10.530 1.035 10.540 1.229 ;
        RECT 10.540 1.045 10.550 1.229 ;
        RECT 10.550 1.055 10.560 1.229 ;
        RECT 10.560 1.060 10.566 1.230 ;
        RECT 10.405 0.910 10.415 1.144 ;
        RECT 10.415 0.920 10.425 1.154 ;
        RECT 10.425 0.930 10.435 1.164 ;
        RECT 10.435 0.940 10.445 1.174 ;
        RECT 10.445 0.950 10.455 1.184 ;
        RECT 10.455 0.960 10.465 1.194 ;
        RECT 10.465 0.970 10.475 1.204 ;
        RECT 10.475 0.980 10.485 1.214 ;
        RECT 10.485 0.985 10.491 1.225 ;
        RECT 10.330 0.900 10.340 1.070 ;
        RECT 10.340 0.900 10.350 1.080 ;
        RECT 10.350 0.900 10.360 1.090 ;
        RECT 10.360 0.900 10.370 1.100 ;
        RECT 10.370 0.900 10.380 1.110 ;
        RECT 10.380 0.900 10.390 1.120 ;
        RECT 10.390 0.900 10.400 1.130 ;
        RECT 10.400 0.900 10.406 1.140 ;
  END 
END FFSDQSRHDMXHT

MACRO FFSDQSRHD2XHT
  CLASS  CORE ;
  FOREIGN FFSDQSRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.350 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.490 0.720 13.660 2.960 ;
        RECT 13.490 1.615 13.840 2.055 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.870 1.240 1.605 1.540 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.675 1.460 6.120 1.955 ;
        RECT 5.675 1.460 6.315 1.695 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.520 1.735 0.690 2.100 ;
        RECT 0.815 1.930 1.290 2.365 ;
        RECT 1.400 1.735 1.570 2.100 ;
        RECT 0.520 1.930 1.570 2.100 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.060 ;
        RECT 2.465 -0.300 2.765 0.515 ;
        RECT 3.340 -0.300 3.640 0.715 ;
        RECT 5.870 -0.300 6.170 1.195 ;
        RECT 8.795 -0.300 8.965 1.360 ;
        RECT 10.740 -0.300 11.040 0.815 ;
        RECT 12.905 -0.300 13.205 1.055 ;
        RECT 13.945 -0.300 14.245 1.055 ;
        RECT 0.000 -0.300 14.350 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.970 1.670 3.360 2.015 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.290 1.610 2.770 2.015 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 12.330 1.330 12.770 1.755 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.915 0.895 3.990 ;
        RECT 2.515 2.895 3.495 3.990 ;
        RECT 5.980 2.995 6.960 3.990 ;
        RECT 8.650 2.995 8.950 3.990 ;
        RECT 10.690 2.750 11.330 3.990 ;
        RECT 12.905 2.295 13.205 3.990 ;
        RECT 13.945 2.295 14.245 3.990 ;
        RECT 0.000 3.390 14.350 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.890 0.275 2.735 ;
        RECT 0.105 2.225 0.340 2.735 ;
        RECT 0.105 0.890 0.405 1.060 ;
        RECT 0.105 2.565 1.340 2.735 ;
        RECT 1.170 2.565 1.340 3.210 ;
        RECT 1.170 3.040 1.995 3.210 ;
        RECT 2.790 1.125 3.420 1.295 ;
        RECT 3.550 1.125 3.590 2.365 ;
        RECT 2.855 2.195 3.590 2.365 ;
        RECT 3.725 1.535 3.755 1.835 ;
        RECT 3.720 1.535 3.726 1.835 ;
        RECT 3.590 1.410 3.600 2.364 ;
        RECT 3.600 1.420 3.610 2.364 ;
        RECT 3.610 1.430 3.620 2.364 ;
        RECT 3.620 1.440 3.630 2.364 ;
        RECT 3.630 1.450 3.640 2.364 ;
        RECT 3.640 1.460 3.650 2.364 ;
        RECT 3.650 1.470 3.660 2.364 ;
        RECT 3.660 1.480 3.670 2.364 ;
        RECT 3.670 1.490 3.680 2.364 ;
        RECT 3.680 1.500 3.690 2.364 ;
        RECT 3.690 1.510 3.700 2.364 ;
        RECT 3.700 1.520 3.710 2.364 ;
        RECT 3.710 1.530 3.720 2.364 ;
        RECT 3.420 1.125 3.430 1.475 ;
        RECT 3.430 1.125 3.440 1.485 ;
        RECT 3.440 1.125 3.450 1.495 ;
        RECT 3.450 1.125 3.460 1.505 ;
        RECT 3.460 1.125 3.470 1.515 ;
        RECT 3.470 1.125 3.480 1.525 ;
        RECT 3.480 1.125 3.490 1.535 ;
        RECT 3.490 1.125 3.500 1.545 ;
        RECT 3.500 1.125 3.510 1.555 ;
        RECT 3.510 1.125 3.520 1.565 ;
        RECT 3.520 1.125 3.530 1.575 ;
        RECT 3.530 1.125 3.540 1.585 ;
        RECT 3.540 1.125 3.550 1.595 ;
        RECT 1.515 0.885 1.985 1.055 ;
        RECT 1.815 0.885 1.985 2.715 ;
        RECT 1.580 2.405 1.985 2.715 ;
        RECT 1.580 2.545 4.490 2.715 ;
        RECT 4.320 1.405 4.490 2.760 ;
        RECT 4.345 0.960 4.515 1.575 ;
        RECT 4.320 1.405 4.515 1.575 ;
        RECT 6.510 0.960 6.715 1.260 ;
        RECT 6.545 0.960 6.715 2.115 ;
        RECT 6.375 1.945 6.715 2.115 ;
        RECT 6.545 1.565 7.275 1.735 ;
        RECT 5.045 0.960 5.215 2.465 ;
        RECT 5.020 2.140 5.215 2.465 ;
        RECT 7.075 2.090 7.245 2.465 ;
        RECT 5.020 2.295 7.245 2.465 ;
        RECT 7.470 1.680 7.640 2.260 ;
        RECT 7.075 2.090 7.640 2.260 ;
        RECT 7.715 1.550 7.885 1.850 ;
        RECT 7.470 1.680 7.885 1.850 ;
        RECT 7.055 0.920 7.225 1.345 ;
        RECT 8.095 0.920 8.265 1.345 ;
        RECT 7.055 1.175 8.265 1.345 ;
        RECT 6.585 0.480 6.885 0.730 ;
        RECT 7.510 0.560 7.810 0.955 ;
        RECT 7.820 2.045 8.045 2.215 ;
        RECT 6.585 0.560 8.615 0.730 ;
        RECT 8.445 0.560 8.615 1.710 ;
        RECT 8.325 1.540 9.210 1.710 ;
        RECT 8.155 1.540 8.165 2.170 ;
        RECT 8.165 1.540 8.175 2.160 ;
        RECT 8.175 1.540 8.185 2.150 ;
        RECT 8.185 1.540 8.195 2.140 ;
        RECT 8.195 1.540 8.205 2.130 ;
        RECT 8.205 1.540 8.215 2.120 ;
        RECT 8.215 1.540 8.225 2.110 ;
        RECT 8.225 1.540 8.235 2.100 ;
        RECT 8.235 1.540 8.245 2.090 ;
        RECT 8.245 1.540 8.255 2.080 ;
        RECT 8.255 1.540 8.265 2.070 ;
        RECT 8.265 1.540 8.275 2.060 ;
        RECT 8.275 1.540 8.285 2.050 ;
        RECT 8.285 1.540 8.295 2.040 ;
        RECT 8.295 1.540 8.305 2.030 ;
        RECT 8.305 1.540 8.315 2.020 ;
        RECT 8.315 1.540 8.325 2.010 ;
        RECT 8.120 1.970 8.130 2.204 ;
        RECT 8.130 1.960 8.140 2.194 ;
        RECT 8.140 1.950 8.150 2.184 ;
        RECT 8.150 1.940 8.156 2.180 ;
        RECT 8.045 2.045 8.055 2.215 ;
        RECT 8.055 2.035 8.065 2.215 ;
        RECT 8.065 2.025 8.075 2.215 ;
        RECT 8.075 2.015 8.085 2.215 ;
        RECT 8.085 2.005 8.095 2.215 ;
        RECT 8.095 1.995 8.105 2.215 ;
        RECT 8.105 1.985 8.115 2.215 ;
        RECT 8.115 1.975 8.121 2.215 ;
        RECT 3.770 1.125 4.105 1.295 ;
        RECT 3.935 0.610 4.105 2.280 ;
        RECT 3.900 1.980 4.105 2.280 ;
        RECT 4.670 1.780 4.840 2.815 ;
        RECT 4.695 0.610 4.865 1.950 ;
        RECT 4.670 1.780 4.865 1.950 ;
        RECT 4.760 2.645 5.060 2.845 ;
        RECT 5.160 0.555 5.460 0.780 ;
        RECT 3.935 0.610 5.460 0.780 ;
        RECT 7.510 2.460 7.680 2.815 ;
        RECT 4.670 2.645 7.680 2.815 ;
        RECT 7.510 2.460 8.135 2.630 ;
        RECT 8.375 2.295 9.190 2.465 ;
        RECT 9.985 1.610 10.155 2.630 ;
        RECT 9.430 2.460 10.155 2.630 ;
        RECT 9.355 2.395 9.365 2.629 ;
        RECT 9.365 2.405 9.375 2.629 ;
        RECT 9.375 2.415 9.385 2.629 ;
        RECT 9.385 2.425 9.395 2.629 ;
        RECT 9.395 2.435 9.405 2.629 ;
        RECT 9.405 2.445 9.415 2.629 ;
        RECT 9.415 2.455 9.425 2.629 ;
        RECT 9.425 2.460 9.431 2.630 ;
        RECT 9.265 2.305 9.275 2.539 ;
        RECT 9.275 2.315 9.285 2.549 ;
        RECT 9.285 2.325 9.295 2.559 ;
        RECT 9.295 2.335 9.305 2.569 ;
        RECT 9.305 2.345 9.315 2.579 ;
        RECT 9.315 2.355 9.325 2.589 ;
        RECT 9.325 2.365 9.335 2.599 ;
        RECT 9.335 2.375 9.345 2.609 ;
        RECT 9.345 2.385 9.355 2.619 ;
        RECT 9.190 2.295 9.200 2.465 ;
        RECT 9.200 2.295 9.210 2.475 ;
        RECT 9.210 2.295 9.220 2.485 ;
        RECT 9.220 2.295 9.230 2.495 ;
        RECT 9.230 2.295 9.240 2.505 ;
        RECT 9.240 2.295 9.250 2.515 ;
        RECT 9.250 2.295 9.260 2.525 ;
        RECT 9.260 2.295 9.266 2.535 ;
        RECT 8.300 2.295 8.310 2.529 ;
        RECT 8.310 2.295 8.320 2.519 ;
        RECT 8.320 2.295 8.330 2.509 ;
        RECT 8.330 2.295 8.340 2.499 ;
        RECT 8.340 2.295 8.350 2.489 ;
        RECT 8.350 2.295 8.360 2.479 ;
        RECT 8.360 2.295 8.370 2.469 ;
        RECT 8.370 2.295 8.376 2.465 ;
        RECT 8.210 2.385 8.220 2.619 ;
        RECT 8.220 2.375 8.230 2.609 ;
        RECT 8.230 2.365 8.240 2.599 ;
        RECT 8.240 2.355 8.250 2.589 ;
        RECT 8.250 2.345 8.260 2.579 ;
        RECT 8.260 2.335 8.270 2.569 ;
        RECT 8.270 2.325 8.280 2.559 ;
        RECT 8.280 2.315 8.290 2.549 ;
        RECT 8.290 2.305 8.300 2.539 ;
        RECT 8.135 2.460 8.145 2.630 ;
        RECT 8.145 2.450 8.155 2.630 ;
        RECT 8.155 2.440 8.165 2.630 ;
        RECT 8.165 2.430 8.175 2.630 ;
        RECT 8.175 2.420 8.185 2.630 ;
        RECT 8.185 2.410 8.195 2.630 ;
        RECT 8.195 2.400 8.205 2.630 ;
        RECT 8.205 2.390 8.211 2.630 ;
        RECT 7.960 3.040 8.300 3.210 ;
        RECT 8.550 2.645 9.035 2.815 ;
        RECT 10.030 1.195 10.240 1.365 ;
        RECT 9.380 2.915 10.335 3.085 ;
        RECT 10.335 1.225 10.345 3.085 ;
        RECT 10.345 1.235 10.355 3.085 ;
        RECT 10.355 1.245 10.365 3.085 ;
        RECT 10.365 1.255 10.375 3.085 ;
        RECT 10.375 1.265 10.385 3.085 ;
        RECT 10.385 1.275 10.395 3.085 ;
        RECT 10.395 1.285 10.405 3.085 ;
        RECT 10.405 1.295 10.415 3.085 ;
        RECT 10.415 1.305 10.425 3.085 ;
        RECT 10.425 1.315 10.435 3.085 ;
        RECT 10.435 1.325 10.445 3.085 ;
        RECT 10.445 1.335 10.455 3.085 ;
        RECT 10.455 1.345 10.465 3.085 ;
        RECT 10.465 1.355 10.475 3.085 ;
        RECT 10.475 1.365 10.485 3.085 ;
        RECT 10.485 1.375 10.495 3.085 ;
        RECT 10.495 1.385 10.505 3.085 ;
        RECT 10.330 1.215 10.336 1.455 ;
        RECT 10.240 1.195 10.250 1.365 ;
        RECT 10.250 1.195 10.260 1.375 ;
        RECT 10.260 1.195 10.270 1.385 ;
        RECT 10.270 1.195 10.280 1.395 ;
        RECT 10.280 1.195 10.290 1.405 ;
        RECT 10.290 1.195 10.300 1.415 ;
        RECT 10.300 1.195 10.310 1.425 ;
        RECT 10.310 1.195 10.320 1.435 ;
        RECT 10.320 1.195 10.330 1.445 ;
        RECT 9.305 2.850 9.315 3.084 ;
        RECT 9.315 2.860 9.325 3.084 ;
        RECT 9.325 2.870 9.335 3.084 ;
        RECT 9.335 2.880 9.345 3.084 ;
        RECT 9.345 2.890 9.355 3.084 ;
        RECT 9.355 2.900 9.365 3.084 ;
        RECT 9.365 2.910 9.375 3.084 ;
        RECT 9.375 2.915 9.381 3.085 ;
        RECT 9.110 2.655 9.120 2.889 ;
        RECT 9.120 2.665 9.130 2.899 ;
        RECT 9.130 2.675 9.140 2.909 ;
        RECT 9.140 2.685 9.150 2.919 ;
        RECT 9.150 2.695 9.160 2.929 ;
        RECT 9.160 2.705 9.170 2.939 ;
        RECT 9.170 2.715 9.180 2.949 ;
        RECT 9.180 2.725 9.190 2.959 ;
        RECT 9.190 2.735 9.200 2.969 ;
        RECT 9.200 2.745 9.210 2.979 ;
        RECT 9.210 2.755 9.220 2.989 ;
        RECT 9.220 2.765 9.230 2.999 ;
        RECT 9.230 2.775 9.240 3.009 ;
        RECT 9.240 2.785 9.250 3.019 ;
        RECT 9.250 2.795 9.260 3.029 ;
        RECT 9.260 2.805 9.270 3.039 ;
        RECT 9.270 2.815 9.280 3.049 ;
        RECT 9.280 2.825 9.290 3.059 ;
        RECT 9.290 2.835 9.300 3.069 ;
        RECT 9.300 2.840 9.306 3.080 ;
        RECT 9.035 2.645 9.045 2.815 ;
        RECT 9.045 2.645 9.055 2.825 ;
        RECT 9.055 2.645 9.065 2.835 ;
        RECT 9.065 2.645 9.075 2.845 ;
        RECT 9.075 2.645 9.085 2.855 ;
        RECT 9.085 2.645 9.095 2.865 ;
        RECT 9.095 2.645 9.105 2.875 ;
        RECT 9.105 2.645 9.111 2.885 ;
        RECT 8.475 2.645 8.485 2.879 ;
        RECT 8.485 2.645 8.495 2.869 ;
        RECT 8.495 2.645 8.505 2.859 ;
        RECT 8.505 2.645 8.515 2.849 ;
        RECT 8.515 2.645 8.525 2.839 ;
        RECT 8.525 2.645 8.535 2.829 ;
        RECT 8.535 2.645 8.545 2.819 ;
        RECT 8.545 2.645 8.551 2.815 ;
        RECT 8.470 2.650 8.476 2.890 ;
        RECT 8.300 2.820 8.310 3.210 ;
        RECT 8.310 2.810 8.320 3.210 ;
        RECT 8.320 2.800 8.330 3.210 ;
        RECT 8.330 2.790 8.340 3.210 ;
        RECT 8.340 2.780 8.350 3.210 ;
        RECT 8.350 2.770 8.360 3.210 ;
        RECT 8.360 2.760 8.370 3.210 ;
        RECT 8.370 2.750 8.380 3.210 ;
        RECT 8.380 2.740 8.390 3.210 ;
        RECT 8.390 2.730 8.400 3.210 ;
        RECT 8.400 2.720 8.410 3.210 ;
        RECT 8.410 2.710 8.420 3.210 ;
        RECT 8.420 2.700 8.430 3.210 ;
        RECT 8.430 2.690 8.440 3.210 ;
        RECT 8.440 2.680 8.450 3.210 ;
        RECT 8.450 2.670 8.460 3.210 ;
        RECT 8.460 2.660 8.470 3.210 ;
        RECT 11.035 1.515 11.205 1.815 ;
        RECT 11.035 1.645 11.975 1.815 ;
        RECT 11.805 0.980 11.975 2.215 ;
        RECT 11.805 0.980 12.105 1.150 ;
        RECT 11.805 2.045 12.375 2.215 ;
        RECT 11.315 0.630 11.485 1.215 ;
        RECT 11.315 0.630 12.525 0.800 ;
        RECT 12.355 0.630 12.525 1.150 ;
        RECT 12.355 0.980 12.655 1.150 ;
        RECT 9.635 0.785 9.805 2.280 ;
        RECT 9.635 0.785 10.375 0.955 ;
        RECT 10.660 0.995 10.855 1.165 ;
        RECT 10.685 0.995 10.855 2.565 ;
        RECT 11.895 2.395 12.195 2.855 ;
        RECT 12.555 1.935 12.725 2.565 ;
        RECT 10.685 2.395 12.725 2.565 ;
        RECT 13.140 1.530 13.310 2.115 ;
        RECT 12.555 1.935 13.310 2.115 ;
        RECT 10.585 0.930 10.595 1.164 ;
        RECT 10.595 0.940 10.605 1.164 ;
        RECT 10.605 0.950 10.615 1.164 ;
        RECT 10.615 0.960 10.625 1.164 ;
        RECT 10.625 0.970 10.635 1.164 ;
        RECT 10.635 0.980 10.645 1.164 ;
        RECT 10.645 0.990 10.655 1.164 ;
        RECT 10.655 0.995 10.661 1.165 ;
        RECT 10.450 0.795 10.460 1.029 ;
        RECT 10.460 0.805 10.470 1.039 ;
        RECT 10.470 0.815 10.480 1.049 ;
        RECT 10.480 0.825 10.490 1.059 ;
        RECT 10.490 0.835 10.500 1.069 ;
        RECT 10.500 0.845 10.510 1.079 ;
        RECT 10.510 0.855 10.520 1.089 ;
        RECT 10.520 0.865 10.530 1.099 ;
        RECT 10.530 0.875 10.540 1.109 ;
        RECT 10.540 0.885 10.550 1.119 ;
        RECT 10.550 0.895 10.560 1.129 ;
        RECT 10.560 0.905 10.570 1.139 ;
        RECT 10.570 0.915 10.580 1.149 ;
        RECT 10.580 0.920 10.586 1.160 ;
        RECT 10.375 0.785 10.385 0.955 ;
        RECT 10.385 0.785 10.395 0.965 ;
        RECT 10.395 0.785 10.405 0.975 ;
        RECT 10.405 0.785 10.415 0.985 ;
        RECT 10.415 0.785 10.425 0.995 ;
        RECT 10.425 0.785 10.435 1.005 ;
        RECT 10.435 0.785 10.445 1.015 ;
        RECT 10.445 0.785 10.451 1.025 ;
  END 
END FFSDQSRHD2XHT

MACRO FFSDQSRHD1XHT
  CLASS  CORE ;
  FOREIGN FFSDQSRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.530 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.190 0.720 13.430 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 1.290 1.605 1.540 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.760 1.560 6.385 1.955 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.520 1.735 0.690 2.100 ;
        RECT 0.815 1.930 1.230 2.360 ;
        RECT 1.400 1.735 1.570 2.100 ;
        RECT 0.520 1.930 1.570 2.100 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.995 ;
        RECT 2.435 -0.300 2.735 0.785 ;
        RECT 3.295 -0.300 3.595 0.745 ;
        RECT 5.970 -0.300 6.270 1.130 ;
        RECT 8.765 -0.300 8.935 1.220 ;
        RECT 10.645 -0.300 10.945 0.795 ;
        RECT 12.605 -0.300 12.905 0.715 ;
        RECT 0.000 -0.300 13.530 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.965 1.550 3.305 2.015 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.290 1.610 2.775 2.015 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 12.275 1.540 12.640 2.015 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 2.905 0.895 3.990 ;
        RECT 2.540 2.895 3.520 3.990 ;
        RECT 6.145 2.995 7.125 3.990 ;
        RECT 8.675 2.995 8.975 3.990 ;
        RECT 10.700 2.315 11.000 3.990 ;
        RECT 12.605 2.975 12.905 3.990 ;
        RECT 0.000 3.390 13.530 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.170 0.340 2.470 ;
        RECT 0.105 0.825 0.275 2.470 ;
        RECT 0.170 2.170 0.340 2.725 ;
        RECT 0.105 0.825 0.405 0.995 ;
        RECT 0.170 2.555 1.305 2.725 ;
        RECT 1.135 2.555 1.305 3.210 ;
        RECT 1.135 3.040 1.995 3.210 ;
        RECT 2.825 1.125 3.750 1.295 ;
        RECT 3.580 1.125 3.750 2.365 ;
        RECT 2.825 2.195 3.750 2.365 ;
        RECT 1.580 0.725 1.750 1.055 ;
        RECT 1.580 0.885 1.985 1.055 ;
        RECT 1.815 0.885 1.985 2.715 ;
        RECT 1.580 2.370 1.985 2.715 ;
        RECT 1.580 2.545 3.730 2.715 ;
        RECT 3.665 2.610 4.615 2.725 ;
        RECT 3.675 2.610 4.615 2.735 ;
        RECT 3.685 2.610 4.615 2.745 ;
        RECT 3.695 2.610 4.615 2.755 ;
        RECT 3.705 2.610 4.615 2.765 ;
        RECT 3.715 2.610 4.615 2.775 ;
        RECT 3.720 2.545 3.730 2.780 ;
        RECT 1.580 2.555 3.740 2.715 ;
        RECT 1.580 2.565 3.750 2.715 ;
        RECT 1.580 2.575 3.760 2.715 ;
        RECT 1.580 2.585 3.770 2.715 ;
        RECT 1.580 2.595 3.780 2.715 ;
        RECT 3.720 2.610 4.615 2.779 ;
        RECT 1.580 2.605 3.790 2.715 ;
        RECT 4.445 0.895 4.615 2.780 ;
        RECT 3.790 2.610 4.615 2.780 ;
        RECT 6.585 0.960 6.755 2.115 ;
        RECT 6.490 0.960 6.790 1.130 ;
        RECT 6.585 1.500 7.360 1.670 ;
        RECT 5.145 0.895 5.315 2.465 ;
        RECT 7.540 1.680 7.710 2.465 ;
        RECT 5.145 2.295 7.710 2.465 ;
        RECT 7.775 1.550 7.945 1.850 ;
        RECT 7.540 1.680 7.945 1.850 ;
        RECT 7.000 0.960 7.300 1.230 ;
        RECT 7.000 1.060 8.235 1.230 ;
        RECT 8.065 1.060 8.235 1.360 ;
        RECT 6.630 0.480 6.930 0.695 ;
        RECT 7.890 2.045 8.015 2.215 ;
        RECT 8.125 1.580 8.190 2.215 ;
        RECT 6.630 0.525 8.585 0.695 ;
        RECT 8.415 0.525 8.585 1.750 ;
        RECT 8.295 1.580 9.180 1.750 ;
        RECT 8.190 1.580 8.200 2.104 ;
        RECT 8.200 1.580 8.210 2.094 ;
        RECT 8.210 1.580 8.220 2.084 ;
        RECT 8.220 1.580 8.230 2.074 ;
        RECT 8.230 1.580 8.240 2.064 ;
        RECT 8.240 1.580 8.250 2.054 ;
        RECT 8.250 1.580 8.260 2.044 ;
        RECT 8.260 1.580 8.270 2.034 ;
        RECT 8.270 1.580 8.280 2.024 ;
        RECT 8.280 1.580 8.290 2.014 ;
        RECT 8.290 1.580 8.296 2.010 ;
        RECT 8.015 2.045 8.025 2.215 ;
        RECT 8.025 2.035 8.035 2.215 ;
        RECT 8.035 2.025 8.045 2.215 ;
        RECT 8.045 2.015 8.055 2.215 ;
        RECT 8.055 2.005 8.065 2.215 ;
        RECT 8.065 1.995 8.075 2.215 ;
        RECT 8.075 1.985 8.085 2.215 ;
        RECT 8.085 1.975 8.095 2.215 ;
        RECT 8.095 1.965 8.105 2.215 ;
        RECT 8.105 1.955 8.115 2.215 ;
        RECT 8.115 1.945 8.125 2.215 ;
        RECT 3.930 0.545 4.100 2.430 ;
        RECT 4.795 0.545 4.965 2.835 ;
        RECT 3.930 0.545 5.560 0.715 ;
        RECT 4.795 2.645 8.020 2.815 ;
        RECT 8.445 2.295 9.205 2.465 ;
        RECT 9.380 2.395 10.105 2.565 ;
        RECT 9.935 2.395 10.105 2.770 ;
        RECT 9.305 2.330 9.315 2.564 ;
        RECT 9.315 2.340 9.325 2.564 ;
        RECT 9.325 2.350 9.335 2.564 ;
        RECT 9.335 2.360 9.345 2.564 ;
        RECT 9.345 2.370 9.355 2.564 ;
        RECT 9.355 2.380 9.365 2.564 ;
        RECT 9.365 2.390 9.375 2.564 ;
        RECT 9.375 2.395 9.381 2.565 ;
        RECT 9.280 2.305 9.290 2.539 ;
        RECT 9.290 2.315 9.300 2.549 ;
        RECT 9.300 2.320 9.306 2.560 ;
        RECT 9.205 2.295 9.215 2.465 ;
        RECT 9.215 2.295 9.225 2.475 ;
        RECT 9.225 2.295 9.235 2.485 ;
        RECT 9.235 2.295 9.245 2.495 ;
        RECT 9.245 2.295 9.255 2.505 ;
        RECT 9.255 2.295 9.265 2.515 ;
        RECT 9.265 2.295 9.275 2.525 ;
        RECT 9.275 2.295 9.281 2.535 ;
        RECT 8.370 2.295 8.380 2.529 ;
        RECT 8.380 2.295 8.390 2.519 ;
        RECT 8.390 2.295 8.400 2.509 ;
        RECT 8.400 2.295 8.410 2.499 ;
        RECT 8.410 2.295 8.420 2.489 ;
        RECT 8.420 2.295 8.430 2.479 ;
        RECT 8.430 2.295 8.440 2.469 ;
        RECT 8.440 2.295 8.446 2.465 ;
        RECT 8.095 2.570 8.105 2.804 ;
        RECT 8.105 2.560 8.115 2.794 ;
        RECT 8.115 2.550 8.125 2.784 ;
        RECT 8.125 2.540 8.135 2.774 ;
        RECT 8.135 2.530 8.145 2.764 ;
        RECT 8.145 2.520 8.155 2.754 ;
        RECT 8.155 2.510 8.165 2.744 ;
        RECT 8.165 2.500 8.175 2.734 ;
        RECT 8.175 2.490 8.185 2.724 ;
        RECT 8.185 2.480 8.195 2.714 ;
        RECT 8.195 2.470 8.205 2.704 ;
        RECT 8.205 2.460 8.215 2.694 ;
        RECT 8.215 2.450 8.225 2.684 ;
        RECT 8.225 2.440 8.235 2.674 ;
        RECT 8.235 2.430 8.245 2.664 ;
        RECT 8.245 2.420 8.255 2.654 ;
        RECT 8.255 2.410 8.265 2.644 ;
        RECT 8.265 2.400 8.275 2.634 ;
        RECT 8.275 2.390 8.285 2.624 ;
        RECT 8.285 2.380 8.295 2.614 ;
        RECT 8.295 2.370 8.305 2.604 ;
        RECT 8.305 2.360 8.315 2.594 ;
        RECT 8.315 2.350 8.325 2.584 ;
        RECT 8.325 2.340 8.335 2.574 ;
        RECT 8.335 2.330 8.345 2.564 ;
        RECT 8.345 2.320 8.355 2.554 ;
        RECT 8.355 2.310 8.365 2.544 ;
        RECT 8.365 2.300 8.371 2.540 ;
        RECT 8.020 2.645 8.030 2.815 ;
        RECT 8.030 2.635 8.040 2.815 ;
        RECT 8.040 2.625 8.050 2.815 ;
        RECT 8.050 2.615 8.060 2.815 ;
        RECT 8.060 2.605 8.070 2.815 ;
        RECT 8.070 2.595 8.080 2.815 ;
        RECT 8.080 2.585 8.090 2.815 ;
        RECT 8.090 2.575 8.096 2.815 ;
        RECT 7.960 3.040 8.325 3.210 ;
        RECT 8.595 2.645 9.050 2.815 ;
        RECT 9.225 2.745 9.665 2.915 ;
        RECT 9.495 2.745 9.665 3.120 ;
        RECT 9.955 1.270 10.255 1.440 ;
        RECT 10.085 1.270 10.255 1.825 ;
        RECT 10.085 1.655 10.455 1.825 ;
        RECT 10.285 1.655 10.455 3.120 ;
        RECT 9.495 2.950 10.455 3.120 ;
        RECT 9.150 2.680 9.160 2.914 ;
        RECT 9.160 2.690 9.170 2.914 ;
        RECT 9.170 2.700 9.180 2.914 ;
        RECT 9.180 2.710 9.190 2.914 ;
        RECT 9.190 2.720 9.200 2.914 ;
        RECT 9.200 2.730 9.210 2.914 ;
        RECT 9.210 2.740 9.220 2.914 ;
        RECT 9.220 2.745 9.226 2.915 ;
        RECT 9.125 2.655 9.135 2.889 ;
        RECT 9.135 2.665 9.145 2.899 ;
        RECT 9.145 2.670 9.151 2.910 ;
        RECT 9.050 2.645 9.060 2.815 ;
        RECT 9.060 2.645 9.070 2.825 ;
        RECT 9.070 2.645 9.080 2.835 ;
        RECT 9.080 2.645 9.090 2.845 ;
        RECT 9.090 2.645 9.100 2.855 ;
        RECT 9.100 2.645 9.110 2.865 ;
        RECT 9.110 2.645 9.120 2.875 ;
        RECT 9.120 2.645 9.126 2.885 ;
        RECT 8.520 2.645 8.530 2.879 ;
        RECT 8.530 2.645 8.540 2.869 ;
        RECT 8.540 2.645 8.550 2.859 ;
        RECT 8.550 2.645 8.560 2.849 ;
        RECT 8.560 2.645 8.570 2.839 ;
        RECT 8.570 2.645 8.580 2.829 ;
        RECT 8.580 2.645 8.590 2.819 ;
        RECT 8.590 2.645 8.596 2.815 ;
        RECT 8.495 2.670 8.505 2.904 ;
        RECT 8.505 2.660 8.515 2.894 ;
        RECT 8.515 2.650 8.521 2.890 ;
        RECT 8.325 2.840 8.335 3.210 ;
        RECT 8.335 2.830 8.345 3.210 ;
        RECT 8.345 2.820 8.355 3.210 ;
        RECT 8.355 2.810 8.365 3.210 ;
        RECT 8.365 2.800 8.375 3.210 ;
        RECT 8.375 2.790 8.385 3.210 ;
        RECT 8.385 2.780 8.395 3.210 ;
        RECT 8.395 2.770 8.405 3.210 ;
        RECT 8.405 2.760 8.415 3.210 ;
        RECT 8.415 2.750 8.425 3.210 ;
        RECT 8.425 2.740 8.435 3.210 ;
        RECT 8.435 2.730 8.445 3.210 ;
        RECT 8.445 2.720 8.455 3.210 ;
        RECT 8.455 2.710 8.465 3.210 ;
        RECT 8.465 2.700 8.475 3.210 ;
        RECT 8.475 2.690 8.485 3.210 ;
        RECT 8.485 2.680 8.495 3.210 ;
        RECT 10.985 1.460 11.155 1.760 ;
        RECT 11.595 1.110 11.895 1.630 ;
        RECT 10.985 1.460 11.895 1.630 ;
        RECT 11.725 1.110 11.895 2.405 ;
        RECT 11.725 2.235 12.295 2.405 ;
        RECT 11.205 0.760 11.375 1.280 ;
        RECT 11.075 1.110 11.375 1.280 ;
        RECT 11.205 0.760 12.285 0.930 ;
        RECT 12.115 0.760 12.285 1.280 ;
        RECT 12.115 1.110 12.415 1.280 ;
        RECT 9.545 0.900 9.715 2.215 ;
        RECT 9.545 2.045 9.845 2.215 ;
        RECT 9.545 0.900 10.330 1.070 ;
        RECT 10.565 1.060 10.805 1.230 ;
        RECT 10.635 1.060 10.805 2.110 ;
        RECT 10.635 1.940 11.390 2.110 ;
        RECT 11.220 1.940 11.390 2.795 ;
        RECT 11.815 2.625 12.115 2.855 ;
        RECT 12.840 1.610 13.010 2.795 ;
        RECT 11.220 2.625 13.010 2.795 ;
        RECT 10.490 0.995 10.500 1.229 ;
        RECT 10.500 1.005 10.510 1.229 ;
        RECT 10.510 1.015 10.520 1.229 ;
        RECT 10.520 1.025 10.530 1.229 ;
        RECT 10.530 1.035 10.540 1.229 ;
        RECT 10.540 1.045 10.550 1.229 ;
        RECT 10.550 1.055 10.560 1.229 ;
        RECT 10.560 1.060 10.566 1.230 ;
        RECT 10.405 0.910 10.415 1.144 ;
        RECT 10.415 0.920 10.425 1.154 ;
        RECT 10.425 0.930 10.435 1.164 ;
        RECT 10.435 0.940 10.445 1.174 ;
        RECT 10.445 0.950 10.455 1.184 ;
        RECT 10.455 0.960 10.465 1.194 ;
        RECT 10.465 0.970 10.475 1.204 ;
        RECT 10.475 0.980 10.485 1.214 ;
        RECT 10.485 0.985 10.491 1.225 ;
        RECT 10.330 0.900 10.340 1.070 ;
        RECT 10.340 0.900 10.350 1.080 ;
        RECT 10.350 0.900 10.360 1.090 ;
        RECT 10.360 0.900 10.370 1.100 ;
        RECT 10.370 0.900 10.380 1.110 ;
        RECT 10.380 0.900 10.390 1.120 ;
        RECT 10.390 0.900 10.400 1.130 ;
        RECT 10.400 0.900 10.406 1.140 ;
  END 
END FFSDQSRHD1XHT

MACRO FFSDQSHDMXHT
  CLASS  CORE ;
  FOREIGN FFSDQSHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.480 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.140 1.060 11.380 1.360 ;
        RECT 11.170 1.060 11.380 2.435 ;
        RECT 11.140 1.980 11.380 2.435 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.595 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.425 -0.300 2.725 0.595 ;
        RECT 3.355 -0.300 3.655 0.595 ;
        RECT 6.035 -0.300 6.335 0.745 ;
        RECT 7.275 -0.300 7.445 0.850 ;
        RECT 9.260 -0.300 9.430 0.640 ;
        RECT 10.555 -0.300 10.855 1.145 ;
        RECT 0.000 -0.300 11.480 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.850 1.525 3.340 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.640 0.520 7.810 1.910 ;
        RECT 6.995 1.610 7.810 1.910 ;
        RECT 7.640 0.520 9.015 0.690 ;
        RECT 8.845 0.520 9.015 1.145 ;
        RECT 9.705 0.540 9.875 1.145 ;
        RECT 8.845 0.920 9.875 1.145 ;
        RECT 9.705 0.540 10.165 0.710 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.355 2.735 2.655 3.990 ;
        RECT 3.235 2.675 3.405 3.990 ;
        RECT 5.965 3.160 6.265 3.990 ;
        RECT 7.175 3.160 7.475 3.990 ;
        RECT 9.280 2.770 9.450 3.990 ;
        RECT 9.920 2.880 10.090 3.990 ;
        RECT 10.590 2.770 10.760 3.990 ;
        RECT 0.000 3.390 11.480 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.525 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.150 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.975 0.775 2.145 1.035 ;
        RECT 1.530 0.865 2.145 1.035 ;
        RECT 1.975 0.775 4.620 0.945 ;
        RECT 4.450 0.775 4.620 2.280 ;
        RECT 5.150 0.900 5.320 2.280 ;
        RECT 5.150 1.600 6.465 1.770 ;
        RECT 6.645 1.060 6.815 2.215 ;
        RECT 6.515 2.045 6.815 2.215 ;
        RECT 6.645 1.060 7.460 1.360 ;
        RECT 2.835 1.125 3.695 1.295 ;
        RECT 2.815 2.190 3.755 2.360 ;
        RECT 3.525 1.125 3.695 2.360 ;
        RECT 3.585 1.525 3.755 2.980 ;
        RECT 3.525 1.525 3.820 1.825 ;
        RECT 3.585 2.810 8.155 2.980 ;
        RECT 3.875 1.125 4.195 1.295 ;
        RECT 3.940 1.980 4.195 2.280 ;
        RECT 4.000 1.125 4.195 2.630 ;
        RECT 4.800 0.535 4.970 2.630 ;
        RECT 4.800 0.535 5.595 0.705 ;
        RECT 7.990 1.645 8.160 2.630 ;
        RECT 8.020 1.245 8.190 1.815 ;
        RECT 7.990 1.645 8.190 1.815 ;
        RECT 4.000 2.460 8.830 2.630 ;
        RECT 8.660 2.460 8.830 2.760 ;
        RECT 9.015 1.325 10.280 1.495 ;
        RECT 10.110 0.890 10.280 2.215 ;
        RECT 9.795 2.045 10.280 2.215 ;
        RECT 8.415 0.870 8.585 2.215 ;
        RECT 8.295 0.870 8.595 1.040 ;
        RECT 8.340 2.045 8.640 2.215 ;
        RECT 9.120 1.675 9.290 2.590 ;
        RECT 8.415 1.675 9.795 1.845 ;
        RECT 10.790 1.610 10.960 2.590 ;
        RECT 9.120 2.420 10.960 2.590 ;
        RECT 10.790 1.610 10.970 1.910 ;
  END 
END FFSDQSHDMXHT

MACRO FFSDQSHDLXHT
  CLASS  CORE ;
  FOREIGN FFSDQSHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.070 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.535 1.060 10.970 1.360 ;
        RECT 10.760 1.060 10.970 2.480 ;
        RECT 10.730 1.980 10.970 2.480 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.525 2.980 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.435 -0.300 2.735 0.595 ;
        RECT 3.325 -0.300 3.625 0.595 ;
        RECT 5.945 -0.300 6.245 0.745 ;
        RECT 7.150 -0.300 7.320 0.850 ;
        RECT 9.105 -0.300 9.275 0.640 ;
        RECT 10.470 -0.300 10.770 0.655 ;
        RECT 0.000 -0.300 11.070 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.760 1.525 3.250 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.040 1.290 2.440 1.800 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.560 0.520 7.730 1.910 ;
        RECT 6.885 1.610 7.730 1.910 ;
        RECT 7.560 0.520 8.890 0.690 ;
        RECT 8.720 0.520 8.890 1.145 ;
        RECT 9.580 0.540 9.750 1.145 ;
        RECT 8.720 0.920 9.750 1.145 ;
        RECT 9.580 0.540 10.010 0.710 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.620 2.715 3.260 3.990 ;
        RECT 5.855 3.160 6.155 3.990 ;
        RECT 7.085 3.160 7.385 3.990 ;
        RECT 9.090 2.770 9.390 3.990 ;
        RECT 10.115 2.770 10.415 3.990 ;
        RECT 0.000 3.390 11.070 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.525 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 2.930 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.530 0.865 1.720 1.185 ;
        RECT 1.750 0.775 1.920 1.035 ;
        RECT 1.530 0.865 1.920 1.035 ;
        RECT 1.750 0.775 4.530 0.945 ;
        RECT 4.360 0.775 4.530 2.280 ;
        RECT 5.060 0.900 5.230 2.280 ;
        RECT 5.060 1.595 6.355 1.765 ;
        RECT 6.535 1.060 6.705 2.215 ;
        RECT 6.405 2.045 6.705 2.215 ;
        RECT 6.535 1.060 7.380 1.360 ;
        RECT 2.745 1.125 3.605 1.295 ;
        RECT 2.775 2.190 3.635 2.360 ;
        RECT 3.435 1.125 3.605 2.360 ;
        RECT 3.465 1.525 3.635 2.980 ;
        RECT 3.435 1.525 3.730 1.825 ;
        RECT 3.465 2.810 8.030 2.980 ;
        RECT 3.785 1.125 4.105 1.295 ;
        RECT 3.935 1.125 4.105 2.630 ;
        RECT 3.815 2.395 4.105 2.630 ;
        RECT 4.710 0.535 4.880 2.630 ;
        RECT 4.710 0.535 5.505 0.705 ;
        RECT 7.910 1.210 8.080 2.630 ;
        RECT 3.815 2.460 8.690 2.630 ;
        RECT 8.520 2.460 8.690 2.760 ;
        RECT 8.860 1.325 10.155 1.495 ;
        RECT 9.985 0.890 10.155 2.215 ;
        RECT 9.655 2.045 10.155 2.215 ;
        RECT 8.140 0.870 8.460 1.040 ;
        RECT 8.290 0.870 8.460 2.280 ;
        RECT 8.290 1.675 8.465 2.280 ;
        RECT 8.995 1.675 9.165 2.590 ;
        RECT 8.290 1.675 9.640 1.845 ;
        RECT 10.380 1.560 10.550 2.590 ;
        RECT 8.995 2.420 10.550 2.590 ;
        RECT 10.380 1.560 10.580 1.860 ;
  END 
END FFSDQSHDLXHT

MACRO FFSDQSHD2XHT
  CLASS  CORE ;
  FOREIGN FFSDQSHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.300 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.440 0.720 11.610 2.960 ;
        RECT 11.440 1.650 11.790 2.015 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.265 -0.300 2.565 0.595 ;
        RECT 3.325 -0.300 3.625 0.595 ;
        RECT 5.885 -0.300 6.185 0.905 ;
        RECT 7.375 -0.300 7.675 0.715 ;
        RECT 9.350 -0.300 9.650 0.795 ;
        RECT 10.855 -0.300 11.155 1.055 ;
        RECT 11.895 -0.300 12.195 1.055 ;
        RECT 0.000 -0.300 12.300 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.730 1.525 3.220 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.265 0.960 7.435 1.565 ;
        RECT 7.160 1.265 7.435 1.565 ;
        RECT 7.855 0.590 8.025 1.130 ;
        RECT 7.265 0.960 8.025 1.130 ;
        RECT 7.855 0.590 9.140 0.760 ;
        RECT 8.970 0.590 9.140 1.145 ;
        RECT 9.860 0.920 10.230 1.145 ;
        RECT 10.060 0.525 10.230 1.145 ;
        RECT 8.970 0.975 10.230 1.145 ;
        RECT 10.060 0.525 10.415 0.695 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.620 2.780 3.260 3.990 ;
        RECT 5.910 3.095 6.210 3.990 ;
        RECT 7.010 3.095 7.650 3.990 ;
        RECT 9.505 2.850 9.805 3.990 ;
        RECT 10.515 2.975 11.155 3.990 ;
        RECT 11.895 2.295 12.195 3.990 ;
        RECT 0.000 3.390 12.300 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.575 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.150 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.945 0.775 2.115 1.035 ;
        RECT 1.530 0.865 2.115 1.035 ;
        RECT 1.945 0.775 4.500 0.945 ;
        RECT 4.330 0.775 4.500 2.280 ;
        RECT 5.030 0.910 5.200 2.280 ;
        RECT 6.120 1.675 6.420 1.865 ;
        RECT 5.030 1.695 6.420 1.865 ;
        RECT 5.625 1.245 5.925 1.515 ;
        RECT 5.625 1.245 6.980 1.415 ;
        RECT 6.810 0.670 6.980 2.215 ;
        RECT 6.460 2.045 6.980 2.215 ;
        RECT 6.810 0.670 7.030 0.970 ;
        RECT 7.655 1.610 7.825 1.915 ;
        RECT 6.810 1.745 7.825 1.915 ;
        RECT 2.775 1.125 3.575 1.295 ;
        RECT 2.775 2.190 3.635 2.360 ;
        RECT 3.405 1.125 3.575 2.360 ;
        RECT 3.465 1.525 3.635 3.035 ;
        RECT 3.405 1.525 3.700 1.825 ;
        RECT 3.465 2.865 5.525 3.035 ;
        RECT 5.765 2.745 8.115 2.915 ;
        RECT 7.935 2.745 8.115 3.185 ;
        RECT 7.935 3.015 8.910 3.185 ;
        RECT 5.645 2.745 5.655 3.025 ;
        RECT 5.655 2.745 5.665 3.015 ;
        RECT 5.665 2.745 5.675 3.005 ;
        RECT 5.675 2.745 5.685 2.995 ;
        RECT 5.685 2.745 5.695 2.985 ;
        RECT 5.695 2.745 5.705 2.975 ;
        RECT 5.705 2.745 5.715 2.965 ;
        RECT 5.715 2.745 5.725 2.955 ;
        RECT 5.725 2.745 5.735 2.945 ;
        RECT 5.735 2.745 5.745 2.935 ;
        RECT 5.745 2.745 5.755 2.925 ;
        RECT 5.755 2.745 5.765 2.915 ;
        RECT 5.525 2.865 5.535 3.035 ;
        RECT 5.535 2.855 5.545 3.035 ;
        RECT 5.545 2.845 5.555 3.035 ;
        RECT 5.555 2.835 5.565 3.035 ;
        RECT 5.565 2.825 5.575 3.035 ;
        RECT 5.575 2.815 5.585 3.035 ;
        RECT 5.585 2.805 5.595 3.035 ;
        RECT 5.595 2.795 5.605 3.035 ;
        RECT 5.605 2.785 5.615 3.035 ;
        RECT 5.615 2.775 5.625 3.035 ;
        RECT 5.625 2.765 5.635 3.035 ;
        RECT 5.635 2.755 5.645 3.035 ;
        RECT 3.755 1.125 4.075 1.295 ;
        RECT 3.905 1.125 4.075 2.685 ;
        RECT 3.820 1.980 4.075 2.685 ;
        RECT 4.680 0.535 4.850 2.685 ;
        RECT 3.820 2.515 5.265 2.685 ;
        RECT 4.680 0.535 5.445 0.705 ;
        RECT 8.135 1.290 8.305 2.565 ;
        RECT 5.505 2.395 9.000 2.565 ;
        RECT 8.830 2.395 9.000 2.770 ;
        RECT 5.385 2.395 5.395 2.675 ;
        RECT 5.395 2.395 5.405 2.665 ;
        RECT 5.405 2.395 5.415 2.655 ;
        RECT 5.415 2.395 5.425 2.645 ;
        RECT 5.425 2.395 5.435 2.635 ;
        RECT 5.435 2.395 5.445 2.625 ;
        RECT 5.445 2.395 5.455 2.615 ;
        RECT 5.455 2.395 5.465 2.605 ;
        RECT 5.465 2.395 5.475 2.595 ;
        RECT 5.475 2.395 5.485 2.585 ;
        RECT 5.485 2.395 5.495 2.575 ;
        RECT 5.495 2.395 5.505 2.565 ;
        RECT 5.265 2.515 5.275 2.685 ;
        RECT 5.275 2.505 5.285 2.685 ;
        RECT 5.285 2.495 5.295 2.685 ;
        RECT 5.295 2.485 5.305 2.685 ;
        RECT 5.305 2.475 5.315 2.685 ;
        RECT 5.315 2.465 5.325 2.685 ;
        RECT 5.325 2.455 5.335 2.685 ;
        RECT 5.335 2.445 5.345 2.685 ;
        RECT 5.345 2.435 5.355 2.685 ;
        RECT 5.355 2.425 5.365 2.685 ;
        RECT 5.365 2.415 5.375 2.685 ;
        RECT 5.375 2.405 5.385 2.685 ;
        RECT 8.975 1.325 10.580 1.495 ;
        RECT 10.410 0.875 10.580 2.215 ;
        RECT 10.065 2.045 10.580 2.215 ;
        RECT 8.265 0.940 8.730 1.110 ;
        RECT 8.560 0.940 8.730 2.215 ;
        RECT 8.560 1.675 8.795 2.215 ;
        RECT 8.560 2.045 8.860 2.215 ;
        RECT 8.560 1.675 9.805 1.845 ;
        RECT 9.635 1.675 9.805 2.610 ;
        RECT 9.950 2.440 10.120 2.740 ;
        RECT 11.090 1.610 11.260 2.610 ;
        RECT 9.635 2.440 11.260 2.610 ;
  END 
END FFSDQSHD2XHT

MACRO FFSDQRHDMXHT
  CLASS  CORE ;
  FOREIGN FFSDQRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.300 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.960 1.060 12.200 2.455 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.960 1.610 8.510 2.010 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.415 -0.300 2.715 0.595 ;
        RECT 3.325 -0.300 3.625 0.595 ;
        RECT 5.945 -0.300 6.245 1.145 ;
        RECT 6.985 -0.300 7.285 0.595 ;
        RECT 8.055 -0.300 8.225 0.810 ;
        RECT 9.995 -0.300 10.295 0.525 ;
        RECT 11.410 -0.300 11.580 1.210 ;
        RECT 0.000 -0.300 12.300 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.740 1.525 3.230 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.625 2.740 3.265 3.990 ;
        RECT 5.965 3.195 6.265 3.990 ;
        RECT 8.095 3.195 8.395 3.990 ;
        RECT 10.035 2.810 10.335 3.990 ;
        RECT 11.345 2.745 11.645 3.990 ;
        RECT 0.000 3.390 12.300 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.555 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.005 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.980 0.775 2.150 1.035 ;
        RECT 1.530 0.865 2.150 1.035 ;
        RECT 1.980 0.775 4.510 0.945 ;
        RECT 4.275 0.585 4.510 0.945 ;
        RECT 4.340 0.585 4.510 2.280 ;
        RECT 4.340 1.960 4.520 2.280 ;
        RECT 4.340 1.970 4.530 2.280 ;
        RECT 4.340 1.980 4.540 2.280 ;
        RECT 5.070 0.910 5.210 2.280 ;
        RECT 6.165 1.675 6.465 1.865 ;
        RECT 5.390 1.695 6.465 1.865 ;
        RECT 5.240 1.555 5.250 1.865 ;
        RECT 5.250 1.565 5.260 1.865 ;
        RECT 5.260 1.575 5.270 1.865 ;
        RECT 5.270 1.585 5.280 1.865 ;
        RECT 5.280 1.595 5.290 1.865 ;
        RECT 5.290 1.605 5.300 1.865 ;
        RECT 5.300 1.615 5.310 1.865 ;
        RECT 5.310 1.625 5.320 1.865 ;
        RECT 5.320 1.635 5.330 1.865 ;
        RECT 5.330 1.645 5.340 1.865 ;
        RECT 5.340 1.655 5.350 1.865 ;
        RECT 5.350 1.665 5.360 1.865 ;
        RECT 5.360 1.675 5.370 1.865 ;
        RECT 5.370 1.685 5.380 1.865 ;
        RECT 5.380 1.695 5.390 1.865 ;
        RECT 5.210 1.525 5.220 2.279 ;
        RECT 5.220 1.535 5.230 2.279 ;
        RECT 5.230 1.545 5.240 2.279 ;
        RECT 5.040 0.910 5.050 1.640 ;
        RECT 5.050 0.910 5.060 1.650 ;
        RECT 5.060 0.910 5.070 1.660 ;
        RECT 5.685 1.325 5.985 1.515 ;
        RECT 6.580 0.775 6.815 1.495 ;
        RECT 5.685 1.325 6.815 1.495 ;
        RECT 6.645 0.775 6.815 2.215 ;
        RECT 6.645 2.045 7.185 2.215 ;
        RECT 7.470 0.480 7.640 0.945 ;
        RECT 6.580 0.775 7.640 0.945 ;
        RECT 2.805 1.125 3.585 1.295 ;
        RECT 2.785 2.190 3.645 2.360 ;
        RECT 3.415 1.125 3.585 2.360 ;
        RECT 3.475 1.525 3.645 2.985 ;
        RECT 3.415 1.525 3.730 1.825 ;
        RECT 8.390 2.745 8.560 2.985 ;
        RECT 3.475 2.815 8.560 2.985 ;
        RECT 8.390 2.745 9.135 2.915 ;
        RECT 3.860 1.980 4.145 2.280 ;
        RECT 3.845 1.125 4.145 1.295 ;
        RECT 3.975 1.125 4.145 2.635 ;
        RECT 3.915 1.980 4.145 2.635 ;
        RECT 4.700 1.755 4.890 1.829 ;
        RECT 4.710 1.755 4.890 1.839 ;
        RECT 4.690 0.535 4.860 1.819 ;
        RECT 4.690 1.735 4.870 1.819 ;
        RECT 4.690 1.745 4.880 1.819 ;
        RECT 4.720 1.755 4.890 2.635 ;
        RECT 4.690 0.535 5.485 0.705 ;
        RECT 8.035 2.395 8.205 2.635 ;
        RECT 3.915 2.465 8.205 2.635 ;
        RECT 8.775 1.330 8.945 2.565 ;
        RECT 8.755 1.330 9.055 1.500 ;
        RECT 8.035 2.395 9.650 2.565 ;
        RECT 9.480 2.395 9.650 2.795 ;
        RECT 6.995 1.590 7.740 1.760 ;
        RECT 7.570 1.125 7.740 2.280 ;
        RECT 8.405 0.605 8.575 1.295 ;
        RECT 7.545 1.125 8.575 1.295 ;
        RECT 9.620 0.605 9.790 0.945 ;
        RECT 8.405 0.605 9.790 0.775 ;
        RECT 9.620 0.775 11.200 0.945 ;
        RECT 11.030 0.775 11.200 1.745 ;
        RECT 9.850 1.125 10.020 1.560 ;
        RECT 9.850 1.125 10.850 1.295 ;
        RECT 10.680 1.125 10.850 2.215 ;
        RECT 10.680 2.045 11.255 2.215 ;
        RECT 9.045 0.955 9.405 1.125 ;
        RECT 9.235 0.955 9.405 2.215 ;
        RECT 9.150 2.045 10.500 2.215 ;
        RECT 10.330 1.610 10.500 2.565 ;
        RECT 11.610 1.560 11.780 2.565 ;
        RECT 10.330 2.395 11.780 2.565 ;
  END 
END FFSDQRHDMXHT

MACRO FFSDQRHDLXHT
  CLASS  CORE ;
  FOREIGN FFSDQRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.300 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.960 1.060 12.200 2.440 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.960 1.535 8.510 2.010 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.350 2.980 ;
        RECT 1.180 2.810 1.350 3.110 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.435 -0.300 2.735 0.595 ;
        RECT 3.405 -0.300 3.705 0.595 ;
        RECT 5.905 -0.300 6.205 0.675 ;
        RECT 6.985 -0.300 7.285 0.595 ;
        RECT 8.055 -0.300 8.225 0.810 ;
        RECT 9.995 -0.300 10.295 0.525 ;
        RECT 11.410 -0.300 11.580 1.360 ;
        RECT 0.000 -0.300 12.300 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.790 1.525 3.280 1.950 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.830 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.630 2.660 3.270 3.990 ;
        RECT 5.965 3.195 6.265 3.990 ;
        RECT 8.095 3.195 8.395 3.990 ;
        RECT 10.035 2.810 10.335 3.990 ;
        RECT 11.345 2.810 11.645 3.990 ;
        RECT 0.000 3.390 12.300 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.555 0.650 ;
        RECT 1.180 2.460 1.880 2.630 ;
        RECT 1.710 2.460 1.880 2.825 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.530 0.865 1.720 1.185 ;
        RECT 2.005 0.775 2.175 1.035 ;
        RECT 1.530 0.865 2.175 1.035 ;
        RECT 2.005 0.775 4.590 0.945 ;
        RECT 4.355 0.645 4.590 0.945 ;
        RECT 4.420 0.645 4.590 2.280 ;
        RECT 5.120 0.900 5.290 2.280 ;
        RECT 6.225 1.675 6.525 1.865 ;
        RECT 5.120 1.695 6.525 1.865 ;
        RECT 5.745 1.325 6.045 1.515 ;
        RECT 6.550 0.775 6.875 1.495 ;
        RECT 5.745 1.325 6.875 1.495 ;
        RECT 6.705 0.775 6.875 2.215 ;
        RECT 6.705 2.045 7.185 2.215 ;
        RECT 7.470 0.480 7.640 0.945 ;
        RECT 6.550 0.775 7.640 0.945 ;
        RECT 2.825 1.125 3.635 1.295 ;
        RECT 2.805 2.130 3.665 2.300 ;
        RECT 3.465 1.125 3.635 2.300 ;
        RECT 3.495 1.525 3.665 3.015 ;
        RECT 3.465 1.525 3.760 1.825 ;
        RECT 8.390 2.745 8.560 3.015 ;
        RECT 3.495 2.845 8.560 3.015 ;
        RECT 8.390 2.745 8.975 2.915 ;
        RECT 3.975 1.125 4.145 2.635 ;
        RECT 3.845 2.400 4.145 2.635 ;
        RECT 3.865 1.125 4.165 1.295 ;
        RECT 4.770 0.535 4.940 2.635 ;
        RECT 4.770 0.535 5.565 0.705 ;
        RECT 8.035 2.395 8.205 2.635 ;
        RECT 3.845 2.465 8.205 2.635 ;
        RECT 8.755 1.330 8.925 2.565 ;
        RECT 8.755 1.330 9.055 1.500 ;
        RECT 9.415 2.395 9.650 2.595 ;
        RECT 8.035 2.395 9.650 2.565 ;
        RECT 9.415 2.425 9.715 2.595 ;
        RECT 7.055 1.585 7.740 1.755 ;
        RECT 7.570 1.125 7.740 2.280 ;
        RECT 8.405 0.605 8.575 1.295 ;
        RECT 7.545 1.125 8.575 1.295 ;
        RECT 9.620 0.605 9.790 0.945 ;
        RECT 8.405 0.605 9.790 0.775 ;
        RECT 9.620 0.775 11.200 0.945 ;
        RECT 11.030 0.775 11.200 1.760 ;
        RECT 9.850 1.125 10.020 1.560 ;
        RECT 9.850 1.125 10.850 1.295 ;
        RECT 10.680 1.125 10.850 2.215 ;
        RECT 10.680 2.045 11.255 2.215 ;
        RECT 9.045 0.955 9.405 1.125 ;
        RECT 9.235 0.955 9.405 2.215 ;
        RECT 9.150 2.045 10.500 2.215 ;
        RECT 10.330 1.610 10.500 2.630 ;
        RECT 11.610 1.540 11.780 2.630 ;
        RECT 10.330 2.460 11.780 2.630 ;
  END 
END FFSDQRHDLXHT

MACRO FFSDQRHD2XHT
  CLASS  CORE ;
  FOREIGN FFSDQRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.120 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 12.260 0.720 12.430 2.960 ;
        RECT 12.260 1.645 12.610 2.015 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 8.105 1.540 8.585 2.130 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.355 -0.300 2.655 0.595 ;
        RECT 3.415 -0.300 3.715 0.595 ;
        RECT 6.070 -0.300 6.370 1.055 ;
        RECT 7.140 -0.300 7.440 0.595 ;
        RECT 8.310 -0.300 8.480 0.780 ;
        RECT 10.145 -0.300 10.445 0.595 ;
        RECT 11.630 -0.300 11.930 1.055 ;
        RECT 12.715 -0.300 13.015 1.055 ;
        RECT 0.000 -0.300 13.120 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.880 1.525 3.395 1.950 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.355 2.345 2.655 3.990 ;
        RECT 3.290 2.620 3.460 3.990 ;
        RECT 6.085 3.140 6.385 3.990 ;
        RECT 8.245 3.095 8.545 3.990 ;
        RECT 10.245 2.810 10.545 3.990 ;
        RECT 11.675 2.975 11.975 3.990 ;
        RECT 12.715 2.295 13.015 3.990 ;
        RECT 0.000 3.390 13.120 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.555 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.150 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.980 0.775 2.150 1.035 ;
        RECT 1.530 0.865 2.150 1.035 ;
        RECT 1.980 0.775 4.675 0.945 ;
        RECT 4.505 0.775 4.675 2.280 ;
        RECT 5.205 0.910 5.375 2.280 ;
        RECT 6.280 1.675 6.580 1.865 ;
        RECT 5.205 1.695 6.580 1.865 ;
        RECT 5.800 1.325 6.100 1.515 ;
        RECT 5.800 1.325 6.930 1.495 ;
        RECT 6.655 0.775 6.825 1.495 ;
        RECT 6.760 1.325 6.930 2.215 ;
        RECT 6.760 2.045 7.410 2.215 ;
        RECT 7.620 0.480 7.790 0.945 ;
        RECT 6.655 0.775 7.790 0.945 ;
        RECT 2.865 1.125 3.750 1.295 ;
        RECT 2.865 2.130 3.810 2.300 ;
        RECT 3.580 1.125 3.750 2.300 ;
        RECT 3.640 1.525 3.810 3.035 ;
        RECT 3.580 1.525 3.875 1.825 ;
        RECT 5.750 2.815 5.820 3.035 ;
        RECT 5.740 2.825 9.115 2.915 ;
        RECT 5.760 2.805 5.820 3.035 ;
        RECT 5.730 2.835 9.115 2.915 ;
        RECT 5.770 2.795 5.820 3.035 ;
        RECT 5.720 2.845 9.115 2.915 ;
        RECT 3.640 2.865 5.820 3.035 ;
        RECT 3.640 2.865 5.830 3.024 ;
        RECT 3.640 2.865 5.840 3.014 ;
        RECT 3.640 2.865 5.850 3.004 ;
        RECT 3.640 2.865 5.860 2.994 ;
        RECT 3.640 2.865 5.870 2.984 ;
        RECT 3.640 2.865 5.880 2.974 ;
        RECT 3.640 2.865 5.890 2.964 ;
        RECT 5.775 2.790 8.075 2.960 ;
        RECT 5.710 2.855 9.115 2.915 ;
        RECT 7.905 2.745 8.075 2.960 ;
        RECT 7.905 2.745 9.115 2.915 ;
        RECT 8.945 2.745 9.115 3.210 ;
        RECT 8.945 3.040 9.775 3.210 ;
        RECT 3.930 1.125 4.250 1.295 ;
        RECT 4.080 1.125 4.250 2.685 ;
        RECT 3.995 1.980 4.250 2.685 ;
        RECT 4.855 0.535 5.025 2.685 ;
        RECT 5.490 2.465 5.560 2.685 ;
        RECT 5.480 2.475 9.800 2.565 ;
        RECT 5.500 2.455 5.560 2.685 ;
        RECT 5.470 2.485 9.800 2.565 ;
        RECT 5.510 2.445 5.560 2.685 ;
        RECT 5.460 2.495 9.800 2.565 ;
        RECT 3.995 2.515 5.560 2.685 ;
        RECT 3.995 2.515 5.570 2.674 ;
        RECT 3.995 2.515 5.580 2.664 ;
        RECT 3.995 2.515 5.590 2.654 ;
        RECT 3.995 2.515 5.600 2.644 ;
        RECT 3.995 2.515 5.610 2.634 ;
        RECT 4.855 0.535 5.620 0.705 ;
        RECT 3.995 2.515 5.620 2.624 ;
        RECT 3.995 2.515 5.630 2.614 ;
        RECT 5.515 2.440 7.720 2.610 ;
        RECT 5.450 2.505 9.800 2.565 ;
        RECT 7.550 2.395 7.720 2.610 ;
        RECT 8.905 1.355 9.075 2.565 ;
        RECT 8.905 1.355 9.205 1.525 ;
        RECT 7.550 2.395 9.800 2.565 ;
        RECT 9.630 2.395 9.800 2.795 ;
        RECT 7.110 1.575 7.925 1.745 ;
        RECT 7.755 1.125 7.925 2.215 ;
        RECT 7.625 2.045 7.925 2.215 ;
        RECT 8.295 0.960 8.465 1.295 ;
        RECT 7.695 1.125 8.465 1.295 ;
        RECT 8.295 0.960 8.830 1.130 ;
        RECT 8.660 0.635 8.830 1.130 ;
        RECT 9.780 0.635 9.950 0.945 ;
        RECT 8.660 0.635 9.950 0.805 ;
        RECT 9.780 0.775 11.415 0.945 ;
        RECT 11.245 0.775 11.415 1.670 ;
        RECT 10.725 1.125 11.065 1.495 ;
        RECT 9.935 1.325 11.065 1.495 ;
        RECT 10.895 1.125 11.065 2.215 ;
        RECT 10.895 2.045 11.465 2.215 ;
        RECT 9.195 0.985 9.600 1.155 ;
        RECT 9.430 0.985 9.600 2.215 ;
        RECT 9.300 2.045 9.600 2.215 ;
        RECT 9.430 1.675 10.715 1.845 ;
        RECT 10.545 1.675 10.715 2.630 ;
        RECT 11.910 1.610 12.080 2.630 ;
        RECT 10.545 2.460 12.080 2.630 ;
  END 
END FFSDQRHD2XHT

MACRO FFSDQRHD1XHT
  CLASS  CORE ;
  FOREIGN FFSDQRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.300 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.960 0.720 12.200 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.960 1.610 8.510 2.010 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.385 -0.300 2.685 0.595 ;
        RECT 3.335 -0.300 3.635 0.595 ;
        RECT 5.945 -0.300 6.245 1.145 ;
        RECT 6.985 -0.300 7.285 0.595 ;
        RECT 8.055 -0.300 8.225 0.810 ;
        RECT 9.995 -0.300 10.295 0.525 ;
        RECT 11.440 -0.300 11.610 1.120 ;
        RECT 0.000 -0.300 12.300 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.740 1.525 3.230 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.565 2.740 3.235 3.990 ;
        RECT 5.965 3.195 6.265 3.990 ;
        RECT 8.095 3.195 8.395 3.990 ;
        RECT 10.035 2.810 10.335 3.990 ;
        RECT 11.375 2.975 11.675 3.990 ;
        RECT 0.000 3.390 12.300 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.575 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.150 ;
        RECT 1.530 0.885 1.700 2.280 ;
        RECT 1.970 0.775 2.140 1.055 ;
        RECT 1.530 0.885 2.140 1.055 ;
        RECT 1.970 0.775 4.510 0.945 ;
        RECT 4.340 0.775 4.510 2.280 ;
        RECT 5.040 0.900 5.210 2.280 ;
        RECT 6.165 1.675 6.465 1.865 ;
        RECT 5.040 1.695 6.465 1.865 ;
        RECT 5.685 1.325 5.985 1.515 ;
        RECT 6.580 0.775 6.815 1.495 ;
        RECT 5.685 1.325 6.815 1.495 ;
        RECT 6.645 0.775 6.815 2.215 ;
        RECT 6.645 2.045 7.185 2.215 ;
        RECT 7.470 0.480 7.640 0.945 ;
        RECT 6.580 0.775 7.640 0.945 ;
        RECT 2.785 1.125 3.585 1.295 ;
        RECT 2.785 2.190 3.645 2.360 ;
        RECT 3.415 1.125 3.585 2.360 ;
        RECT 3.475 1.525 3.645 3.015 ;
        RECT 3.415 1.525 3.710 1.825 ;
        RECT 8.545 2.745 8.715 3.015 ;
        RECT 3.475 2.845 8.715 3.015 ;
        RECT 8.545 2.745 9.135 2.915 ;
        RECT 3.830 1.980 4.085 2.280 ;
        RECT 3.765 1.125 4.085 1.295 ;
        RECT 3.890 1.125 4.085 2.665 ;
        RECT 3.850 1.980 4.085 2.665 ;
        RECT 4.690 0.535 4.860 2.665 ;
        RECT 4.690 0.535 5.485 0.705 ;
        RECT 8.035 2.395 8.205 2.665 ;
        RECT 3.850 2.495 8.205 2.665 ;
        RECT 8.775 1.330 8.945 2.565 ;
        RECT 8.755 1.330 9.055 1.500 ;
        RECT 8.035 2.395 9.650 2.565 ;
        RECT 9.480 2.395 9.650 2.795 ;
        RECT 6.995 1.600 7.740 1.770 ;
        RECT 7.570 1.125 7.740 2.280 ;
        RECT 8.405 0.605 8.575 1.295 ;
        RECT 7.545 1.125 8.575 1.295 ;
        RECT 9.620 0.605 9.790 0.945 ;
        RECT 8.405 0.605 9.790 0.775 ;
        RECT 9.620 0.775 11.200 0.945 ;
        RECT 11.030 0.775 11.200 1.715 ;
        RECT 9.850 1.125 10.020 1.560 ;
        RECT 9.850 1.125 10.850 1.295 ;
        RECT 10.680 1.125 10.850 2.215 ;
        RECT 10.680 2.045 11.255 2.215 ;
        RECT 9.045 0.955 9.405 1.125 ;
        RECT 9.235 0.955 9.405 2.215 ;
        RECT 9.150 2.045 10.500 2.215 ;
        RECT 10.330 1.610 10.500 2.630 ;
        RECT 11.610 1.540 11.780 2.630 ;
        RECT 10.330 2.460 11.780 2.630 ;
  END 
END FFSDQRHD1XHT

MACRO FFSDQHDMXHT
  CLASS  CORE ;
  FOREIGN FFSDQHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.320 1.060 10.560 1.360 ;
        RECT 10.350 1.060 10.560 2.440 ;
        RECT 10.320 1.980 10.560 2.440 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.415 -0.300 2.715 0.595 ;
        RECT 3.325 -0.300 3.625 0.595 ;
        RECT 5.815 -0.300 6.115 0.595 ;
        RECT 6.755 -0.300 7.055 0.595 ;
        RECT 8.655 -0.300 8.955 1.110 ;
        RECT 9.735 -0.300 10.035 1.145 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.740 1.525 3.230 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.630 2.740 3.270 3.990 ;
        RECT 6.000 3.160 6.980 3.990 ;
        RECT 8.710 2.745 8.880 3.990 ;
        RECT 9.705 2.775 10.005 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.555 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.150 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.975 0.775 2.145 1.035 ;
        RECT 1.530 0.865 2.145 1.035 ;
        RECT 1.975 0.775 4.510 0.945 ;
        RECT 4.275 0.550 4.510 0.945 ;
        RECT 4.340 0.550 4.510 2.280 ;
        RECT 4.340 1.960 4.520 2.280 ;
        RECT 4.340 1.970 4.530 2.280 ;
        RECT 4.340 1.980 4.540 2.280 ;
        RECT 5.070 0.910 5.210 2.280 ;
        RECT 6.185 1.675 6.485 1.865 ;
        RECT 5.390 1.695 6.485 1.865 ;
        RECT 5.240 1.555 5.250 1.865 ;
        RECT 5.250 1.565 5.260 1.865 ;
        RECT 5.260 1.575 5.270 1.865 ;
        RECT 5.270 1.585 5.280 1.865 ;
        RECT 5.280 1.595 5.290 1.865 ;
        RECT 5.290 1.605 5.300 1.865 ;
        RECT 5.300 1.615 5.310 1.865 ;
        RECT 5.310 1.625 5.320 1.865 ;
        RECT 5.320 1.635 5.330 1.865 ;
        RECT 5.330 1.645 5.340 1.865 ;
        RECT 5.340 1.655 5.350 1.865 ;
        RECT 5.350 1.665 5.360 1.865 ;
        RECT 5.360 1.675 5.370 1.865 ;
        RECT 5.370 1.685 5.380 1.865 ;
        RECT 5.380 1.695 5.390 1.865 ;
        RECT 5.210 1.525 5.220 2.279 ;
        RECT 5.220 1.535 5.230 2.279 ;
        RECT 5.230 1.545 5.240 2.279 ;
        RECT 5.040 0.910 5.050 1.590 ;
        RECT 5.050 0.910 5.060 1.600 ;
        RECT 5.060 0.910 5.070 1.610 ;
        RECT 5.685 1.325 5.985 1.515 ;
        RECT 6.430 0.910 6.600 1.495 ;
        RECT 5.685 1.325 7.165 1.495 ;
        RECT 6.995 1.325 7.165 2.215 ;
        RECT 6.365 2.045 7.165 2.215 ;
        RECT 2.805 1.125 3.665 1.295 ;
        RECT 2.785 2.190 3.680 2.360 ;
        RECT 3.475 1.125 3.665 2.980 ;
        RECT 3.415 1.125 3.665 2.360 ;
        RECT 3.475 1.525 3.680 2.980 ;
        RECT 3.415 1.525 3.735 1.825 ;
        RECT 3.475 2.810 7.635 2.980 ;
        RECT 3.860 1.980 4.085 2.280 ;
        RECT 3.915 1.125 4.085 2.630 ;
        RECT 3.845 1.125 4.145 1.295 ;
        RECT 4.700 1.790 4.890 1.869 ;
        RECT 4.710 1.790 4.890 1.879 ;
        RECT 4.690 0.535 4.860 1.859 ;
        RECT 4.690 1.770 4.870 1.859 ;
        RECT 4.690 1.780 4.880 1.859 ;
        RECT 4.720 1.790 4.890 2.630 ;
        RECT 4.690 0.535 5.485 0.705 ;
        RECT 7.345 0.500 7.515 2.630 ;
        RECT 7.345 0.500 7.745 0.670 ;
        RECT 7.345 2.440 8.150 2.630 ;
        RECT 3.915 2.460 8.150 2.630 ;
        RECT 7.980 2.440 8.150 2.770 ;
        RECT 8.405 1.460 9.495 1.630 ;
        RECT 9.290 0.875 9.460 1.630 ;
        RECT 9.325 1.460 9.495 2.215 ;
        RECT 9.195 2.045 9.495 2.215 ;
        RECT 7.770 0.875 7.940 2.215 ;
        RECT 7.695 2.045 8.905 2.215 ;
        RECT 8.735 2.045 8.905 2.565 ;
        RECT 9.080 2.395 9.250 2.780 ;
        RECT 9.970 1.520 10.140 2.565 ;
        RECT 8.735 2.395 10.140 2.565 ;
        RECT 9.970 1.520 10.160 1.820 ;
  END 
END FFSDQHDMXHT

MACRO FFSDQHDLXHT
  CLASS  CORE ;
  FOREIGN FFSDQHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.320 1.060 10.560 2.445 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.350 2.980 ;
        RECT 1.180 2.810 1.350 3.110 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.375 -0.300 2.675 0.595 ;
        RECT 3.405 -0.300 3.705 0.595 ;
        RECT 5.875 -0.300 6.175 0.595 ;
        RECT 6.835 -0.300 7.135 0.565 ;
        RECT 8.715 -0.300 9.015 0.560 ;
        RECT 9.705 -0.300 10.005 1.295 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.790 1.525 3.280 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.265 2.735 2.565 3.990 ;
        RECT 3.175 2.675 3.345 3.990 ;
        RECT 6.060 3.160 7.040 3.990 ;
        RECT 8.710 2.745 8.880 3.990 ;
        RECT 9.705 2.745 10.005 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.555 0.650 ;
        RECT 1.180 2.460 1.880 2.630 ;
        RECT 1.710 2.460 1.880 2.835 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.530 0.865 1.720 1.185 ;
        RECT 2.000 0.775 2.170 1.035 ;
        RECT 1.530 0.865 2.170 1.035 ;
        RECT 2.000 0.775 4.570 0.945 ;
        RECT 4.335 0.485 4.570 0.945 ;
        RECT 4.400 0.485 4.570 2.280 ;
        RECT 5.100 0.900 5.270 2.280 ;
        RECT 6.235 1.675 6.535 1.865 ;
        RECT 5.100 1.695 6.535 1.865 ;
        RECT 5.745 1.325 6.045 1.515 ;
        RECT 6.510 0.900 6.680 1.495 ;
        RECT 5.745 1.325 7.225 1.495 ;
        RECT 7.055 1.325 7.225 2.215 ;
        RECT 6.425 2.045 7.225 2.215 ;
        RECT 2.825 1.125 3.635 1.295 ;
        RECT 2.805 2.190 3.695 2.360 ;
        RECT 3.465 1.125 3.635 2.360 ;
        RECT 3.525 1.525 3.695 3.020 ;
        RECT 3.465 1.525 3.760 1.825 ;
        RECT 5.245 2.810 5.545 3.020 ;
        RECT 3.525 2.850 5.545 3.020 ;
        RECT 5.245 2.810 7.695 2.980 ;
        RECT 3.955 1.125 4.135 2.670 ;
        RECT 3.910 2.370 4.135 2.670 ;
        RECT 3.865 1.125 4.165 1.295 ;
        RECT 4.750 0.535 4.920 2.630 ;
        RECT 4.750 0.535 5.545 0.705 ;
        RECT 7.425 0.500 7.595 2.630 ;
        RECT 7.425 0.500 7.875 0.670 ;
        RECT 7.425 2.440 8.230 2.630 ;
        RECT 3.910 2.460 8.230 2.630 ;
        RECT 8.060 2.440 8.230 2.740 ;
        RECT 8.475 1.435 9.495 1.605 ;
        RECT 9.260 0.875 9.430 1.605 ;
        RECT 9.325 1.435 9.495 2.215 ;
        RECT 9.195 2.045 9.495 2.215 ;
        RECT 7.850 0.875 8.020 2.215 ;
        RECT 7.775 2.045 8.965 2.215 ;
        RECT 8.795 2.045 8.965 2.565 ;
        RECT 9.080 2.395 9.250 2.695 ;
        RECT 9.970 1.540 10.140 2.565 ;
        RECT 8.795 2.395 10.140 2.565 ;
  END 
END FFSDQHDLXHT

MACRO FFSDQHD2XHT
  CLASS  CORE ;
  FOREIGN FFSDQHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.480 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.620 0.720 10.790 2.960 ;
        RECT 10.620 1.645 10.970 2.015 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.595 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.385 -0.300 2.685 0.595 ;
        RECT 3.490 -0.300 3.790 0.595 ;
        RECT 6.085 -0.300 6.385 0.595 ;
        RECT 7.145 -0.300 7.445 1.055 ;
        RECT 8.890 -0.300 9.060 0.780 ;
        RECT 10.035 -0.300 10.335 1.055 ;
        RECT 11.075 -0.300 11.375 1.055 ;
        RECT 0.000 -0.300 11.480 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.970 1.525 3.505 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.385 2.345 2.685 3.990 ;
        RECT 3.400 2.675 3.570 3.990 ;
        RECT 6.195 3.160 6.495 3.990 ;
        RECT 7.115 3.095 7.415 3.990 ;
        RECT 9.010 2.810 9.180 3.990 ;
        RECT 10.035 2.975 10.335 3.990 ;
        RECT 11.075 2.295 11.375 3.990 ;
        RECT 0.000 3.390 11.480 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.555 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.150 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.970 0.775 2.140 1.035 ;
        RECT 1.530 0.865 2.140 1.035 ;
        RECT 1.970 0.775 4.785 0.945 ;
        RECT 4.615 0.775 4.785 2.280 ;
        RECT 5.315 0.910 5.485 2.280 ;
        RECT 6.455 1.675 6.755 1.865 ;
        RECT 5.315 1.695 6.755 1.865 ;
        RECT 5.910 1.325 6.210 1.515 ;
        RECT 6.700 0.910 6.870 1.495 ;
        RECT 5.910 1.325 7.535 1.495 ;
        RECT 7.365 1.325 7.535 2.215 ;
        RECT 6.635 2.045 7.535 2.215 ;
        RECT 2.920 1.125 3.860 1.295 ;
        RECT 2.920 2.190 3.920 2.360 ;
        RECT 3.690 1.125 3.860 2.360 ;
        RECT 3.750 1.525 3.920 3.035 ;
        RECT 3.690 1.525 3.985 1.825 ;
        RECT 3.750 2.865 5.810 3.035 ;
        RECT 6.050 2.745 7.765 2.915 ;
        RECT 7.595 2.745 7.765 3.145 ;
        RECT 7.595 2.975 8.615 3.145 ;
        RECT 8.315 2.975 8.615 3.210 ;
        RECT 5.930 2.745 5.940 3.025 ;
        RECT 5.940 2.745 5.950 3.015 ;
        RECT 5.950 2.745 5.960 3.005 ;
        RECT 5.960 2.745 5.970 2.995 ;
        RECT 5.970 2.745 5.980 2.985 ;
        RECT 5.980 2.745 5.990 2.975 ;
        RECT 5.990 2.745 6.000 2.965 ;
        RECT 6.000 2.745 6.010 2.955 ;
        RECT 6.010 2.745 6.020 2.945 ;
        RECT 6.020 2.745 6.030 2.935 ;
        RECT 6.030 2.745 6.040 2.925 ;
        RECT 6.040 2.745 6.050 2.915 ;
        RECT 5.810 2.865 5.820 3.035 ;
        RECT 5.820 2.855 5.830 3.035 ;
        RECT 5.830 2.845 5.840 3.035 ;
        RECT 5.840 2.835 5.850 3.035 ;
        RECT 5.850 2.825 5.860 3.035 ;
        RECT 5.860 2.815 5.870 3.035 ;
        RECT 5.870 2.805 5.880 3.035 ;
        RECT 5.880 2.795 5.890 3.035 ;
        RECT 5.890 2.785 5.900 3.035 ;
        RECT 5.900 2.775 5.910 3.035 ;
        RECT 5.910 2.765 5.920 3.035 ;
        RECT 5.920 2.755 5.930 3.035 ;
        RECT 8.805 1.610 9.760 1.780 ;
        RECT 9.590 1.060 9.760 2.280 ;
        RECT 4.040 1.125 4.360 1.295 ;
        RECT 4.165 1.125 4.360 2.685 ;
        RECT 4.105 1.980 4.360 2.685 ;
        RECT 4.965 0.535 5.135 2.685 ;
        RECT 4.105 2.515 5.590 2.685 ;
        RECT 4.965 0.535 5.730 0.705 ;
        RECT 7.715 0.710 7.850 2.565 ;
        RECT 5.790 2.395 7.850 2.565 ;
        RECT 7.995 2.455 8.550 2.625 ;
        RECT 7.885 0.710 8.655 0.880 ;
        RECT 8.380 2.455 8.550 2.795 ;
        RECT 8.485 0.710 8.655 1.140 ;
        RECT 9.240 0.480 9.410 1.140 ;
        RECT 8.485 0.970 9.410 1.140 ;
        RECT 9.240 0.480 9.820 0.650 ;
        RECT 7.910 2.380 7.920 2.624 ;
        RECT 7.920 2.390 7.930 2.624 ;
        RECT 7.930 2.400 7.940 2.624 ;
        RECT 7.940 2.410 7.950 2.624 ;
        RECT 7.950 2.420 7.960 2.624 ;
        RECT 7.960 2.430 7.970 2.624 ;
        RECT 7.970 2.440 7.980 2.624 ;
        RECT 7.980 2.450 7.990 2.624 ;
        RECT 7.990 2.455 7.996 2.625 ;
        RECT 7.885 2.355 7.895 2.599 ;
        RECT 7.895 2.365 7.905 2.609 ;
        RECT 7.905 2.370 7.911 2.620 ;
        RECT 7.850 0.710 7.860 2.564 ;
        RECT 7.860 0.710 7.870 2.574 ;
        RECT 7.870 0.710 7.880 2.584 ;
        RECT 7.880 0.710 7.886 2.594 ;
        RECT 5.710 2.395 5.720 2.635 ;
        RECT 5.720 2.395 5.730 2.625 ;
        RECT 5.730 2.395 5.740 2.615 ;
        RECT 5.740 2.395 5.750 2.605 ;
        RECT 5.750 2.395 5.760 2.595 ;
        RECT 5.760 2.395 5.770 2.585 ;
        RECT 5.770 2.395 5.780 2.575 ;
        RECT 5.780 2.395 5.790 2.565 ;
        RECT 5.670 2.435 5.680 2.675 ;
        RECT 5.680 2.425 5.690 2.665 ;
        RECT 5.690 2.415 5.700 2.655 ;
        RECT 5.700 2.405 5.710 2.645 ;
        RECT 5.590 2.515 5.600 2.685 ;
        RECT 5.600 2.505 5.610 2.685 ;
        RECT 5.610 2.495 5.620 2.685 ;
        RECT 5.620 2.485 5.630 2.685 ;
        RECT 5.630 2.475 5.640 2.685 ;
        RECT 5.640 2.465 5.650 2.685 ;
        RECT 5.650 2.455 5.660 2.685 ;
        RECT 5.660 2.445 5.670 2.685 ;
        RECT 8.130 1.060 8.300 2.230 ;
        RECT 8.065 2.060 9.410 2.230 ;
        RECT 9.240 2.060 9.410 2.630 ;
        RECT 9.380 2.460 9.550 2.770 ;
        RECT 10.270 1.610 10.440 2.630 ;
        RECT 9.240 2.460 10.440 2.630 ;
  END 
END FFSDQHD2XHT

MACRO FFSDQHD1XHT
  CLASS  CORE ;
  FOREIGN FFSDQHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.320 0.720 10.560 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.595 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.385 -0.300 2.685 0.595 ;
        RECT 3.335 -0.300 3.635 0.595 ;
        RECT 5.815 -0.300 6.115 0.595 ;
        RECT 6.755 -0.300 7.055 0.565 ;
        RECT 8.645 -0.300 8.945 0.630 ;
        RECT 9.735 -0.300 10.035 1.055 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.740 1.525 3.230 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.625 2.740 3.265 3.990 ;
        RECT 5.995 3.160 6.975 3.990 ;
        RECT 8.660 2.745 8.830 3.990 ;
        RECT 9.735 2.975 10.035 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.555 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.150 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.980 0.775 2.150 1.035 ;
        RECT 1.530 0.865 2.150 1.035 ;
        RECT 1.980 0.775 4.510 0.945 ;
        RECT 4.340 0.775 4.510 2.280 ;
        RECT 5.040 0.900 5.210 2.280 ;
        RECT 6.185 1.675 6.495 1.865 ;
        RECT 5.040 1.695 6.495 1.865 ;
        RECT 5.685 1.325 5.985 1.515 ;
        RECT 6.430 0.910 6.600 1.495 ;
        RECT 5.685 1.325 7.165 1.495 ;
        RECT 6.995 1.325 7.165 2.215 ;
        RECT 6.365 2.045 7.165 2.215 ;
        RECT 2.785 1.125 3.585 1.295 ;
        RECT 2.785 2.190 3.645 2.360 ;
        RECT 3.415 1.125 3.585 2.360 ;
        RECT 3.475 1.525 3.645 2.980 ;
        RECT 3.415 1.525 3.710 1.825 ;
        RECT 3.475 2.810 7.745 2.980 ;
        RECT 3.830 1.980 4.085 2.280 ;
        RECT 3.765 1.125 4.085 1.295 ;
        RECT 3.890 1.125 4.085 2.630 ;
        RECT 3.850 1.980 4.085 2.630 ;
        RECT 4.690 0.535 4.860 2.630 ;
        RECT 4.690 0.535 5.485 0.705 ;
        RECT 7.345 0.500 7.515 2.630 ;
        RECT 7.345 0.500 7.745 0.670 ;
        RECT 7.345 2.440 8.190 2.630 ;
        RECT 3.850 2.460 8.190 2.630 ;
        RECT 8.020 2.440 8.190 2.770 ;
        RECT 8.405 1.380 9.445 1.550 ;
        RECT 9.240 0.945 9.410 1.550 ;
        RECT 9.275 1.380 9.445 2.215 ;
        RECT 9.145 2.045 9.445 2.215 ;
        RECT 7.760 0.945 7.930 2.215 ;
        RECT 7.695 2.045 8.905 2.215 ;
        RECT 8.735 2.045 8.905 2.565 ;
        RECT 9.030 2.395 9.200 2.780 ;
        RECT 9.970 1.520 10.140 2.565 ;
        RECT 8.735 2.395 10.140 2.565 ;
  END 
END FFSDQHD1XHT

MACRO FFSDNSRHDMXHT
  CLASS  CORE ;
  FOREIGN FFSDNSRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.760 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.965 1.550 3.305 2.015 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.405 0.830 14.575 2.280 ;
        RECT 14.405 0.830 14.660 1.230 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.220 0.820 13.705 1.295 ;
        RECT 13.535 0.820 13.705 2.215 ;
        RECT 13.300 2.045 13.705 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.325 0.855 1.545 1.460 ;
        RECT 0.855 1.290 1.545 1.460 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.840 1.540 6.385 2.110 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.455 1.640 0.625 1.945 ;
        RECT 0.815 1.775 1.290 2.365 ;
        RECT 1.370 1.640 1.540 1.945 ;
        RECT 0.455 1.775 1.540 1.945 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.060 ;
        RECT 2.610 -0.300 3.595 0.785 ;
        RECT 5.970 -0.300 6.270 1.130 ;
        RECT 8.765 -0.300 8.935 1.345 ;
        RECT 10.745 -0.300 11.045 0.860 ;
        RECT 12.715 -0.300 13.015 0.720 ;
        RECT 13.885 -0.300 14.055 1.210 ;
        RECT 0.000 -0.300 14.760 0.300 ;
    END
  END GND
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.290 1.610 2.775 2.015 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 12.315 1.540 12.760 1.950 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.545 2.975 0.845 3.990 ;
        RECT 2.475 2.995 3.455 3.990 ;
        RECT 6.170 2.995 7.150 3.990 ;
        RECT 8.700 2.995 9.000 3.990 ;
        RECT 10.800 2.365 11.100 3.990 ;
        RECT 12.665 2.830 12.965 3.990 ;
        RECT 13.790 2.925 14.090 3.990 ;
        RECT 0.000 3.390 14.760 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.130 0.340 2.430 ;
        RECT 0.105 0.890 0.275 2.430 ;
        RECT 0.170 2.130 0.340 2.795 ;
        RECT 0.105 0.890 0.405 1.060 ;
        RECT 0.170 2.625 1.305 2.795 ;
        RECT 1.135 2.625 1.305 3.115 ;
        RECT 1.135 2.945 1.995 3.115 ;
        RECT 2.805 1.125 3.750 1.295 ;
        RECT 3.580 1.125 3.750 2.365 ;
        RECT 2.825 2.195 3.750 2.365 ;
        RECT 1.725 0.825 1.985 1.125 ;
        RECT 1.815 0.825 1.985 2.715 ;
        RECT 1.580 2.150 1.985 2.715 ;
        RECT 4.445 1.045 4.615 2.715 ;
        RECT 1.580 2.545 4.615 2.715 ;
        RECT 3.930 0.695 4.100 2.310 ;
        RECT 3.930 0.695 5.545 0.865 ;
        RECT 5.375 0.695 5.545 2.245 ;
        RECT 6.555 0.895 6.755 1.195 ;
        RECT 6.585 0.895 6.755 2.115 ;
        RECT 6.585 1.445 7.345 1.745 ;
        RECT 5.025 1.045 5.195 2.595 ;
        RECT 5.025 2.425 5.705 2.595 ;
        RECT 7.525 1.680 7.695 2.465 ;
        RECT 5.910 2.295 7.695 2.465 ;
        RECT 7.775 1.550 7.945 1.850 ;
        RECT 7.525 1.680 7.945 1.850 ;
        RECT 5.835 2.295 5.845 2.529 ;
        RECT 5.845 2.295 5.855 2.519 ;
        RECT 5.855 2.295 5.865 2.509 ;
        RECT 5.865 2.295 5.875 2.499 ;
        RECT 5.875 2.295 5.885 2.489 ;
        RECT 5.885 2.295 5.895 2.479 ;
        RECT 5.895 2.295 5.905 2.469 ;
        RECT 5.905 2.295 5.911 2.465 ;
        RECT 5.780 2.350 5.790 2.584 ;
        RECT 5.790 2.340 5.800 2.574 ;
        RECT 5.800 2.330 5.810 2.564 ;
        RECT 5.810 2.320 5.820 2.554 ;
        RECT 5.820 2.310 5.830 2.544 ;
        RECT 5.830 2.300 5.836 2.540 ;
        RECT 5.705 2.425 5.715 2.595 ;
        RECT 5.715 2.415 5.725 2.595 ;
        RECT 5.725 2.405 5.735 2.595 ;
        RECT 5.735 2.395 5.745 2.595 ;
        RECT 5.745 2.385 5.755 2.595 ;
        RECT 5.755 2.375 5.765 2.595 ;
        RECT 5.765 2.365 5.775 2.595 ;
        RECT 5.775 2.355 5.781 2.595 ;
        RECT 7.000 0.960 7.300 1.215 ;
        RECT 7.000 1.045 8.235 1.215 ;
        RECT 8.065 1.045 8.235 1.345 ;
        RECT 6.990 0.525 7.160 0.730 ;
        RECT 6.630 0.525 7.160 0.695 ;
        RECT 7.890 2.045 8.015 2.215 ;
        RECT 8.125 1.535 8.190 2.215 ;
        RECT 6.990 0.560 8.585 0.730 ;
        RECT 8.415 0.560 8.585 1.705 ;
        RECT 8.295 1.535 9.210 1.705 ;
        RECT 8.190 1.535 8.200 2.105 ;
        RECT 8.200 1.535 8.210 2.095 ;
        RECT 8.210 1.535 8.220 2.085 ;
        RECT 8.220 1.535 8.230 2.075 ;
        RECT 8.230 1.535 8.240 2.065 ;
        RECT 8.240 1.535 8.250 2.055 ;
        RECT 8.250 1.535 8.260 2.045 ;
        RECT 8.260 1.535 8.270 2.035 ;
        RECT 8.270 1.535 8.280 2.025 ;
        RECT 8.280 1.535 8.290 2.015 ;
        RECT 8.290 1.535 8.296 2.009 ;
        RECT 8.015 2.045 8.025 2.215 ;
        RECT 8.025 2.035 8.035 2.215 ;
        RECT 8.035 2.025 8.045 2.215 ;
        RECT 8.045 2.015 8.055 2.215 ;
        RECT 8.055 2.005 8.065 2.215 ;
        RECT 8.065 1.995 8.075 2.215 ;
        RECT 8.075 1.985 8.085 2.215 ;
        RECT 8.085 1.975 8.095 2.215 ;
        RECT 8.095 1.965 8.105 2.215 ;
        RECT 8.105 1.955 8.115 2.215 ;
        RECT 8.115 1.945 8.125 2.215 ;
        RECT 3.655 2.895 5.735 3.065 ;
        RECT 7.875 2.425 8.045 2.815 ;
        RECT 6.095 2.645 8.045 2.815 ;
        RECT 7.875 2.425 8.240 2.595 ;
        RECT 8.445 2.295 9.260 2.465 ;
        RECT 10.100 1.810 10.270 2.565 ;
        RECT 9.435 2.395 10.270 2.565 ;
        RECT 9.360 2.330 9.370 2.564 ;
        RECT 9.370 2.340 9.380 2.564 ;
        RECT 9.380 2.350 9.390 2.564 ;
        RECT 9.390 2.360 9.400 2.564 ;
        RECT 9.400 2.370 9.410 2.564 ;
        RECT 9.410 2.380 9.420 2.564 ;
        RECT 9.420 2.390 9.430 2.564 ;
        RECT 9.430 2.395 9.436 2.565 ;
        RECT 9.335 2.305 9.345 2.539 ;
        RECT 9.345 2.315 9.355 2.549 ;
        RECT 9.355 2.320 9.361 2.560 ;
        RECT 9.260 2.295 9.270 2.465 ;
        RECT 9.270 2.295 9.280 2.475 ;
        RECT 9.280 2.295 9.290 2.485 ;
        RECT 9.290 2.295 9.300 2.495 ;
        RECT 9.300 2.295 9.310 2.505 ;
        RECT 9.310 2.295 9.320 2.515 ;
        RECT 9.320 2.295 9.330 2.525 ;
        RECT 9.330 2.295 9.336 2.535 ;
        RECT 8.370 2.295 8.380 2.529 ;
        RECT 8.380 2.295 8.390 2.519 ;
        RECT 8.390 2.295 8.400 2.509 ;
        RECT 8.400 2.295 8.410 2.499 ;
        RECT 8.410 2.295 8.420 2.489 ;
        RECT 8.420 2.295 8.430 2.479 ;
        RECT 8.430 2.295 8.440 2.469 ;
        RECT 8.440 2.295 8.446 2.465 ;
        RECT 8.315 2.350 8.325 2.584 ;
        RECT 8.325 2.340 8.335 2.574 ;
        RECT 8.335 2.330 8.345 2.564 ;
        RECT 8.345 2.320 8.355 2.554 ;
        RECT 8.355 2.310 8.365 2.544 ;
        RECT 8.365 2.300 8.371 2.540 ;
        RECT 8.240 2.425 8.250 2.595 ;
        RECT 8.250 2.415 8.260 2.595 ;
        RECT 8.260 2.405 8.270 2.595 ;
        RECT 8.270 2.395 8.280 2.595 ;
        RECT 8.280 2.385 8.290 2.595 ;
        RECT 8.290 2.375 8.300 2.595 ;
        RECT 8.300 2.365 8.310 2.595 ;
        RECT 8.310 2.355 8.316 2.595 ;
        RECT 5.985 2.645 5.995 2.915 ;
        RECT 5.995 2.645 6.005 2.905 ;
        RECT 6.005 2.645 6.015 2.895 ;
        RECT 6.015 2.645 6.025 2.885 ;
        RECT 6.025 2.645 6.035 2.875 ;
        RECT 6.035 2.645 6.045 2.865 ;
        RECT 6.045 2.645 6.055 2.855 ;
        RECT 6.055 2.645 6.065 2.845 ;
        RECT 6.065 2.645 6.075 2.835 ;
        RECT 6.075 2.645 6.085 2.825 ;
        RECT 6.085 2.645 6.095 2.815 ;
        RECT 5.845 2.785 5.855 3.055 ;
        RECT 5.855 2.775 5.865 3.045 ;
        RECT 5.865 2.765 5.875 3.035 ;
        RECT 5.875 2.755 5.885 3.025 ;
        RECT 5.885 2.745 5.895 3.015 ;
        RECT 5.895 2.735 5.905 3.005 ;
        RECT 5.905 2.725 5.915 2.995 ;
        RECT 5.915 2.715 5.925 2.985 ;
        RECT 5.925 2.705 5.935 2.975 ;
        RECT 5.935 2.695 5.945 2.965 ;
        RECT 5.945 2.685 5.955 2.955 ;
        RECT 5.955 2.675 5.965 2.945 ;
        RECT 5.965 2.665 5.975 2.935 ;
        RECT 5.975 2.655 5.985 2.925 ;
        RECT 5.735 2.895 5.745 3.065 ;
        RECT 5.745 2.885 5.755 3.065 ;
        RECT 5.755 2.875 5.765 3.065 ;
        RECT 5.765 2.865 5.775 3.065 ;
        RECT 5.775 2.855 5.785 3.065 ;
        RECT 5.785 2.845 5.795 3.065 ;
        RECT 5.795 2.835 5.805 3.065 ;
        RECT 5.805 2.825 5.815 3.065 ;
        RECT 5.815 2.815 5.825 3.065 ;
        RECT 5.825 2.805 5.835 3.065 ;
        RECT 5.835 2.795 5.845 3.065 ;
        RECT 8.235 2.835 8.355 3.210 ;
        RECT 7.410 3.040 8.355 3.210 ;
        RECT 8.620 2.645 9.105 2.815 ;
        RECT 10.055 1.270 10.295 1.440 ;
        RECT 9.280 2.745 10.450 2.915 ;
        RECT 10.450 1.360 10.460 2.914 ;
        RECT 10.460 1.370 10.470 2.914 ;
        RECT 10.470 1.380 10.480 2.914 ;
        RECT 10.480 1.390 10.490 2.914 ;
        RECT 10.490 1.400 10.500 2.914 ;
        RECT 10.500 1.410 10.510 2.914 ;
        RECT 10.510 1.420 10.520 2.914 ;
        RECT 10.520 1.430 10.530 2.914 ;
        RECT 10.530 1.440 10.540 2.914 ;
        RECT 10.540 1.450 10.550 2.914 ;
        RECT 10.550 1.460 10.560 2.914 ;
        RECT 10.560 1.470 10.570 2.914 ;
        RECT 10.570 1.480 10.580 2.914 ;
        RECT 10.580 1.490 10.590 2.914 ;
        RECT 10.590 1.500 10.600 2.914 ;
        RECT 10.600 1.510 10.610 2.914 ;
        RECT 10.610 1.520 10.620 2.914 ;
        RECT 10.370 1.280 10.380 1.514 ;
        RECT 10.380 1.290 10.390 1.524 ;
        RECT 10.390 1.300 10.400 1.534 ;
        RECT 10.400 1.310 10.410 1.544 ;
        RECT 10.410 1.320 10.420 1.554 ;
        RECT 10.420 1.330 10.430 1.564 ;
        RECT 10.430 1.340 10.440 1.574 ;
        RECT 10.440 1.350 10.450 1.584 ;
        RECT 10.295 1.270 10.305 1.440 ;
        RECT 10.305 1.270 10.315 1.450 ;
        RECT 10.315 1.270 10.325 1.460 ;
        RECT 10.325 1.270 10.335 1.470 ;
        RECT 10.335 1.270 10.345 1.480 ;
        RECT 10.345 1.270 10.355 1.490 ;
        RECT 10.355 1.270 10.365 1.500 ;
        RECT 10.365 1.270 10.371 1.510 ;
        RECT 9.205 2.680 9.215 2.914 ;
        RECT 9.215 2.690 9.225 2.914 ;
        RECT 9.225 2.700 9.235 2.914 ;
        RECT 9.235 2.710 9.245 2.914 ;
        RECT 9.245 2.720 9.255 2.914 ;
        RECT 9.255 2.730 9.265 2.914 ;
        RECT 9.265 2.740 9.275 2.914 ;
        RECT 9.275 2.745 9.281 2.915 ;
        RECT 9.180 2.655 9.190 2.889 ;
        RECT 9.190 2.665 9.200 2.899 ;
        RECT 9.200 2.670 9.206 2.910 ;
        RECT 9.105 2.645 9.115 2.815 ;
        RECT 9.115 2.645 9.125 2.825 ;
        RECT 9.125 2.645 9.135 2.835 ;
        RECT 9.135 2.645 9.145 2.845 ;
        RECT 9.145 2.645 9.155 2.855 ;
        RECT 9.155 2.645 9.165 2.865 ;
        RECT 9.165 2.645 9.175 2.875 ;
        RECT 9.175 2.645 9.181 2.885 ;
        RECT 8.545 2.645 8.555 2.879 ;
        RECT 8.555 2.645 8.565 2.869 ;
        RECT 8.565 2.645 8.575 2.859 ;
        RECT 8.575 2.645 8.585 2.849 ;
        RECT 8.585 2.645 8.595 2.839 ;
        RECT 8.595 2.645 8.605 2.829 ;
        RECT 8.605 2.645 8.615 2.819 ;
        RECT 8.615 2.645 8.621 2.815 ;
        RECT 8.405 2.785 8.415 3.019 ;
        RECT 8.415 2.775 8.425 3.009 ;
        RECT 8.425 2.765 8.435 2.999 ;
        RECT 8.435 2.755 8.445 2.989 ;
        RECT 8.445 2.745 8.455 2.979 ;
        RECT 8.455 2.735 8.465 2.969 ;
        RECT 8.465 2.725 8.475 2.959 ;
        RECT 8.475 2.715 8.485 2.949 ;
        RECT 8.485 2.705 8.495 2.939 ;
        RECT 8.495 2.695 8.505 2.929 ;
        RECT 8.505 2.685 8.515 2.919 ;
        RECT 8.515 2.675 8.525 2.909 ;
        RECT 8.525 2.665 8.535 2.899 ;
        RECT 8.535 2.655 8.545 2.889 ;
        RECT 8.355 2.835 8.365 3.209 ;
        RECT 8.365 2.825 8.375 3.209 ;
        RECT 8.375 2.815 8.385 3.209 ;
        RECT 8.385 2.805 8.395 3.209 ;
        RECT 8.395 2.795 8.405 3.209 ;
        RECT 11.355 0.760 11.525 1.280 ;
        RECT 11.225 1.110 11.525 1.280 ;
        RECT 11.355 0.760 12.435 0.930 ;
        RECT 12.265 0.760 12.435 1.280 ;
        RECT 12.265 1.110 12.565 1.280 ;
        RECT 11.150 1.460 11.320 1.760 ;
        RECT 11.745 1.110 12.045 1.630 ;
        RECT 11.150 1.460 12.045 1.630 ;
        RECT 11.875 1.110 12.045 2.300 ;
        RECT 12.940 1.540 13.110 2.300 ;
        RECT 11.875 2.130 13.110 2.300 ;
        RECT 12.940 1.540 13.355 1.840 ;
        RECT 9.620 0.900 9.790 2.215 ;
        RECT 9.620 2.045 9.920 2.215 ;
        RECT 9.620 0.900 10.430 1.070 ;
        RECT 10.645 1.040 10.970 1.210 ;
        RECT 10.800 1.040 10.970 2.110 ;
        RECT 10.800 1.940 11.530 2.110 ;
        RECT 11.360 1.940 11.530 2.650 ;
        RECT 11.935 2.480 12.235 2.855 ;
        RECT 14.055 1.515 14.225 2.650 ;
        RECT 11.360 2.480 14.225 2.650 ;
        RECT 10.570 0.975 10.580 1.209 ;
        RECT 10.580 0.985 10.590 1.209 ;
        RECT 10.590 0.995 10.600 1.209 ;
        RECT 10.600 1.005 10.610 1.209 ;
        RECT 10.610 1.015 10.620 1.209 ;
        RECT 10.620 1.025 10.630 1.209 ;
        RECT 10.630 1.035 10.640 1.209 ;
        RECT 10.640 1.040 10.646 1.210 ;
        RECT 10.505 0.910 10.515 1.144 ;
        RECT 10.515 0.920 10.525 1.154 ;
        RECT 10.525 0.930 10.535 1.164 ;
        RECT 10.535 0.940 10.545 1.174 ;
        RECT 10.545 0.950 10.555 1.184 ;
        RECT 10.555 0.960 10.565 1.194 ;
        RECT 10.565 0.965 10.571 1.205 ;
        RECT 10.430 0.900 10.440 1.070 ;
        RECT 10.440 0.900 10.450 1.080 ;
        RECT 10.450 0.900 10.460 1.090 ;
        RECT 10.460 0.900 10.470 1.100 ;
        RECT 10.470 0.900 10.480 1.110 ;
        RECT 10.480 0.900 10.490 1.120 ;
        RECT 10.490 0.900 10.500 1.130 ;
        RECT 10.500 0.900 10.506 1.140 ;
  END 
END FFSDNSRHDMXHT

MACRO FFSDNSRHD2XHT
  CLASS  CORE ;
  FOREIGN FFSDNSRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.990 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.825 1.530 3.245 1.950 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 15.130 1.180 15.480 1.350 ;
        RECT 15.270 0.710 15.300 2.895 ;
        RECT 15.130 0.710 15.300 1.350 ;
        RECT 15.270 1.180 15.365 2.895 ;
        RECT 15.065 2.010 15.365 2.895 ;
        RECT 15.270 1.180 15.480 2.170 ;
        RECT 15.065 2.010 15.480 2.170 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.040 0.720 14.260 1.360 ;
        RECT 14.040 1.190 14.525 1.360 ;
        RECT 14.355 1.190 14.525 2.300 ;
        RECT 14.025 2.130 14.525 2.300 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.255 0.920 1.605 1.425 ;
        RECT 0.825 1.255 1.605 1.425 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.060 1.485 6.230 1.950 ;
        RECT 5.745 1.740 6.230 1.950 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.455 1.610 1.200 1.950 ;
        RECT 0.455 1.675 1.575 1.845 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.955 ;
        RECT 2.535 -0.300 3.515 0.735 ;
        RECT 5.855 -0.300 6.155 1.140 ;
        RECT 8.780 -0.300 8.950 1.020 ;
        RECT 10.820 -0.300 11.120 0.740 ;
        RECT 13.130 -0.300 13.770 1.055 ;
        RECT 14.545 -0.300 14.845 0.715 ;
        RECT 15.650 -0.300 15.820 1.120 ;
        RECT 0.000 -0.300 15.990 0.300 ;
    END
  END GND
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 0.855 2.360 1.675 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 13.155 1.325 13.325 1.840 ;
        RECT 13.155 1.325 13.525 1.540 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 2.715 0.835 3.990 ;
        RECT 2.425 3.045 2.725 3.990 ;
        RECT 3.445 2.830 3.615 3.990 ;
        RECT 6.020 2.995 7.000 3.990 ;
        RECT 8.710 2.995 9.010 3.990 ;
        RECT 10.695 2.960 10.995 3.990 ;
        RECT 12.535 3.015 12.835 3.990 ;
        RECT 13.505 2.975 13.805 3.990 ;
        RECT 14.545 2.975 14.845 3.990 ;
        RECT 15.650 2.230 15.820 3.990 ;
        RECT 0.000 3.390 15.990 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.785 0.275 2.335 ;
        RECT 0.105 0.785 0.405 0.955 ;
        RECT 0.105 2.165 1.250 2.335 ;
        RECT 1.080 2.165 1.250 3.085 ;
        RECT 1.080 2.915 2.035 3.085 ;
        RECT 2.755 1.125 3.620 1.295 ;
        RECT 3.450 1.125 3.620 2.300 ;
        RECT 2.830 2.130 3.620 2.300 ;
        RECT 3.450 1.530 3.820 1.830 ;
        RECT 1.545 0.565 1.955 0.735 ;
        RECT 1.785 0.565 1.955 2.650 ;
        RECT 1.520 2.280 1.955 2.650 ;
        RECT 4.380 0.905 4.550 2.650 ;
        RECT 1.520 2.480 4.550 2.650 ;
        RECT 4.380 2.130 4.680 2.430 ;
        RECT 3.805 1.120 4.170 1.295 ;
        RECT 4.000 0.555 4.170 2.280 ;
        RECT 4.565 0.500 4.865 0.725 ;
        RECT 4.000 0.555 5.555 0.725 ;
        RECT 5.260 1.370 5.430 2.035 ;
        RECT 5.385 0.555 5.555 1.540 ;
        RECT 5.260 1.370 5.555 1.540 ;
        RECT 6.400 0.960 6.610 1.260 ;
        RECT 6.410 0.960 6.610 2.115 ;
        RECT 6.410 1.435 6.710 2.115 ;
        RECT 6.410 1.435 7.330 1.605 ;
        RECT 4.860 0.970 5.030 2.465 ;
        RECT 4.860 0.970 5.205 1.140 ;
        RECT 4.860 2.295 7.325 2.465 ;
        RECT 7.665 1.675 7.860 1.845 ;
        RECT 7.560 1.675 7.570 1.939 ;
        RECT 7.570 1.675 7.580 1.929 ;
        RECT 7.580 1.675 7.590 1.919 ;
        RECT 7.590 1.675 7.600 1.909 ;
        RECT 7.600 1.675 7.610 1.899 ;
        RECT 7.610 1.675 7.620 1.889 ;
        RECT 7.620 1.675 7.630 1.879 ;
        RECT 7.630 1.675 7.640 1.869 ;
        RECT 7.640 1.675 7.650 1.859 ;
        RECT 7.650 1.675 7.660 1.849 ;
        RECT 7.660 1.675 7.666 1.845 ;
        RECT 7.495 1.755 7.505 2.005 ;
        RECT 7.505 1.745 7.515 1.995 ;
        RECT 7.515 1.735 7.525 1.985 ;
        RECT 7.525 1.725 7.535 1.975 ;
        RECT 7.535 1.715 7.545 1.965 ;
        RECT 7.545 1.705 7.555 1.955 ;
        RECT 7.555 1.695 7.561 1.949 ;
        RECT 7.325 1.925 7.335 2.465 ;
        RECT 7.335 1.915 7.345 2.465 ;
        RECT 7.345 1.905 7.355 2.465 ;
        RECT 7.355 1.895 7.365 2.465 ;
        RECT 7.365 1.885 7.375 2.465 ;
        RECT 7.375 1.875 7.385 2.465 ;
        RECT 7.385 1.865 7.395 2.465 ;
        RECT 7.395 1.855 7.405 2.465 ;
        RECT 7.405 1.845 7.415 2.465 ;
        RECT 7.415 1.835 7.425 2.465 ;
        RECT 7.425 1.825 7.435 2.465 ;
        RECT 7.435 1.815 7.445 2.465 ;
        RECT 7.445 1.805 7.455 2.465 ;
        RECT 7.455 1.795 7.465 2.465 ;
        RECT 7.465 1.785 7.475 2.465 ;
        RECT 7.475 1.775 7.485 2.465 ;
        RECT 7.485 1.765 7.495 2.465 ;
        RECT 6.885 1.025 7.185 1.230 ;
        RECT 6.885 1.060 8.220 1.230 ;
        RECT 8.050 1.060 8.220 1.360 ;
        RECT 6.545 0.480 6.845 0.780 ;
        RECT 7.435 0.610 7.605 0.880 ;
        RECT 6.545 0.610 7.605 0.780 ;
        RECT 7.740 2.045 7.950 2.215 ;
        RECT 7.435 0.710 8.570 0.880 ;
        RECT 8.400 0.710 8.570 1.755 ;
        RECT 8.400 1.580 9.250 1.755 ;
        RECT 8.210 1.585 9.250 1.755 ;
        RECT 8.040 1.585 8.050 2.205 ;
        RECT 8.050 1.585 8.060 2.195 ;
        RECT 8.060 1.585 8.070 2.185 ;
        RECT 8.070 1.585 8.080 2.175 ;
        RECT 8.080 1.585 8.090 2.165 ;
        RECT 8.090 1.585 8.100 2.155 ;
        RECT 8.100 1.585 8.110 2.145 ;
        RECT 8.110 1.585 8.120 2.135 ;
        RECT 8.120 1.585 8.130 2.125 ;
        RECT 8.130 1.585 8.140 2.115 ;
        RECT 8.140 1.585 8.150 2.105 ;
        RECT 8.150 1.585 8.160 2.095 ;
        RECT 8.160 1.585 8.170 2.085 ;
        RECT 8.170 1.585 8.180 2.075 ;
        RECT 8.180 1.585 8.190 2.065 ;
        RECT 8.190 1.585 8.200 2.055 ;
        RECT 8.200 1.585 8.210 2.045 ;
        RECT 7.950 2.045 7.960 2.215 ;
        RECT 7.960 2.035 7.970 2.215 ;
        RECT 7.970 2.025 7.980 2.215 ;
        RECT 7.980 2.015 7.990 2.215 ;
        RECT 7.990 2.005 8.000 2.215 ;
        RECT 8.000 1.995 8.010 2.215 ;
        RECT 8.010 1.985 8.020 2.215 ;
        RECT 8.020 1.975 8.030 2.215 ;
        RECT 8.030 1.965 8.040 2.215 ;
        RECT 3.815 2.830 3.985 3.130 ;
        RECT 4.810 2.645 4.980 3.000 ;
        RECT 3.815 2.830 4.980 3.000 ;
        RECT 4.810 2.645 7.880 2.815 ;
        RECT 8.305 2.295 9.315 2.465 ;
        RECT 9.645 2.550 9.975 2.720 ;
        RECT 10.075 1.700 10.085 2.684 ;
        RECT 10.085 1.700 10.095 2.674 ;
        RECT 10.095 1.700 10.105 2.664 ;
        RECT 10.105 1.700 10.115 2.654 ;
        RECT 10.115 1.700 10.125 2.644 ;
        RECT 10.125 1.700 10.135 2.634 ;
        RECT 10.135 1.700 10.145 2.624 ;
        RECT 10.145 1.700 10.155 2.614 ;
        RECT 10.155 1.700 10.165 2.604 ;
        RECT 10.165 1.700 10.175 2.594 ;
        RECT 10.175 1.700 10.185 2.584 ;
        RECT 10.185 1.700 10.195 2.574 ;
        RECT 10.195 1.700 10.205 2.564 ;
        RECT 10.205 1.700 10.215 2.554 ;
        RECT 10.215 1.700 10.225 2.544 ;
        RECT 10.225 1.700 10.235 2.534 ;
        RECT 10.235 1.700 10.245 2.524 ;
        RECT 10.050 2.475 10.060 2.709 ;
        RECT 10.060 2.465 10.070 2.699 ;
        RECT 10.070 2.455 10.076 2.695 ;
        RECT 9.975 2.550 9.985 2.720 ;
        RECT 9.985 2.540 9.995 2.720 ;
        RECT 9.995 2.530 10.005 2.720 ;
        RECT 10.005 2.520 10.015 2.720 ;
        RECT 10.015 2.510 10.025 2.720 ;
        RECT 10.025 2.500 10.035 2.720 ;
        RECT 10.035 2.490 10.045 2.720 ;
        RECT 10.045 2.480 10.051 2.720 ;
        RECT 9.570 2.485 9.580 2.719 ;
        RECT 9.580 2.495 9.590 2.719 ;
        RECT 9.590 2.505 9.600 2.719 ;
        RECT 9.600 2.515 9.610 2.719 ;
        RECT 9.610 2.525 9.620 2.719 ;
        RECT 9.620 2.535 9.630 2.719 ;
        RECT 9.630 2.545 9.640 2.719 ;
        RECT 9.640 2.550 9.646 2.720 ;
        RECT 9.390 2.305 9.400 2.539 ;
        RECT 9.400 2.315 9.410 2.549 ;
        RECT 9.410 2.325 9.420 2.559 ;
        RECT 9.420 2.335 9.430 2.569 ;
        RECT 9.430 2.345 9.440 2.579 ;
        RECT 9.440 2.355 9.450 2.589 ;
        RECT 9.450 2.365 9.460 2.599 ;
        RECT 9.460 2.375 9.470 2.609 ;
        RECT 9.470 2.385 9.480 2.619 ;
        RECT 9.480 2.395 9.490 2.629 ;
        RECT 9.490 2.405 9.500 2.639 ;
        RECT 9.500 2.415 9.510 2.649 ;
        RECT 9.510 2.425 9.520 2.659 ;
        RECT 9.520 2.435 9.530 2.669 ;
        RECT 9.530 2.445 9.540 2.679 ;
        RECT 9.540 2.455 9.550 2.689 ;
        RECT 9.550 2.465 9.560 2.699 ;
        RECT 9.560 2.475 9.570 2.709 ;
        RECT 9.315 2.295 9.325 2.465 ;
        RECT 9.325 2.295 9.335 2.475 ;
        RECT 9.335 2.295 9.345 2.485 ;
        RECT 9.345 2.295 9.355 2.495 ;
        RECT 9.355 2.295 9.365 2.505 ;
        RECT 9.365 2.295 9.375 2.515 ;
        RECT 9.375 2.295 9.385 2.525 ;
        RECT 9.385 2.295 9.391 2.535 ;
        RECT 8.230 2.295 8.240 2.529 ;
        RECT 8.240 2.295 8.250 2.519 ;
        RECT 8.250 2.295 8.260 2.509 ;
        RECT 8.260 2.295 8.270 2.499 ;
        RECT 8.270 2.295 8.280 2.489 ;
        RECT 8.280 2.295 8.290 2.479 ;
        RECT 8.290 2.295 8.300 2.469 ;
        RECT 8.300 2.295 8.306 2.465 ;
        RECT 7.955 2.570 7.965 2.804 ;
        RECT 7.965 2.560 7.975 2.794 ;
        RECT 7.975 2.550 7.985 2.784 ;
        RECT 7.985 2.540 7.995 2.774 ;
        RECT 7.995 2.530 8.005 2.764 ;
        RECT 8.005 2.520 8.015 2.754 ;
        RECT 8.015 2.510 8.025 2.744 ;
        RECT 8.025 2.500 8.035 2.734 ;
        RECT 8.035 2.490 8.045 2.724 ;
        RECT 8.045 2.480 8.055 2.714 ;
        RECT 8.055 2.470 8.065 2.704 ;
        RECT 8.065 2.460 8.075 2.694 ;
        RECT 8.075 2.450 8.085 2.684 ;
        RECT 8.085 2.440 8.095 2.674 ;
        RECT 8.095 2.430 8.105 2.664 ;
        RECT 8.105 2.420 8.115 2.654 ;
        RECT 8.115 2.410 8.125 2.644 ;
        RECT 8.125 2.400 8.135 2.634 ;
        RECT 8.135 2.390 8.145 2.624 ;
        RECT 8.145 2.380 8.155 2.614 ;
        RECT 8.155 2.370 8.165 2.604 ;
        RECT 8.165 2.360 8.175 2.594 ;
        RECT 8.175 2.350 8.185 2.584 ;
        RECT 8.185 2.340 8.195 2.574 ;
        RECT 8.195 2.330 8.205 2.564 ;
        RECT 8.205 2.320 8.215 2.554 ;
        RECT 8.215 2.310 8.225 2.544 ;
        RECT 8.225 2.300 8.231 2.540 ;
        RECT 7.880 2.645 7.890 2.815 ;
        RECT 7.890 2.635 7.900 2.815 ;
        RECT 7.900 2.625 7.910 2.815 ;
        RECT 7.910 2.615 7.920 2.815 ;
        RECT 7.920 2.605 7.930 2.815 ;
        RECT 7.930 2.595 7.940 2.815 ;
        RECT 7.940 2.585 7.950 2.815 ;
        RECT 7.950 2.575 7.956 2.815 ;
        RECT 8.020 3.040 8.360 3.210 ;
        RECT 8.485 2.645 8.530 3.210 ;
        RECT 8.580 2.645 9.125 2.815 ;
        RECT 9.470 2.915 10.240 3.085 ;
        RECT 10.130 1.285 10.425 1.455 ;
        RECT 10.425 1.285 10.435 2.965 ;
        RECT 10.435 1.285 10.445 2.955 ;
        RECT 10.445 1.285 10.455 2.945 ;
        RECT 10.455 1.285 10.465 2.935 ;
        RECT 10.465 1.285 10.475 2.925 ;
        RECT 10.475 1.285 10.485 2.915 ;
        RECT 10.485 1.285 10.495 2.905 ;
        RECT 10.495 1.285 10.505 2.895 ;
        RECT 10.505 1.285 10.515 2.885 ;
        RECT 10.515 1.285 10.525 2.875 ;
        RECT 10.525 1.285 10.535 2.865 ;
        RECT 10.535 1.285 10.545 2.855 ;
        RECT 10.545 1.285 10.555 2.845 ;
        RECT 10.555 1.285 10.565 2.835 ;
        RECT 10.565 1.285 10.575 2.825 ;
        RECT 10.575 1.285 10.585 2.815 ;
        RECT 10.585 1.285 10.595 2.805 ;
        RECT 10.315 2.840 10.325 3.074 ;
        RECT 10.325 2.830 10.335 3.064 ;
        RECT 10.335 2.820 10.345 3.054 ;
        RECT 10.345 2.810 10.355 3.044 ;
        RECT 10.355 2.800 10.365 3.034 ;
        RECT 10.365 2.790 10.375 3.024 ;
        RECT 10.375 2.780 10.385 3.014 ;
        RECT 10.385 2.770 10.395 3.004 ;
        RECT 10.395 2.760 10.405 2.994 ;
        RECT 10.405 2.750 10.415 2.984 ;
        RECT 10.415 2.740 10.425 2.974 ;
        RECT 10.240 2.915 10.250 3.085 ;
        RECT 10.250 2.905 10.260 3.085 ;
        RECT 10.260 2.895 10.270 3.085 ;
        RECT 10.270 2.885 10.280 3.085 ;
        RECT 10.280 2.875 10.290 3.085 ;
        RECT 10.290 2.865 10.300 3.085 ;
        RECT 10.300 2.855 10.310 3.085 ;
        RECT 10.310 2.845 10.316 3.085 ;
        RECT 9.395 2.850 9.405 3.084 ;
        RECT 9.405 2.860 9.415 3.084 ;
        RECT 9.415 2.870 9.425 3.084 ;
        RECT 9.425 2.880 9.435 3.084 ;
        RECT 9.435 2.890 9.445 3.084 ;
        RECT 9.445 2.900 9.455 3.084 ;
        RECT 9.455 2.910 9.465 3.084 ;
        RECT 9.465 2.915 9.471 3.085 ;
        RECT 9.200 2.655 9.210 2.889 ;
        RECT 9.210 2.665 9.220 2.899 ;
        RECT 9.220 2.675 9.230 2.909 ;
        RECT 9.230 2.685 9.240 2.919 ;
        RECT 9.240 2.695 9.250 2.929 ;
        RECT 9.250 2.705 9.260 2.939 ;
        RECT 9.260 2.715 9.270 2.949 ;
        RECT 9.270 2.725 9.280 2.959 ;
        RECT 9.280 2.735 9.290 2.969 ;
        RECT 9.290 2.745 9.300 2.979 ;
        RECT 9.300 2.755 9.310 2.989 ;
        RECT 9.310 2.765 9.320 2.999 ;
        RECT 9.320 2.775 9.330 3.009 ;
        RECT 9.330 2.785 9.340 3.019 ;
        RECT 9.340 2.795 9.350 3.029 ;
        RECT 9.350 2.805 9.360 3.039 ;
        RECT 9.360 2.815 9.370 3.049 ;
        RECT 9.370 2.825 9.380 3.059 ;
        RECT 9.380 2.835 9.390 3.069 ;
        RECT 9.390 2.840 9.396 3.080 ;
        RECT 9.125 2.645 9.135 2.815 ;
        RECT 9.135 2.645 9.145 2.825 ;
        RECT 9.145 2.645 9.155 2.835 ;
        RECT 9.155 2.645 9.165 2.845 ;
        RECT 9.165 2.645 9.175 2.855 ;
        RECT 9.175 2.645 9.185 2.865 ;
        RECT 9.185 2.645 9.195 2.875 ;
        RECT 9.195 2.645 9.201 2.885 ;
        RECT 8.530 2.645 8.540 2.855 ;
        RECT 8.540 2.645 8.550 2.845 ;
        RECT 8.550 2.645 8.560 2.835 ;
        RECT 8.560 2.645 8.570 2.825 ;
        RECT 8.570 2.645 8.580 2.815 ;
        RECT 8.360 2.770 8.370 3.210 ;
        RECT 8.370 2.760 8.380 3.210 ;
        RECT 8.380 2.750 8.390 3.210 ;
        RECT 8.390 2.740 8.400 3.210 ;
        RECT 8.400 2.730 8.410 3.210 ;
        RECT 8.410 2.720 8.420 3.210 ;
        RECT 8.420 2.710 8.430 3.210 ;
        RECT 8.430 2.700 8.440 3.210 ;
        RECT 8.440 2.690 8.450 3.210 ;
        RECT 8.450 2.680 8.460 3.210 ;
        RECT 8.460 2.670 8.470 3.210 ;
        RECT 8.470 2.660 8.480 3.210 ;
        RECT 8.480 2.650 8.486 3.210 ;
        RECT 11.525 1.565 12.200 1.735 ;
        RECT 12.030 1.565 12.200 2.070 ;
        RECT 12.030 1.900 12.625 2.070 ;
        RECT 11.345 0.545 12.855 0.715 ;
        RECT 11.125 1.125 11.295 1.425 ;
        RECT 11.985 2.275 12.160 2.585 ;
        RECT 11.615 2.415 12.160 2.585 ;
        RECT 11.955 0.895 12.255 1.370 ;
        RECT 11.125 1.200 12.975 1.370 ;
        RECT 12.805 1.200 12.975 2.445 ;
        RECT 11.985 2.275 13.835 2.445 ;
        RECT 13.665 1.780 13.835 2.445 ;
        RECT 13.940 1.540 14.110 1.950 ;
        RECT 13.665 1.780 14.110 1.950 ;
        RECT 9.710 0.720 9.880 1.105 ;
        RECT 9.725 0.935 9.895 2.370 ;
        RECT 9.710 0.935 10.945 1.105 ;
        RECT 10.775 0.935 10.945 2.215 ;
        RECT 11.265 2.045 11.435 2.935 ;
        RECT 10.775 2.045 11.735 2.215 ;
        RECT 11.265 2.765 12.280 2.935 ;
        RECT 14.705 1.530 14.875 2.795 ;
        RECT 12.495 2.625 14.875 2.795 ;
        RECT 14.705 1.530 15.090 1.830 ;
        RECT 12.420 2.625 12.430 2.859 ;
        RECT 12.430 2.625 12.440 2.849 ;
        RECT 12.440 2.625 12.450 2.839 ;
        RECT 12.450 2.625 12.460 2.829 ;
        RECT 12.460 2.625 12.470 2.819 ;
        RECT 12.470 2.625 12.480 2.809 ;
        RECT 12.480 2.625 12.490 2.799 ;
        RECT 12.490 2.625 12.496 2.795 ;
        RECT 12.355 2.690 12.365 2.924 ;
        RECT 12.365 2.680 12.375 2.914 ;
        RECT 12.375 2.670 12.385 2.904 ;
        RECT 12.385 2.660 12.395 2.894 ;
        RECT 12.395 2.650 12.405 2.884 ;
        RECT 12.405 2.640 12.415 2.874 ;
        RECT 12.415 2.630 12.421 2.870 ;
        RECT 12.280 2.765 12.290 2.935 ;
        RECT 12.290 2.755 12.300 2.935 ;
        RECT 12.300 2.745 12.310 2.935 ;
        RECT 12.310 2.735 12.320 2.935 ;
        RECT 12.320 2.725 12.330 2.935 ;
        RECT 12.330 2.715 12.340 2.935 ;
        RECT 12.340 2.705 12.350 2.935 ;
        RECT 12.350 2.695 12.356 2.935 ;
  END 
END FFSDNSRHD2XHT

MACRO FFSDNSRHD1XHT
  CLASS  CORE ;
  FOREIGN FFSDNSRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.760 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.965 1.550 3.305 2.015 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.970 0.915 14.575 1.130 ;
        RECT 14.405 0.720 14.575 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.110 0.920 13.535 1.130 ;
        RECT 13.365 0.720 13.535 1.360 ;
        RECT 13.365 1.150 13.780 1.360 ;
        RECT 13.610 1.150 13.780 2.215 ;
        RECT 13.300 2.045 13.780 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.325 0.855 1.545 1.455 ;
        RECT 0.855 1.285 1.545 1.455 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.760 1.735 6.385 2.110 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.455 1.635 0.625 1.945 ;
        RECT 0.455 1.770 1.290 1.945 ;
        RECT 0.815 1.770 1.290 2.365 ;
        RECT 1.370 1.635 1.540 1.940 ;
        RECT 0.455 1.770 1.540 1.940 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.060 ;
        RECT 2.595 -0.300 2.895 0.785 ;
        RECT 3.295 -0.300 3.595 0.745 ;
        RECT 5.970 -0.300 6.270 1.130 ;
        RECT 8.765 -0.300 8.935 1.220 ;
        RECT 10.745 -0.300 11.045 0.860 ;
        RECT 12.715 -0.300 13.015 0.695 ;
        RECT 13.820 -0.300 14.120 0.715 ;
        RECT 0.000 -0.300 14.760 0.300 ;
    END
  END GND
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.290 1.610 2.775 2.015 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 12.305 1.540 12.760 1.950 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.545 2.970 0.845 3.990 ;
        RECT 2.505 2.995 3.485 3.990 ;
        RECT 6.180 2.995 7.160 3.990 ;
        RECT 8.700 2.995 9.000 3.990 ;
        RECT 10.800 2.365 11.100 3.990 ;
        RECT 12.665 2.830 12.965 3.990 ;
        RECT 13.820 2.975 14.120 3.990 ;
        RECT 0.000 3.390 14.760 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.125 0.340 2.425 ;
        RECT 0.105 0.890 0.275 2.425 ;
        RECT 0.170 2.125 0.340 2.775 ;
        RECT 0.105 0.890 0.405 1.060 ;
        RECT 0.170 2.605 1.305 2.775 ;
        RECT 1.135 2.605 1.305 3.150 ;
        RECT 1.135 2.980 1.995 3.150 ;
        RECT 2.825 1.125 3.750 1.295 ;
        RECT 3.580 1.125 3.750 2.365 ;
        RECT 2.825 2.195 3.750 2.365 ;
        RECT 1.740 0.825 1.985 1.125 ;
        RECT 1.815 0.825 1.985 2.715 ;
        RECT 1.580 2.200 1.985 2.715 ;
        RECT 4.445 1.045 4.615 2.715 ;
        RECT 1.580 2.545 4.615 2.715 ;
        RECT 3.930 0.695 4.100 2.280 ;
        RECT 3.930 0.695 5.545 0.865 ;
        RECT 5.375 0.695 5.545 2.245 ;
        RECT 6.555 0.895 6.755 1.195 ;
        RECT 6.585 0.895 6.755 2.115 ;
        RECT 6.585 1.445 7.345 1.745 ;
        RECT 5.025 1.045 5.195 2.595 ;
        RECT 5.025 2.425 5.680 2.595 ;
        RECT 7.525 1.680 7.695 2.465 ;
        RECT 5.885 2.295 7.695 2.465 ;
        RECT 7.775 1.550 7.945 1.850 ;
        RECT 7.525 1.680 7.945 1.850 ;
        RECT 5.810 2.295 5.820 2.529 ;
        RECT 5.820 2.295 5.830 2.519 ;
        RECT 5.830 2.295 5.840 2.509 ;
        RECT 5.840 2.295 5.850 2.499 ;
        RECT 5.850 2.295 5.860 2.489 ;
        RECT 5.860 2.295 5.870 2.479 ;
        RECT 5.870 2.295 5.880 2.469 ;
        RECT 5.880 2.295 5.886 2.465 ;
        RECT 5.755 2.350 5.765 2.584 ;
        RECT 5.765 2.340 5.775 2.574 ;
        RECT 5.775 2.330 5.785 2.564 ;
        RECT 5.785 2.320 5.795 2.554 ;
        RECT 5.795 2.310 5.805 2.544 ;
        RECT 5.805 2.300 5.811 2.540 ;
        RECT 5.680 2.425 5.690 2.595 ;
        RECT 5.690 2.415 5.700 2.595 ;
        RECT 5.700 2.405 5.710 2.595 ;
        RECT 5.710 2.395 5.720 2.595 ;
        RECT 5.720 2.385 5.730 2.595 ;
        RECT 5.730 2.375 5.740 2.595 ;
        RECT 5.740 2.365 5.750 2.595 ;
        RECT 5.750 2.355 5.756 2.595 ;
        RECT 7.000 0.960 7.300 1.215 ;
        RECT 7.000 1.045 8.235 1.215 ;
        RECT 8.065 1.045 8.235 1.345 ;
        RECT 7.890 2.045 8.015 2.215 ;
        RECT 8.125 1.535 8.190 2.215 ;
        RECT 6.630 0.525 8.585 0.695 ;
        RECT 8.415 0.525 8.585 1.705 ;
        RECT 8.295 1.535 9.210 1.705 ;
        RECT 8.190 1.535 8.200 2.105 ;
        RECT 8.200 1.535 8.210 2.095 ;
        RECT 8.210 1.535 8.220 2.085 ;
        RECT 8.220 1.535 8.230 2.075 ;
        RECT 8.230 1.535 8.240 2.065 ;
        RECT 8.240 1.535 8.250 2.055 ;
        RECT 8.250 1.535 8.260 2.045 ;
        RECT 8.260 1.535 8.270 2.035 ;
        RECT 8.270 1.535 8.280 2.025 ;
        RECT 8.280 1.535 8.290 2.015 ;
        RECT 8.290 1.535 8.296 2.009 ;
        RECT 8.015 2.045 8.025 2.215 ;
        RECT 8.025 2.035 8.035 2.215 ;
        RECT 8.035 2.025 8.045 2.215 ;
        RECT 8.045 2.015 8.055 2.215 ;
        RECT 8.055 2.005 8.065 2.215 ;
        RECT 8.065 1.995 8.075 2.215 ;
        RECT 8.075 1.985 8.085 2.215 ;
        RECT 8.085 1.975 8.095 2.215 ;
        RECT 8.095 1.965 8.105 2.215 ;
        RECT 8.105 1.955 8.115 2.215 ;
        RECT 8.115 1.945 8.125 2.215 ;
        RECT 3.685 2.895 5.710 3.065 ;
        RECT 7.875 2.415 8.045 2.815 ;
        RECT 6.035 2.645 8.045 2.815 ;
        RECT 7.875 2.415 8.250 2.585 ;
        RECT 8.445 2.295 9.260 2.465 ;
        RECT 10.100 1.810 10.270 2.565 ;
        RECT 9.435 2.395 10.270 2.565 ;
        RECT 9.360 2.330 9.370 2.564 ;
        RECT 9.370 2.340 9.380 2.564 ;
        RECT 9.380 2.350 9.390 2.564 ;
        RECT 9.390 2.360 9.400 2.564 ;
        RECT 9.400 2.370 9.410 2.564 ;
        RECT 9.410 2.380 9.420 2.564 ;
        RECT 9.420 2.390 9.430 2.564 ;
        RECT 9.430 2.395 9.436 2.565 ;
        RECT 9.335 2.305 9.345 2.539 ;
        RECT 9.345 2.315 9.355 2.549 ;
        RECT 9.355 2.320 9.361 2.560 ;
        RECT 9.260 2.295 9.270 2.465 ;
        RECT 9.270 2.295 9.280 2.475 ;
        RECT 9.280 2.295 9.290 2.485 ;
        RECT 9.290 2.295 9.300 2.495 ;
        RECT 9.300 2.295 9.310 2.505 ;
        RECT 9.310 2.295 9.320 2.515 ;
        RECT 9.320 2.295 9.330 2.525 ;
        RECT 9.330 2.295 9.336 2.535 ;
        RECT 8.370 2.295 8.380 2.529 ;
        RECT 8.380 2.295 8.390 2.519 ;
        RECT 8.390 2.295 8.400 2.509 ;
        RECT 8.400 2.295 8.410 2.499 ;
        RECT 8.410 2.295 8.420 2.489 ;
        RECT 8.420 2.295 8.430 2.479 ;
        RECT 8.430 2.295 8.440 2.469 ;
        RECT 8.440 2.295 8.446 2.465 ;
        RECT 8.325 2.340 8.335 2.574 ;
        RECT 8.335 2.330 8.345 2.564 ;
        RECT 8.345 2.320 8.355 2.554 ;
        RECT 8.355 2.310 8.365 2.544 ;
        RECT 8.365 2.300 8.371 2.540 ;
        RECT 8.250 2.415 8.260 2.585 ;
        RECT 8.260 2.405 8.270 2.585 ;
        RECT 8.270 2.395 8.280 2.585 ;
        RECT 8.280 2.385 8.290 2.585 ;
        RECT 8.290 2.375 8.300 2.585 ;
        RECT 8.300 2.365 8.310 2.585 ;
        RECT 8.310 2.355 8.320 2.585 ;
        RECT 8.320 2.345 8.326 2.585 ;
        RECT 5.960 2.645 5.970 2.879 ;
        RECT 5.970 2.645 5.980 2.869 ;
        RECT 5.980 2.645 5.990 2.859 ;
        RECT 5.990 2.645 6.000 2.849 ;
        RECT 6.000 2.645 6.010 2.839 ;
        RECT 6.010 2.645 6.020 2.829 ;
        RECT 6.020 2.645 6.030 2.819 ;
        RECT 6.030 2.645 6.036 2.815 ;
        RECT 5.785 2.820 5.795 3.054 ;
        RECT 5.795 2.810 5.805 3.044 ;
        RECT 5.805 2.800 5.815 3.034 ;
        RECT 5.815 2.790 5.825 3.024 ;
        RECT 5.825 2.780 5.835 3.014 ;
        RECT 5.835 2.770 5.845 3.004 ;
        RECT 5.845 2.760 5.855 2.994 ;
        RECT 5.855 2.750 5.865 2.984 ;
        RECT 5.865 2.740 5.875 2.974 ;
        RECT 5.875 2.730 5.885 2.964 ;
        RECT 5.885 2.720 5.895 2.954 ;
        RECT 5.895 2.710 5.905 2.944 ;
        RECT 5.905 2.700 5.915 2.934 ;
        RECT 5.915 2.690 5.925 2.924 ;
        RECT 5.925 2.680 5.935 2.914 ;
        RECT 5.935 2.670 5.945 2.904 ;
        RECT 5.945 2.660 5.955 2.894 ;
        RECT 5.955 2.650 5.961 2.890 ;
        RECT 5.710 2.895 5.720 3.065 ;
        RECT 5.720 2.885 5.730 3.065 ;
        RECT 5.730 2.875 5.740 3.065 ;
        RECT 5.740 2.865 5.750 3.065 ;
        RECT 5.750 2.855 5.760 3.065 ;
        RECT 5.760 2.845 5.770 3.065 ;
        RECT 5.770 2.835 5.780 3.065 ;
        RECT 5.780 2.825 5.786 3.065 ;
        RECT 8.225 2.765 8.395 3.210 ;
        RECT 7.960 3.040 8.395 3.210 ;
        RECT 8.225 2.765 8.425 2.935 ;
        RECT 8.620 2.645 9.105 2.815 ;
        RECT 10.055 1.270 10.295 1.440 ;
        RECT 9.280 2.745 10.450 2.915 ;
        RECT 10.450 1.360 10.460 2.914 ;
        RECT 10.460 1.370 10.470 2.914 ;
        RECT 10.470 1.380 10.480 2.914 ;
        RECT 10.480 1.390 10.490 2.914 ;
        RECT 10.490 1.400 10.500 2.914 ;
        RECT 10.500 1.410 10.510 2.914 ;
        RECT 10.510 1.420 10.520 2.914 ;
        RECT 10.520 1.430 10.530 2.914 ;
        RECT 10.530 1.440 10.540 2.914 ;
        RECT 10.540 1.450 10.550 2.914 ;
        RECT 10.550 1.460 10.560 2.914 ;
        RECT 10.560 1.470 10.570 2.914 ;
        RECT 10.570 1.480 10.580 2.914 ;
        RECT 10.580 1.490 10.590 2.914 ;
        RECT 10.590 1.500 10.600 2.914 ;
        RECT 10.600 1.510 10.610 2.914 ;
        RECT 10.610 1.520 10.620 2.914 ;
        RECT 10.370 1.280 10.380 1.514 ;
        RECT 10.380 1.290 10.390 1.524 ;
        RECT 10.390 1.300 10.400 1.534 ;
        RECT 10.400 1.310 10.410 1.544 ;
        RECT 10.410 1.320 10.420 1.554 ;
        RECT 10.420 1.330 10.430 1.564 ;
        RECT 10.430 1.340 10.440 1.574 ;
        RECT 10.440 1.350 10.450 1.584 ;
        RECT 10.295 1.270 10.305 1.440 ;
        RECT 10.305 1.270 10.315 1.450 ;
        RECT 10.315 1.270 10.325 1.460 ;
        RECT 10.325 1.270 10.335 1.470 ;
        RECT 10.335 1.270 10.345 1.480 ;
        RECT 10.345 1.270 10.355 1.490 ;
        RECT 10.355 1.270 10.365 1.500 ;
        RECT 10.365 1.270 10.371 1.510 ;
        RECT 9.205 2.680 9.215 2.914 ;
        RECT 9.215 2.690 9.225 2.914 ;
        RECT 9.225 2.700 9.235 2.914 ;
        RECT 9.235 2.710 9.245 2.914 ;
        RECT 9.245 2.720 9.255 2.914 ;
        RECT 9.255 2.730 9.265 2.914 ;
        RECT 9.265 2.740 9.275 2.914 ;
        RECT 9.275 2.745 9.281 2.915 ;
        RECT 9.180 2.655 9.190 2.889 ;
        RECT 9.190 2.665 9.200 2.899 ;
        RECT 9.200 2.670 9.206 2.910 ;
        RECT 9.105 2.645 9.115 2.815 ;
        RECT 9.115 2.645 9.125 2.825 ;
        RECT 9.125 2.645 9.135 2.835 ;
        RECT 9.135 2.645 9.145 2.845 ;
        RECT 9.145 2.645 9.155 2.855 ;
        RECT 9.155 2.645 9.165 2.865 ;
        RECT 9.165 2.645 9.175 2.875 ;
        RECT 9.175 2.645 9.181 2.885 ;
        RECT 8.545 2.645 8.555 2.879 ;
        RECT 8.555 2.645 8.565 2.869 ;
        RECT 8.565 2.645 8.575 2.859 ;
        RECT 8.575 2.645 8.585 2.849 ;
        RECT 8.585 2.645 8.595 2.839 ;
        RECT 8.595 2.645 8.605 2.829 ;
        RECT 8.605 2.645 8.615 2.819 ;
        RECT 8.615 2.645 8.621 2.815 ;
        RECT 8.500 2.690 8.510 2.924 ;
        RECT 8.510 2.680 8.520 2.914 ;
        RECT 8.520 2.670 8.530 2.904 ;
        RECT 8.530 2.660 8.540 2.894 ;
        RECT 8.540 2.650 8.546 2.890 ;
        RECT 8.425 2.765 8.435 2.935 ;
        RECT 8.435 2.755 8.445 2.935 ;
        RECT 8.445 2.745 8.455 2.935 ;
        RECT 8.455 2.735 8.465 2.935 ;
        RECT 8.465 2.725 8.475 2.935 ;
        RECT 8.475 2.715 8.485 2.935 ;
        RECT 8.485 2.705 8.495 2.935 ;
        RECT 8.495 2.695 8.501 2.935 ;
        RECT 11.355 0.760 11.525 1.280 ;
        RECT 11.225 1.110 11.525 1.280 ;
        RECT 11.355 0.760 12.435 0.930 ;
        RECT 12.265 0.760 12.435 1.280 ;
        RECT 12.265 1.110 12.565 1.280 ;
        RECT 11.150 1.465 11.320 1.765 ;
        RECT 11.745 1.110 12.045 1.635 ;
        RECT 11.150 1.465 12.045 1.635 ;
        RECT 11.875 1.110 12.045 2.300 ;
        RECT 12.950 1.540 13.120 2.300 ;
        RECT 11.875 2.130 13.120 2.300 ;
        RECT 12.950 1.540 13.430 1.840 ;
        RECT 9.620 0.900 9.790 2.215 ;
        RECT 9.620 2.045 9.920 2.215 ;
        RECT 9.620 0.900 10.430 1.070 ;
        RECT 10.645 1.040 10.970 1.210 ;
        RECT 10.800 1.040 10.970 2.115 ;
        RECT 10.800 1.945 11.530 2.115 ;
        RECT 11.360 1.945 11.530 2.650 ;
        RECT 11.935 2.480 12.235 2.955 ;
        RECT 13.960 1.535 14.130 2.650 ;
        RECT 11.360 2.480 14.130 2.650 ;
        RECT 13.960 1.535 14.225 1.835 ;
        RECT 10.570 0.975 10.580 1.209 ;
        RECT 10.580 0.985 10.590 1.209 ;
        RECT 10.590 0.995 10.600 1.209 ;
        RECT 10.600 1.005 10.610 1.209 ;
        RECT 10.610 1.015 10.620 1.209 ;
        RECT 10.620 1.025 10.630 1.209 ;
        RECT 10.630 1.035 10.640 1.209 ;
        RECT 10.640 1.040 10.646 1.210 ;
        RECT 10.505 0.910 10.515 1.144 ;
        RECT 10.515 0.920 10.525 1.154 ;
        RECT 10.525 0.930 10.535 1.164 ;
        RECT 10.535 0.940 10.545 1.174 ;
        RECT 10.545 0.950 10.555 1.184 ;
        RECT 10.555 0.960 10.565 1.194 ;
        RECT 10.565 0.965 10.571 1.205 ;
        RECT 10.430 0.900 10.440 1.070 ;
        RECT 10.440 0.900 10.450 1.080 ;
        RECT 10.450 0.900 10.460 1.090 ;
        RECT 10.460 0.900 10.470 1.100 ;
        RECT 10.470 0.900 10.480 1.110 ;
        RECT 10.480 0.900 10.490 1.120 ;
        RECT 10.490 0.900 10.500 1.130 ;
        RECT 10.500 0.900 10.506 1.140 ;
  END 
END FFSDNSRHD1XHT

MACRO FFSDNSHDMXHT
  CLASS  CORE ;
  FOREIGN FFSDNSHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.890 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 3.640 1.525 4.110 2.010 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.550 1.060 11.790 1.360 ;
        RECT 11.580 1.060 11.790 2.450 ;
        RECT 11.550 1.980 11.790 2.450 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.510 1.060 10.680 1.360 ;
        RECT 10.510 1.190 10.970 1.360 ;
        RECT 10.760 1.190 10.970 2.240 ;
        RECT 10.445 2.070 10.970 2.240 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.415 -0.300 2.715 0.595 ;
        RECT 3.335 -0.300 3.635 0.595 ;
        RECT 5.925 -0.300 6.225 0.745 ;
        RECT 7.165 -0.300 7.335 0.850 ;
        RECT 9.150 -0.300 9.320 0.640 ;
        RECT 10.965 -0.300 11.265 0.595 ;
        RECT 0.000 -0.300 11.890 0.300 ;
    END
  END GND
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.530 0.500 7.700 1.910 ;
        RECT 6.885 1.610 7.700 1.910 ;
        RECT 7.530 0.500 8.905 0.670 ;
        RECT 8.735 0.500 8.905 1.145 ;
        RECT 9.595 0.540 9.765 1.145 ;
        RECT 8.735 0.920 9.765 1.145 ;
        RECT 9.595 0.540 10.055 0.710 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.305 2.735 2.605 3.990 ;
        RECT 3.335 2.955 3.635 3.990 ;
        RECT 5.855 3.160 6.155 3.990 ;
        RECT 7.100 3.160 7.400 3.990 ;
        RECT 9.170 2.770 9.340 3.990 ;
        RECT 9.810 2.880 9.980 3.990 ;
        RECT 10.965 2.975 11.265 3.990 ;
        RECT 0.000 3.390 11.890 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.555 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.045 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.975 0.775 2.145 1.035 ;
        RECT 1.530 0.865 2.145 1.035 ;
        RECT 1.975 0.775 4.510 0.945 ;
        RECT 4.275 0.540 4.510 0.945 ;
        RECT 4.340 0.540 4.510 2.280 ;
        RECT 5.040 0.900 5.210 2.280 ;
        RECT 5.040 1.675 6.355 1.845 ;
        RECT 6.535 1.060 6.705 2.215 ;
        RECT 6.405 2.045 6.705 2.215 ;
        RECT 6.535 1.060 7.350 1.360 ;
        RECT 2.825 1.125 2.960 2.710 ;
        RECT 2.825 1.125 3.105 1.295 ;
        RECT 3.055 2.540 3.710 2.710 ;
        RECT 4.065 2.810 8.045 2.980 ;
        RECT 3.980 2.735 3.990 2.979 ;
        RECT 3.990 2.745 4.000 2.979 ;
        RECT 4.000 2.755 4.010 2.979 ;
        RECT 4.010 2.765 4.020 2.979 ;
        RECT 4.020 2.775 4.030 2.979 ;
        RECT 4.030 2.785 4.040 2.979 ;
        RECT 4.040 2.795 4.050 2.979 ;
        RECT 4.050 2.805 4.060 2.979 ;
        RECT 4.060 2.810 4.066 2.980 ;
        RECT 3.795 2.550 3.805 2.794 ;
        RECT 3.805 2.560 3.815 2.804 ;
        RECT 3.815 2.570 3.825 2.814 ;
        RECT 3.825 2.580 3.835 2.824 ;
        RECT 3.835 2.590 3.845 2.834 ;
        RECT 3.845 2.600 3.855 2.844 ;
        RECT 3.855 2.610 3.865 2.854 ;
        RECT 3.865 2.620 3.875 2.864 ;
        RECT 3.875 2.630 3.885 2.874 ;
        RECT 3.885 2.640 3.895 2.884 ;
        RECT 3.895 2.650 3.905 2.894 ;
        RECT 3.905 2.660 3.915 2.904 ;
        RECT 3.915 2.670 3.925 2.914 ;
        RECT 3.925 2.680 3.935 2.924 ;
        RECT 3.935 2.690 3.945 2.934 ;
        RECT 3.945 2.700 3.955 2.944 ;
        RECT 3.955 2.710 3.965 2.954 ;
        RECT 3.965 2.720 3.975 2.964 ;
        RECT 3.975 2.725 3.981 2.975 ;
        RECT 3.710 2.540 3.720 2.710 ;
        RECT 3.720 2.540 3.730 2.720 ;
        RECT 3.730 2.540 3.740 2.730 ;
        RECT 3.740 2.540 3.750 2.740 ;
        RECT 3.750 2.540 3.760 2.750 ;
        RECT 3.760 2.540 3.770 2.760 ;
        RECT 3.770 2.540 3.780 2.770 ;
        RECT 3.780 2.540 3.790 2.780 ;
        RECT 3.790 2.540 3.796 2.790 ;
        RECT 2.960 2.105 2.970 2.709 ;
        RECT 2.970 2.115 2.980 2.709 ;
        RECT 2.980 2.125 2.990 2.709 ;
        RECT 2.990 2.135 3.000 2.709 ;
        RECT 3.000 2.145 3.010 2.709 ;
        RECT 3.010 2.155 3.020 2.709 ;
        RECT 3.020 2.165 3.030 2.709 ;
        RECT 3.030 2.175 3.040 2.709 ;
        RECT 3.040 2.185 3.050 2.709 ;
        RECT 3.050 2.190 3.056 2.710 ;
        RECT 2.765 1.125 2.775 2.279 ;
        RECT 2.775 1.125 2.785 2.289 ;
        RECT 2.785 1.125 2.795 2.299 ;
        RECT 2.795 1.125 2.805 2.309 ;
        RECT 2.805 1.125 2.815 2.319 ;
        RECT 2.815 1.125 2.825 2.329 ;
        RECT 3.140 1.525 3.455 1.825 ;
        RECT 3.285 1.125 3.455 2.360 ;
        RECT 3.285 2.190 3.900 2.360 ;
        RECT 3.285 1.125 4.145 1.295 ;
        RECT 4.690 0.535 4.860 2.630 ;
        RECT 4.690 0.535 5.485 0.705 ;
        RECT 7.880 1.645 8.050 2.630 ;
        RECT 7.910 1.245 8.080 1.815 ;
        RECT 7.880 1.645 8.080 1.815 ;
        RECT 4.245 2.460 8.720 2.630 ;
        RECT 8.550 2.460 8.720 2.795 ;
        RECT 4.170 2.395 4.180 2.629 ;
        RECT 4.180 2.405 4.190 2.629 ;
        RECT 4.190 2.415 4.200 2.629 ;
        RECT 4.200 2.425 4.210 2.629 ;
        RECT 4.210 2.435 4.220 2.629 ;
        RECT 4.220 2.445 4.230 2.629 ;
        RECT 4.230 2.455 4.240 2.629 ;
        RECT 4.240 2.460 4.246 2.630 ;
        RECT 4.065 2.290 4.075 2.524 ;
        RECT 4.075 2.300 4.085 2.534 ;
        RECT 4.085 2.310 4.095 2.544 ;
        RECT 4.095 2.320 4.105 2.554 ;
        RECT 4.105 2.330 4.115 2.564 ;
        RECT 4.115 2.340 4.125 2.574 ;
        RECT 4.125 2.350 4.135 2.584 ;
        RECT 4.135 2.360 4.145 2.594 ;
        RECT 4.145 2.370 4.155 2.604 ;
        RECT 4.155 2.380 4.165 2.614 ;
        RECT 4.165 2.385 4.171 2.625 ;
        RECT 3.900 2.190 3.910 2.360 ;
        RECT 3.910 2.190 3.920 2.370 ;
        RECT 3.920 2.190 3.930 2.380 ;
        RECT 3.930 2.190 3.940 2.390 ;
        RECT 3.940 2.190 3.950 2.400 ;
        RECT 3.950 2.190 3.960 2.410 ;
        RECT 3.960 2.190 3.970 2.420 ;
        RECT 3.970 2.190 3.980 2.430 ;
        RECT 3.980 2.190 3.990 2.440 ;
        RECT 3.990 2.190 4.000 2.450 ;
        RECT 4.000 2.190 4.010 2.460 ;
        RECT 4.010 2.190 4.020 2.470 ;
        RECT 4.020 2.190 4.030 2.480 ;
        RECT 4.030 2.190 4.040 2.490 ;
        RECT 4.040 2.190 4.050 2.500 ;
        RECT 4.050 2.190 4.060 2.510 ;
        RECT 4.060 2.190 4.066 2.520 ;
        RECT 8.905 1.325 10.240 1.495 ;
        RECT 10.000 0.890 10.170 1.495 ;
        RECT 10.070 1.325 10.240 2.215 ;
        RECT 9.655 2.045 10.240 2.215 ;
        RECT 10.070 1.540 10.580 1.840 ;
        RECT 8.305 0.885 8.475 2.215 ;
        RECT 8.185 0.885 8.485 1.055 ;
        RECT 8.230 2.045 8.530 2.215 ;
        RECT 9.010 1.675 9.180 2.590 ;
        RECT 8.305 1.675 9.755 1.845 ;
        RECT 11.200 1.540 11.370 2.590 ;
        RECT 9.010 2.420 11.370 2.590 ;
        RECT 11.200 1.540 11.380 1.840 ;
  END 
END FFSDNSHDMXHT

MACRO FFSDNSHDLXHT
  CLASS  CORE ;
  FOREIGN FFSDNSHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.890 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 3.640 1.525 4.130 2.010 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.550 1.060 11.790 1.360 ;
        RECT 11.580 1.060 11.790 2.430 ;
        RECT 11.550 1.980 11.790 2.430 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.540 1.060 10.710 1.360 ;
        RECT 10.540 1.190 10.970 1.360 ;
        RECT 10.760 1.190 10.970 2.240 ;
        RECT 10.445 2.070 10.970 2.240 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.525 2.980 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.435 -0.300 2.735 0.595 ;
        RECT 3.325 -0.300 3.625 0.595 ;
        RECT 5.945 -0.300 6.245 0.745 ;
        RECT 7.165 -0.300 7.335 0.850 ;
        RECT 9.150 -0.300 9.320 0.640 ;
        RECT 10.995 -0.300 11.295 0.745 ;
        RECT 0.000 -0.300 11.890 0.300 ;
    END
  END GND
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.560 0.500 7.730 1.910 ;
        RECT 6.885 1.610 7.730 1.910 ;
        RECT 7.560 0.500 8.905 0.670 ;
        RECT 8.735 0.500 8.905 1.145 ;
        RECT 9.595 0.540 9.765 1.145 ;
        RECT 8.735 0.920 9.765 1.145 ;
        RECT 9.595 0.540 10.005 0.710 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.450 2.510 2.620 3.990 ;
        RECT 3.300 2.890 3.470 3.990 ;
        RECT 5.855 3.160 6.155 3.990 ;
        RECT 7.100 3.160 7.400 3.990 ;
        RECT 9.075 2.770 9.375 3.990 ;
        RECT 9.655 2.880 9.955 3.990 ;
        RECT 10.965 2.770 11.265 3.990 ;
        RECT 0.000 3.390 11.890 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.515 1.350 2.630 ;
        RECT 1.180 0.515 1.525 0.685 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 2.940 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.530 0.865 1.720 1.185 ;
        RECT 2.030 0.775 2.200 1.035 ;
        RECT 1.530 0.865 2.200 1.035 ;
        RECT 2.030 0.775 4.530 0.945 ;
        RECT 4.360 0.775 4.530 2.280 ;
        RECT 5.060 0.900 5.230 2.280 ;
        RECT 5.060 1.675 6.355 1.845 ;
        RECT 6.535 1.060 6.705 2.215 ;
        RECT 6.440 2.045 6.740 2.215 ;
        RECT 6.535 1.060 7.380 1.360 ;
        RECT 2.745 1.980 3.010 2.280 ;
        RECT 2.745 1.125 2.915 2.280 ;
        RECT 2.840 1.980 3.010 2.710 ;
        RECT 2.745 1.125 3.045 1.295 ;
        RECT 2.840 2.540 3.830 2.710 ;
        RECT 3.660 2.540 3.830 2.980 ;
        RECT 3.660 2.810 8.045 2.980 ;
        RECT 3.160 1.525 3.455 1.825 ;
        RECT 3.285 1.125 3.455 2.360 ;
        RECT 3.285 2.190 4.180 2.360 ;
        RECT 3.285 1.125 4.085 1.295 ;
        RECT 4.010 2.190 4.180 2.630 ;
        RECT 4.710 0.535 4.880 2.630 ;
        RECT 4.710 0.535 5.505 0.705 ;
        RECT 7.910 1.210 8.080 2.630 ;
        RECT 4.010 2.460 8.755 2.630 ;
        RECT 10.030 0.890 10.240 1.495 ;
        RECT 8.905 1.325 10.240 1.495 ;
        RECT 10.070 0.890 10.240 2.215 ;
        RECT 9.655 2.045 10.240 2.215 ;
        RECT 10.070 1.540 10.580 1.840 ;
        RECT 8.305 0.890 8.475 2.280 ;
        RECT 8.295 1.980 8.475 2.280 ;
        RECT 8.185 0.890 8.485 1.060 ;
        RECT 9.010 1.675 9.180 2.590 ;
        RECT 8.305 1.675 9.685 1.845 ;
        RECT 11.200 1.610 11.370 2.590 ;
        RECT 9.010 2.420 11.370 2.590 ;
        RECT 11.200 1.610 11.380 1.910 ;
  END 
END FFSDNSHDLXHT

MACRO FFSDNSHD2XHT
  CLASS  CORE ;
  FOREIGN FFSDNSHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.530 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 3.650 1.525 4.140 2.010 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 12.670 0.720 12.840 2.960 ;
        RECT 12.670 1.670 13.020 2.015 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.580 0.720 11.800 2.215 ;
        RECT 11.565 2.045 11.865 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.460 0.410 3.180 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.470 1.325 1.555 1.845 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.600 -0.300 0.770 0.660 ;
        RECT 2.415 -0.300 2.715 0.595 ;
        RECT 3.365 -0.300 3.665 0.595 ;
        RECT 5.925 -0.300 6.225 0.895 ;
        RECT 7.415 -0.300 7.715 0.715 ;
        RECT 9.580 -0.300 9.880 0.740 ;
        RECT 11.045 -0.300 11.345 0.715 ;
        RECT 12.085 -0.300 12.385 1.055 ;
        RECT 13.125 -0.300 13.425 1.055 ;
        RECT 0.000 -0.300 13.530 0.300 ;
    END
  END GND
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.105 1.270 2.600 1.800 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.305 0.960 7.475 1.565 ;
        RECT 7.200 1.265 7.475 1.565 ;
        RECT 7.895 0.605 8.065 1.130 ;
        RECT 7.305 0.960 8.065 1.130 ;
        RECT 7.895 0.605 9.225 0.775 ;
        RECT 9.055 0.605 9.225 1.145 ;
        RECT 9.875 0.920 10.460 1.145 ;
        RECT 10.290 0.515 10.460 1.145 ;
        RECT 9.055 0.975 10.460 1.145 ;
        RECT 10.290 0.515 10.620 0.685 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.610 2.650 0.780 3.990 ;
        RECT 2.460 2.830 2.630 3.990 ;
        RECT 3.310 2.890 3.480 3.990 ;
        RECT 5.950 3.095 6.250 3.990 ;
        RECT 7.080 3.095 7.720 3.990 ;
        RECT 9.465 2.790 9.765 3.990 ;
        RECT 10.655 2.975 11.295 3.990 ;
        RECT 12.085 2.975 12.385 3.990 ;
        RECT 13.125 2.295 13.425 3.990 ;
        RECT 0.000 3.390 13.530 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 0.275 2.215 ;
        RECT 0.105 2.045 1.230 2.215 ;
        RECT 1.025 0.480 1.195 1.145 ;
        RECT 0.105 0.975 1.195 1.145 ;
        RECT 1.060 2.045 1.230 3.085 ;
        RECT 1.025 0.480 1.555 0.650 ;
        RECT 1.060 2.915 2.035 3.085 ;
        RECT 1.530 2.045 1.700 2.620 ;
        RECT 1.750 0.775 1.925 1.080 ;
        RECT 1.465 0.910 1.925 1.080 ;
        RECT 1.755 0.775 1.925 2.215 ;
        RECT 1.465 2.045 1.925 2.215 ;
        RECT 1.750 0.775 4.540 0.945 ;
        RECT 4.370 0.775 4.540 2.280 ;
        RECT 5.070 0.910 5.240 2.280 ;
        RECT 6.145 1.675 6.460 1.865 ;
        RECT 5.070 1.695 6.460 1.865 ;
        RECT 5.665 1.245 5.965 1.515 ;
        RECT 5.665 1.245 7.020 1.415 ;
        RECT 6.850 0.820 7.020 2.215 ;
        RECT 6.500 2.045 7.020 2.215 ;
        RECT 6.850 0.820 7.080 1.120 ;
        RECT 7.695 1.610 7.865 1.915 ;
        RECT 6.850 1.745 7.865 1.915 ;
        RECT 2.795 1.980 3.050 2.280 ;
        RECT 2.795 1.125 2.990 2.280 ;
        RECT 2.880 1.980 3.050 2.710 ;
        RECT 2.795 1.125 3.115 1.295 ;
        RECT 2.880 2.540 3.840 2.710 ;
        RECT 3.670 2.540 3.840 3.035 ;
        RECT 3.670 2.865 5.565 3.035 ;
        RECT 5.805 2.745 8.510 2.915 ;
        RECT 8.330 2.745 8.510 3.185 ;
        RECT 8.330 3.015 8.950 3.185 ;
        RECT 5.685 2.745 5.695 3.025 ;
        RECT 5.695 2.745 5.705 3.015 ;
        RECT 5.705 2.745 5.715 3.005 ;
        RECT 5.715 2.745 5.725 2.995 ;
        RECT 5.725 2.745 5.735 2.985 ;
        RECT 5.735 2.745 5.745 2.975 ;
        RECT 5.745 2.745 5.755 2.965 ;
        RECT 5.755 2.745 5.765 2.955 ;
        RECT 5.765 2.745 5.775 2.945 ;
        RECT 5.775 2.745 5.785 2.935 ;
        RECT 5.785 2.745 5.795 2.925 ;
        RECT 5.795 2.745 5.805 2.915 ;
        RECT 5.565 2.865 5.575 3.035 ;
        RECT 5.575 2.855 5.585 3.035 ;
        RECT 5.585 2.845 5.595 3.035 ;
        RECT 5.595 2.835 5.605 3.035 ;
        RECT 5.605 2.825 5.615 3.035 ;
        RECT 5.615 2.815 5.625 3.035 ;
        RECT 5.625 2.805 5.635 3.035 ;
        RECT 5.635 2.795 5.645 3.035 ;
        RECT 5.645 2.785 5.655 3.035 ;
        RECT 5.655 2.775 5.665 3.035 ;
        RECT 5.665 2.765 5.675 3.035 ;
        RECT 5.675 2.755 5.685 3.035 ;
        RECT 3.170 1.525 3.465 1.825 ;
        RECT 3.295 1.125 3.465 2.360 ;
        RECT 3.295 2.190 4.190 2.360 ;
        RECT 3.295 1.125 4.095 1.295 ;
        RECT 4.020 2.190 4.190 2.685 ;
        RECT 4.720 0.535 4.890 2.685 ;
        RECT 4.020 2.515 5.305 2.685 ;
        RECT 4.720 0.535 5.485 0.705 ;
        RECT 8.175 1.290 8.345 2.565 ;
        RECT 5.545 2.395 9.040 2.565 ;
        RECT 8.870 2.395 9.040 2.770 ;
        RECT 5.425 2.395 5.435 2.675 ;
        RECT 5.435 2.395 5.445 2.665 ;
        RECT 5.445 2.395 5.455 2.655 ;
        RECT 5.455 2.395 5.465 2.645 ;
        RECT 5.465 2.395 5.475 2.635 ;
        RECT 5.475 2.395 5.485 2.625 ;
        RECT 5.485 2.395 5.495 2.615 ;
        RECT 5.495 2.395 5.505 2.605 ;
        RECT 5.505 2.395 5.515 2.595 ;
        RECT 5.515 2.395 5.525 2.585 ;
        RECT 5.525 2.395 5.535 2.575 ;
        RECT 5.535 2.395 5.545 2.565 ;
        RECT 5.305 2.515 5.315 2.685 ;
        RECT 5.315 2.505 5.325 2.685 ;
        RECT 5.325 2.495 5.335 2.685 ;
        RECT 5.335 2.485 5.345 2.685 ;
        RECT 5.345 2.475 5.355 2.685 ;
        RECT 5.355 2.465 5.365 2.685 ;
        RECT 5.365 2.455 5.375 2.685 ;
        RECT 5.375 2.445 5.385 2.685 ;
        RECT 5.385 2.435 5.395 2.685 ;
        RECT 5.395 2.425 5.405 2.685 ;
        RECT 5.405 2.415 5.415 2.685 ;
        RECT 5.415 2.405 5.425 2.685 ;
        RECT 9.275 1.325 10.810 1.495 ;
        RECT 10.640 1.060 10.810 2.215 ;
        RECT 10.025 2.045 10.810 2.215 ;
        RECT 10.640 1.585 11.400 1.755 ;
        RECT 8.535 0.955 8.835 1.125 ;
        RECT 8.620 0.955 8.835 2.215 ;
        RECT 8.600 2.045 8.900 2.215 ;
        RECT 9.675 1.675 9.845 2.565 ;
        RECT 8.620 1.675 10.090 1.845 ;
        RECT 12.320 1.525 12.490 2.565 ;
        RECT 9.675 2.395 12.490 2.565 ;
  END 
END FFSDNSHD2XHT

MACRO FFSDNSHD1XHT
  CLASS  CORE ;
  FOREIGN FFSDNSHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.890 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 3.650 1.525 4.140 2.010 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.550 0.720 11.790 1.360 ;
        RECT 11.620 0.720 11.790 2.960 ;
        RECT 11.550 1.980 11.790 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.510 0.720 10.680 1.360 ;
        RECT 10.510 1.190 10.970 1.360 ;
        RECT 10.760 1.190 10.970 2.240 ;
        RECT 10.445 2.070 10.970 2.240 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.460 0.410 3.180 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.470 1.325 1.555 1.845 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.415 -0.300 2.715 0.595 ;
        RECT 3.365 -0.300 3.665 0.595 ;
        RECT 6.760 -0.300 7.335 0.780 ;
        RECT 9.080 -0.300 9.250 0.640 ;
        RECT 10.965 -0.300 11.265 0.715 ;
        RECT 0.000 -0.300 11.890 0.300 ;
    END
  END GND
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.210 2.500 2.105 ;
    END
  END TI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.530 0.605 7.700 1.910 ;
        RECT 6.885 1.610 7.700 1.910 ;
        RECT 7.530 0.605 8.900 0.775 ;
        RECT 8.730 0.605 8.900 1.145 ;
        RECT 9.595 0.535 9.765 1.145 ;
        RECT 8.730 0.920 9.765 1.145 ;
        RECT 9.595 0.535 10.055 0.705 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.610 2.715 0.780 3.990 ;
        RECT 2.395 2.895 2.695 3.990 ;
        RECT 3.310 2.890 3.480 3.990 ;
        RECT 5.855 3.160 6.155 3.990 ;
        RECT 7.100 3.160 7.400 3.990 ;
        RECT 9.105 2.770 9.405 3.990 ;
        RECT 9.745 2.940 10.045 3.990 ;
        RECT 10.965 2.975 11.265 3.990 ;
        RECT 0.000 3.390 11.890 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 0.275 2.215 ;
        RECT 0.105 2.045 1.240 2.215 ;
        RECT 1.070 2.045 1.240 3.130 ;
        RECT 1.085 0.480 1.255 1.145 ;
        RECT 0.105 0.975 1.255 1.145 ;
        RECT 1.085 0.480 1.555 0.650 ;
        RECT 1.070 2.960 1.985 3.130 ;
        RECT 1.530 2.045 1.700 2.620 ;
        RECT 1.750 0.775 1.925 1.080 ;
        RECT 1.465 0.910 1.925 1.080 ;
        RECT 1.755 0.775 1.925 2.215 ;
        RECT 1.465 2.045 1.925 2.215 ;
        RECT 1.750 0.775 4.540 0.945 ;
        RECT 4.370 0.775 4.540 2.280 ;
        RECT 5.070 0.900 5.240 2.280 ;
        RECT 5.070 1.675 6.355 1.845 ;
        RECT 6.535 1.060 6.705 2.215 ;
        RECT 6.405 2.045 6.705 2.215 ;
        RECT 6.535 1.060 7.350 1.360 ;
        RECT 2.810 1.980 3.050 2.280 ;
        RECT 2.810 1.125 2.990 2.280 ;
        RECT 2.880 1.980 3.050 2.710 ;
        RECT 2.810 1.125 3.115 1.295 ;
        RECT 2.880 2.540 3.840 2.710 ;
        RECT 3.670 2.540 3.840 2.980 ;
        RECT 3.670 2.810 8.205 2.980 ;
        RECT 3.170 1.525 3.465 1.825 ;
        RECT 3.295 1.125 3.465 2.360 ;
        RECT 3.295 2.190 4.190 2.360 ;
        RECT 3.295 1.125 4.095 1.295 ;
        RECT 4.020 2.190 4.190 2.630 ;
        RECT 4.720 0.535 4.890 2.630 ;
        RECT 4.720 0.535 5.485 0.705 ;
        RECT 7.880 1.645 8.050 2.630 ;
        RECT 7.910 1.245 8.080 1.815 ;
        RECT 7.880 1.645 8.080 1.815 ;
        RECT 4.020 2.460 8.720 2.630 ;
        RECT 8.550 2.460 8.720 2.795 ;
        RECT 8.905 1.325 10.240 1.495 ;
        RECT 10.000 0.890 10.170 1.495 ;
        RECT 10.070 1.325 10.240 2.215 ;
        RECT 9.655 2.045 10.240 2.215 ;
        RECT 10.070 1.540 10.580 1.840 ;
        RECT 8.215 0.955 8.520 1.125 ;
        RECT 8.350 0.955 8.520 2.215 ;
        RECT 8.350 1.675 8.530 2.215 ;
        RECT 8.230 2.045 8.530 2.215 ;
        RECT 9.010 1.675 9.180 2.590 ;
        RECT 8.350 1.675 9.755 1.845 ;
        RECT 11.200 1.610 11.370 2.590 ;
        RECT 9.010 2.420 11.370 2.590 ;
        RECT 11.200 1.610 11.380 1.910 ;
  END 
END FFSDNSHD1XHT

MACRO FFSDNRHDMXHT
  CLASS  CORE ;
  FOREIGN FFSDNRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.120 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 3.635 1.525 4.110 2.010 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 12.780 1.060 13.020 1.360 ;
        RECT 12.850 1.060 13.020 2.445 ;
        RECT 12.780 1.980 13.020 2.445 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.580 0.860 11.910 1.470 ;
        RECT 11.580 1.300 12.250 1.470 ;
        RECT 12.080 1.300 12.250 2.215 ;
        RECT 11.675 2.045 12.250 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 8.030 1.610 8.510 2.010 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.415 -0.300 2.715 0.595 ;
        RECT 3.385 -0.300 3.685 0.595 ;
        RECT 5.895 -0.300 6.195 0.595 ;
        RECT 7.035 -0.300 7.335 0.595 ;
        RECT 8.125 -0.300 8.295 0.810 ;
        RECT 10.065 -0.300 10.365 0.525 ;
        RECT 11.195 -0.300 11.495 0.530 ;
        RECT 12.195 -0.300 12.495 0.595 ;
        RECT 0.000 -0.300 13.120 0.300 ;
    END
  END GND
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.315 2.670 2.615 3.990 ;
        RECT 3.335 2.890 3.635 3.990 ;
        RECT 6.035 3.195 6.335 3.990 ;
        RECT 8.165 3.195 8.465 3.990 ;
        RECT 10.165 2.810 10.465 3.990 ;
        RECT 12.195 2.975 12.495 3.990 ;
        RECT 0.000 3.390 13.120 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.555 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.150 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.980 0.775 2.150 1.035 ;
        RECT 1.530 0.865 2.150 1.035 ;
        RECT 1.980 0.775 4.510 0.945 ;
        RECT 4.275 0.590 4.510 0.945 ;
        RECT 4.340 0.590 4.510 2.280 ;
        RECT 5.040 0.910 5.210 2.280 ;
        RECT 6.235 1.675 6.535 1.865 ;
        RECT 5.040 1.695 6.535 1.865 ;
        RECT 5.685 1.325 5.985 1.515 ;
        RECT 6.510 0.775 6.680 1.495 ;
        RECT 5.685 1.325 6.885 1.495 ;
        RECT 6.715 1.325 6.885 2.215 ;
        RECT 6.715 2.045 7.255 2.215 ;
        RECT 7.540 0.480 7.710 0.945 ;
        RECT 6.510 0.775 7.710 0.945 ;
        RECT 2.795 1.125 2.960 2.710 ;
        RECT 2.795 1.125 3.105 1.295 ;
        RECT 2.990 2.540 3.750 2.710 ;
        RECT 8.460 2.745 8.630 3.015 ;
        RECT 4.140 2.845 8.630 3.015 ;
        RECT 8.460 2.745 9.205 2.915 ;
        RECT 4.055 2.770 4.065 3.014 ;
        RECT 4.065 2.780 4.075 3.014 ;
        RECT 4.075 2.790 4.085 3.014 ;
        RECT 4.085 2.800 4.095 3.014 ;
        RECT 4.095 2.810 4.105 3.014 ;
        RECT 4.105 2.820 4.115 3.014 ;
        RECT 4.115 2.830 4.125 3.014 ;
        RECT 4.125 2.840 4.135 3.014 ;
        RECT 4.135 2.845 4.141 3.015 ;
        RECT 3.835 2.550 3.845 2.794 ;
        RECT 3.845 2.560 3.855 2.804 ;
        RECT 3.855 2.570 3.865 2.814 ;
        RECT 3.865 2.580 3.875 2.824 ;
        RECT 3.875 2.590 3.885 2.834 ;
        RECT 3.885 2.600 3.895 2.844 ;
        RECT 3.895 2.610 3.905 2.854 ;
        RECT 3.905 2.620 3.915 2.864 ;
        RECT 3.915 2.630 3.925 2.874 ;
        RECT 3.925 2.640 3.935 2.884 ;
        RECT 3.935 2.650 3.945 2.894 ;
        RECT 3.945 2.660 3.955 2.904 ;
        RECT 3.955 2.670 3.965 2.914 ;
        RECT 3.965 2.680 3.975 2.924 ;
        RECT 3.975 2.690 3.985 2.934 ;
        RECT 3.985 2.700 3.995 2.944 ;
        RECT 3.995 2.710 4.005 2.954 ;
        RECT 4.005 2.720 4.015 2.964 ;
        RECT 4.015 2.730 4.025 2.974 ;
        RECT 4.025 2.740 4.035 2.984 ;
        RECT 4.035 2.750 4.045 2.994 ;
        RECT 4.045 2.760 4.055 3.004 ;
        RECT 3.750 2.540 3.760 2.710 ;
        RECT 3.760 2.540 3.770 2.720 ;
        RECT 3.770 2.540 3.780 2.730 ;
        RECT 3.780 2.540 3.790 2.740 ;
        RECT 3.790 2.540 3.800 2.750 ;
        RECT 3.800 2.540 3.810 2.760 ;
        RECT 3.810 2.540 3.820 2.770 ;
        RECT 3.820 2.540 3.830 2.780 ;
        RECT 3.830 2.540 3.836 2.790 ;
        RECT 2.960 2.015 2.970 2.709 ;
        RECT 2.970 2.025 2.980 2.709 ;
        RECT 2.980 2.035 2.990 2.709 ;
        RECT 2.765 1.125 2.775 2.199 ;
        RECT 2.775 1.125 2.785 2.209 ;
        RECT 2.785 1.125 2.795 2.219 ;
        RECT 3.140 1.525 3.455 1.825 ;
        RECT 3.285 1.125 3.455 2.360 ;
        RECT 3.285 2.190 3.910 2.360 ;
        RECT 3.285 1.125 4.145 1.295 ;
        RECT 4.690 0.535 4.860 2.635 ;
        RECT 4.690 0.535 5.485 0.705 ;
        RECT 8.105 2.395 8.275 2.635 ;
        RECT 4.270 2.465 8.275 2.635 ;
        RECT 8.825 1.330 8.995 2.565 ;
        RECT 8.825 1.330 9.125 1.500 ;
        RECT 8.105 2.395 9.720 2.565 ;
        RECT 9.550 2.395 9.720 2.695 ;
        RECT 4.185 2.390 4.195 2.634 ;
        RECT 4.195 2.400 4.205 2.634 ;
        RECT 4.205 2.410 4.215 2.634 ;
        RECT 4.215 2.420 4.225 2.634 ;
        RECT 4.225 2.430 4.235 2.634 ;
        RECT 4.235 2.440 4.245 2.634 ;
        RECT 4.245 2.450 4.255 2.634 ;
        RECT 4.255 2.460 4.265 2.634 ;
        RECT 4.265 2.465 4.271 2.635 ;
        RECT 4.065 2.270 4.075 2.514 ;
        RECT 4.075 2.280 4.085 2.524 ;
        RECT 4.085 2.290 4.095 2.534 ;
        RECT 4.095 2.300 4.105 2.544 ;
        RECT 4.105 2.310 4.115 2.554 ;
        RECT 4.115 2.320 4.125 2.564 ;
        RECT 4.125 2.330 4.135 2.574 ;
        RECT 4.135 2.340 4.145 2.584 ;
        RECT 4.145 2.350 4.155 2.594 ;
        RECT 4.155 2.360 4.165 2.604 ;
        RECT 4.165 2.370 4.175 2.614 ;
        RECT 4.175 2.380 4.185 2.624 ;
        RECT 3.910 2.190 3.920 2.360 ;
        RECT 3.920 2.190 3.930 2.370 ;
        RECT 3.930 2.190 3.940 2.380 ;
        RECT 3.940 2.190 3.950 2.390 ;
        RECT 3.950 2.190 3.960 2.400 ;
        RECT 3.960 2.190 3.970 2.410 ;
        RECT 3.970 2.190 3.980 2.420 ;
        RECT 3.980 2.190 3.990 2.430 ;
        RECT 3.990 2.190 4.000 2.440 ;
        RECT 4.000 2.190 4.010 2.450 ;
        RECT 4.010 2.190 4.020 2.460 ;
        RECT 4.020 2.190 4.030 2.470 ;
        RECT 4.030 2.190 4.040 2.480 ;
        RECT 4.040 2.190 4.050 2.490 ;
        RECT 4.050 2.190 4.060 2.500 ;
        RECT 4.060 2.190 4.066 2.510 ;
        RECT 7.065 1.585 7.810 1.755 ;
        RECT 7.640 1.125 7.810 2.280 ;
        RECT 8.475 0.605 8.645 1.295 ;
        RECT 7.615 1.125 8.645 1.295 ;
        RECT 9.690 0.605 9.860 0.945 ;
        RECT 8.475 0.605 9.860 0.775 ;
        RECT 9.690 0.775 11.335 0.945 ;
        RECT 11.165 0.775 11.335 1.515 ;
        RECT 9.805 1.325 10.985 1.495 ;
        RECT 10.615 1.125 10.915 1.495 ;
        RECT 10.815 1.325 10.985 1.865 ;
        RECT 11.150 1.695 11.320 2.280 ;
        RECT 11.600 1.675 11.900 1.865 ;
        RECT 10.815 1.695 11.900 1.865 ;
        RECT 9.115 0.955 9.475 1.125 ;
        RECT 9.305 0.955 9.475 2.215 ;
        RECT 9.220 2.045 9.520 2.215 ;
        RECT 9.305 1.675 10.635 1.845 ;
        RECT 10.465 1.675 10.635 2.630 ;
        RECT 12.430 1.610 12.600 2.630 ;
        RECT 10.465 2.460 12.600 2.630 ;
  END 
END FFSDNRHDMXHT

MACRO FFSDNRHD2XHT
  CLASS  CORE ;
  FOREIGN FFSDNRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.940 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 3.650 1.525 4.140 2.010 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.080 0.720 13.250 2.960 ;
        RECT 13.080 1.650 13.430 2.015 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.990 0.720 12.210 1.600 ;
        RECT 12.005 0.720 12.210 2.280 ;
        RECT 11.990 1.980 12.210 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.460 0.410 3.180 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.900 1.605 8.510 1.775 ;
        RECT 8.300 1.605 8.510 2.055 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.470 1.325 1.555 1.845 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.415 -0.300 2.715 0.595 ;
        RECT 3.365 -0.300 3.665 0.595 ;
        RECT 5.935 -0.300 6.235 1.055 ;
        RECT 7.005 -0.300 7.305 0.595 ;
        RECT 8.110 -0.300 8.410 0.715 ;
        RECT 10.010 -0.300 10.310 0.595 ;
        RECT 11.520 -0.300 11.690 1.120 ;
        RECT 12.495 -0.300 12.795 1.055 ;
        RECT 13.535 -0.300 13.835 1.055 ;
        RECT 0.000 -0.300 13.940 0.300 ;
    END
  END GND
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.105 1.270 2.600 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.610 2.650 0.780 3.990 ;
        RECT 2.425 2.945 2.725 3.990 ;
        RECT 3.310 2.890 3.480 3.990 ;
        RECT 5.935 3.095 6.235 3.990 ;
        RECT 8.085 3.095 8.385 3.990 ;
        RECT 10.110 2.975 10.410 3.990 ;
        RECT 11.455 2.975 11.755 3.990 ;
        RECT 12.495 2.975 12.795 3.990 ;
        RECT 13.535 2.295 13.835 3.990 ;
        RECT 0.000 3.390 13.940 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 0.275 2.215 ;
        RECT 0.105 2.045 1.240 2.215 ;
        RECT 1.050 0.480 1.220 1.145 ;
        RECT 0.105 0.975 1.220 1.145 ;
        RECT 1.070 2.045 1.240 3.135 ;
        RECT 1.050 0.480 1.555 0.650 ;
        RECT 1.070 2.965 1.985 3.135 ;
        RECT 1.530 2.045 1.700 2.620 ;
        RECT 1.750 0.775 1.925 1.080 ;
        RECT 1.465 0.910 1.925 1.080 ;
        RECT 1.755 0.775 1.925 2.215 ;
        RECT 1.465 2.045 1.925 2.215 ;
        RECT 1.750 0.775 4.540 0.945 ;
        RECT 4.370 0.775 4.540 2.280 ;
        RECT 5.070 0.910 5.240 2.280 ;
        RECT 6.145 1.675 6.445 1.865 ;
        RECT 5.070 1.695 6.445 1.865 ;
        RECT 5.665 1.325 5.965 1.515 ;
        RECT 5.665 1.325 6.795 1.495 ;
        RECT 6.520 0.775 6.690 1.495 ;
        RECT 6.625 1.325 6.795 2.215 ;
        RECT 6.625 2.045 7.275 2.215 ;
        RECT 7.485 0.480 7.655 0.945 ;
        RECT 6.520 0.775 7.655 0.945 ;
        RECT 2.795 1.980 3.050 2.280 ;
        RECT 2.795 1.125 2.990 2.280 ;
        RECT 2.880 1.980 3.050 2.710 ;
        RECT 2.795 1.125 3.115 1.295 ;
        RECT 2.880 2.540 3.840 2.710 ;
        RECT 3.670 2.540 3.840 3.050 ;
        RECT 3.670 2.880 5.550 3.050 ;
        RECT 5.805 2.745 8.980 2.915 ;
        RECT 8.810 2.745 8.980 3.210 ;
        RECT 8.810 3.040 9.640 3.210 ;
        RECT 5.685 2.745 5.695 3.025 ;
        RECT 5.695 2.745 5.705 3.015 ;
        RECT 5.705 2.745 5.715 3.005 ;
        RECT 5.715 2.745 5.725 2.995 ;
        RECT 5.725 2.745 5.735 2.985 ;
        RECT 5.735 2.745 5.745 2.975 ;
        RECT 5.745 2.745 5.755 2.965 ;
        RECT 5.755 2.745 5.765 2.955 ;
        RECT 5.765 2.745 5.775 2.945 ;
        RECT 5.775 2.745 5.785 2.935 ;
        RECT 5.785 2.745 5.795 2.925 ;
        RECT 5.795 2.745 5.805 2.915 ;
        RECT 5.670 2.760 5.680 3.040 ;
        RECT 5.680 2.750 5.686 3.034 ;
        RECT 5.550 2.880 5.560 3.050 ;
        RECT 5.560 2.870 5.570 3.050 ;
        RECT 5.570 2.860 5.580 3.050 ;
        RECT 5.580 2.850 5.590 3.050 ;
        RECT 5.590 2.840 5.600 3.050 ;
        RECT 5.600 2.830 5.610 3.050 ;
        RECT 5.610 2.820 5.620 3.050 ;
        RECT 5.620 2.810 5.630 3.050 ;
        RECT 5.630 2.800 5.640 3.050 ;
        RECT 5.640 2.790 5.650 3.050 ;
        RECT 5.650 2.780 5.660 3.050 ;
        RECT 5.660 2.770 5.670 3.050 ;
        RECT 3.170 1.525 3.465 1.825 ;
        RECT 3.295 1.125 3.465 2.360 ;
        RECT 3.295 2.190 4.190 2.360 ;
        RECT 3.295 1.125 4.095 1.295 ;
        RECT 4.020 2.190 4.190 2.635 ;
        RECT 4.720 0.535 4.890 2.700 ;
        RECT 4.635 2.465 4.935 2.700 ;
        RECT 5.395 2.425 5.475 2.635 ;
        RECT 5.385 2.435 9.665 2.565 ;
        RECT 5.405 2.415 5.475 2.635 ;
        RECT 5.375 2.445 9.665 2.565 ;
        RECT 5.415 2.405 5.475 2.635 ;
        RECT 5.365 2.455 9.665 2.565 ;
        RECT 4.020 2.465 5.475 2.635 ;
        RECT 4.720 0.535 5.485 0.705 ;
        RECT 4.020 2.465 5.485 2.625 ;
        RECT 4.020 2.465 5.495 2.615 ;
        RECT 4.020 2.465 5.505 2.605 ;
        RECT 4.020 2.465 5.515 2.595 ;
        RECT 4.020 2.465 5.525 2.585 ;
        RECT 4.020 2.465 5.535 2.575 ;
        RECT 8.770 1.355 8.940 2.565 ;
        RECT 8.770 1.355 9.070 1.525 ;
        RECT 5.425 2.395 9.665 2.565 ;
        RECT 9.495 2.395 9.665 2.795 ;
        RECT 6.975 1.580 7.660 1.750 ;
        RECT 7.490 1.125 7.660 2.215 ;
        RECT 7.490 2.045 7.790 2.215 ;
        RECT 8.195 0.960 8.365 1.295 ;
        RECT 7.490 1.125 8.365 1.295 ;
        RECT 8.195 0.960 8.800 1.130 ;
        RECT 8.630 0.635 8.800 1.130 ;
        RECT 9.645 0.635 9.815 0.945 ;
        RECT 8.630 0.635 9.815 0.805 ;
        RECT 9.645 0.775 11.280 0.945 ;
        RECT 11.110 0.775 11.280 1.490 ;
        RECT 9.750 1.325 10.930 1.495 ;
        RECT 10.560 1.125 10.860 1.495 ;
        RECT 10.760 1.325 10.930 1.845 ;
        RECT 11.095 1.675 11.265 2.280 ;
        RECT 10.760 1.675 11.825 1.845 ;
        RECT 9.060 0.985 9.465 1.155 ;
        RECT 9.295 0.985 9.465 2.215 ;
        RECT 9.165 2.045 9.465 2.215 ;
        RECT 9.295 1.675 10.580 1.845 ;
        RECT 10.410 1.675 10.580 2.630 ;
        RECT 12.730 1.610 12.900 2.630 ;
        RECT 10.410 2.460 12.900 2.630 ;
  END 
END FFSDNRHD2XHT

MACRO FFSDNRHD1XHT
  CLASS  CORE ;
  FOREIGN FFSDNRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.120 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 3.650 1.525 4.140 2.010 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 12.780 0.720 13.020 1.360 ;
        RECT 12.810 0.720 13.020 2.960 ;
        RECT 12.780 1.980 13.020 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.580 0.720 11.910 1.470 ;
        RECT 11.580 1.300 12.250 1.470 ;
        RECT 12.080 1.300 12.250 2.275 ;
        RECT 11.675 2.105 12.250 2.275 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.460 0.410 3.180 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 8.030 1.610 8.510 2.010 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.470 1.325 1.555 1.845 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.415 -0.300 2.715 0.595 ;
        RECT 3.365 -0.300 3.665 0.595 ;
        RECT 5.980 -0.300 6.280 1.145 ;
        RECT 7.055 -0.300 7.355 0.590 ;
        RECT 8.125 -0.300 8.295 0.810 ;
        RECT 10.035 -0.300 10.335 0.525 ;
        RECT 11.195 -0.300 11.495 0.480 ;
        RECT 12.195 -0.300 12.495 1.055 ;
        RECT 0.000 -0.300 13.120 0.300 ;
    END
  END GND
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.105 1.270 2.600 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.610 2.880 0.780 3.990 ;
        RECT 2.425 2.880 2.725 3.990 ;
        RECT 3.310 2.890 3.480 3.990 ;
        RECT 6.035 3.195 6.335 3.990 ;
        RECT 8.165 3.195 8.465 3.990 ;
        RECT 10.165 2.975 10.465 3.990 ;
        RECT 12.195 2.975 12.495 3.990 ;
        RECT 0.000 3.390 13.120 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 0.275 2.215 ;
        RECT 0.105 2.045 1.225 2.215 ;
        RECT 1.055 2.045 1.225 3.185 ;
        RECT 1.085 0.480 1.255 1.145 ;
        RECT 0.105 0.975 1.255 1.145 ;
        RECT 1.085 0.480 1.555 0.650 ;
        RECT 1.055 3.015 1.985 3.185 ;
        RECT 1.530 2.045 1.700 2.620 ;
        RECT 1.750 0.775 1.925 1.120 ;
        RECT 1.465 0.950 1.925 1.120 ;
        RECT 1.755 0.775 1.925 2.215 ;
        RECT 1.465 2.045 1.925 2.215 ;
        RECT 1.750 0.775 4.540 0.945 ;
        RECT 4.370 0.775 4.540 2.280 ;
        RECT 5.070 0.900 5.240 2.280 ;
        RECT 6.235 1.675 6.535 1.865 ;
        RECT 5.070 1.695 6.535 1.865 ;
        RECT 5.715 1.325 6.015 1.515 ;
        RECT 6.650 0.775 6.885 1.495 ;
        RECT 5.715 1.325 6.885 1.495 ;
        RECT 6.715 0.775 6.885 2.215 ;
        RECT 6.715 2.045 7.255 2.215 ;
        RECT 7.540 0.480 7.710 0.945 ;
        RECT 6.650 0.775 7.710 0.945 ;
        RECT 2.795 1.980 3.050 2.280 ;
        RECT 2.795 1.125 2.990 2.280 ;
        RECT 2.880 1.980 3.050 2.710 ;
        RECT 2.795 1.125 3.115 1.295 ;
        RECT 2.880 2.540 3.840 2.710 ;
        RECT 3.670 2.540 3.840 3.015 ;
        RECT 8.460 2.745 8.630 3.015 ;
        RECT 3.670 2.845 8.630 3.015 ;
        RECT 8.460 2.745 9.205 2.915 ;
        RECT 3.170 1.525 3.465 1.825 ;
        RECT 3.295 1.125 3.465 2.360 ;
        RECT 3.295 2.190 4.190 2.360 ;
        RECT 3.295 1.125 4.095 1.295 ;
        RECT 4.020 2.190 4.190 2.665 ;
        RECT 4.720 0.535 4.890 2.665 ;
        RECT 4.720 0.535 5.515 0.705 ;
        RECT 8.105 2.395 8.275 2.665 ;
        RECT 4.020 2.495 8.275 2.665 ;
        RECT 8.825 1.330 8.995 2.565 ;
        RECT 8.825 1.330 9.125 1.500 ;
        RECT 8.105 2.395 9.720 2.565 ;
        RECT 9.550 2.395 9.720 2.795 ;
        RECT 7.065 1.585 7.810 1.755 ;
        RECT 7.640 1.125 7.810 2.280 ;
        RECT 8.475 0.605 8.645 1.295 ;
        RECT 7.615 1.125 8.645 1.295 ;
        RECT 9.690 0.605 9.860 0.945 ;
        RECT 8.475 0.605 9.860 0.775 ;
        RECT 9.690 0.775 11.335 0.945 ;
        RECT 11.165 0.775 11.335 1.575 ;
        RECT 10.615 1.125 10.985 1.495 ;
        RECT 9.855 1.325 10.985 1.495 ;
        RECT 10.815 1.125 10.985 1.925 ;
        RECT 11.150 1.755 11.320 2.280 ;
        RECT 11.600 1.675 11.900 1.925 ;
        RECT 10.815 1.755 11.900 1.925 ;
        RECT 9.115 0.955 9.475 1.125 ;
        RECT 9.305 0.955 9.475 2.215 ;
        RECT 9.220 2.045 9.520 2.215 ;
        RECT 9.305 1.675 10.635 1.845 ;
        RECT 10.465 1.675 10.635 2.630 ;
        RECT 12.430 1.610 12.600 2.630 ;
        RECT 10.465 2.460 12.600 2.630 ;
  END 
END FFSDNRHD1XHT

MACRO FFSDNHDMXHT
  CLASS  CORE ;
  FOREIGN FFSDNHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.070 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 3.635 1.525 4.110 2.010 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.730 1.060 10.970 1.360 ;
        RECT 10.760 1.060 10.970 2.280 ;
        RECT 10.730 1.980 10.970 2.280 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.690 1.060 9.860 1.470 ;
        RECT 9.690 1.290 10.150 1.470 ;
        RECT 9.940 1.290 10.150 2.215 ;
        RECT 9.625 2.045 10.150 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.415 -0.300 2.715 0.595 ;
        RECT 3.335 -0.300 3.635 0.595 ;
        RECT 5.815 -0.300 6.115 0.595 ;
        RECT 6.755 -0.300 7.055 0.595 ;
        RECT 8.655 -0.300 8.955 0.560 ;
        RECT 10.145 -0.300 10.445 0.595 ;
        RECT 0.000 -0.300 11.070 0.300 ;
    END
  END GND
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.265 2.680 2.565 3.990 ;
        RECT 3.265 2.890 3.565 3.990 ;
        RECT 5.925 3.160 6.225 3.990 ;
        RECT 6.755 3.160 7.055 3.990 ;
        RECT 8.600 2.745 8.770 3.990 ;
        RECT 10.145 2.925 10.445 3.990 ;
        RECT 0.000 3.390 11.070 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.555 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.150 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.980 0.775 2.150 1.035 ;
        RECT 1.530 0.865 2.150 1.035 ;
        RECT 1.980 0.775 4.510 0.945 ;
        RECT 4.340 0.480 4.510 2.280 ;
        RECT 5.040 0.900 5.210 2.280 ;
        RECT 6.185 1.675 6.495 1.865 ;
        RECT 5.040 1.695 6.495 1.865 ;
        RECT 5.685 1.325 5.985 1.515 ;
        RECT 6.430 0.900 6.600 1.495 ;
        RECT 5.685 1.325 7.165 1.495 ;
        RECT 6.995 1.325 7.165 2.215 ;
        RECT 6.365 2.045 7.165 2.215 ;
        RECT 2.765 1.125 2.960 2.710 ;
        RECT 2.765 1.125 3.105 1.295 ;
        RECT 2.765 2.540 3.715 2.710 ;
        RECT 4.075 2.810 7.635 2.980 ;
        RECT 3.985 2.730 3.995 2.980 ;
        RECT 3.995 2.740 4.005 2.980 ;
        RECT 4.005 2.750 4.015 2.980 ;
        RECT 4.015 2.760 4.025 2.980 ;
        RECT 4.025 2.770 4.035 2.980 ;
        RECT 4.035 2.780 4.045 2.980 ;
        RECT 4.045 2.790 4.055 2.980 ;
        RECT 4.055 2.800 4.065 2.980 ;
        RECT 4.065 2.810 4.075 2.980 ;
        RECT 3.805 2.550 3.815 2.800 ;
        RECT 3.815 2.560 3.825 2.810 ;
        RECT 3.825 2.570 3.835 2.820 ;
        RECT 3.835 2.580 3.845 2.830 ;
        RECT 3.845 2.590 3.855 2.840 ;
        RECT 3.855 2.600 3.865 2.850 ;
        RECT 3.865 2.610 3.875 2.860 ;
        RECT 3.875 2.620 3.885 2.870 ;
        RECT 3.885 2.630 3.895 2.880 ;
        RECT 3.895 2.640 3.905 2.890 ;
        RECT 3.905 2.650 3.915 2.900 ;
        RECT 3.915 2.660 3.925 2.910 ;
        RECT 3.925 2.670 3.935 2.920 ;
        RECT 3.935 2.680 3.945 2.930 ;
        RECT 3.945 2.690 3.955 2.940 ;
        RECT 3.955 2.700 3.965 2.950 ;
        RECT 3.965 2.710 3.975 2.960 ;
        RECT 3.975 2.720 3.985 2.970 ;
        RECT 3.715 2.540 3.725 2.710 ;
        RECT 3.725 2.540 3.735 2.720 ;
        RECT 3.735 2.540 3.745 2.730 ;
        RECT 3.745 2.540 3.755 2.740 ;
        RECT 3.755 2.540 3.765 2.750 ;
        RECT 3.765 2.540 3.775 2.760 ;
        RECT 3.775 2.540 3.785 2.770 ;
        RECT 3.785 2.540 3.795 2.780 ;
        RECT 3.795 2.540 3.805 2.790 ;
        RECT 3.170 1.525 3.455 1.825 ;
        RECT 3.285 1.125 3.455 2.360 ;
        RECT 3.265 1.525 3.455 2.360 ;
        RECT 3.265 2.190 3.905 2.360 ;
        RECT 3.285 1.125 4.145 1.295 ;
        RECT 4.690 0.535 4.860 2.630 ;
        RECT 4.690 0.535 5.485 0.705 ;
        RECT 7.345 0.500 7.515 2.630 ;
        RECT 7.345 0.500 7.745 0.670 ;
        RECT 7.345 2.440 8.150 2.630 ;
        RECT 4.260 2.460 8.150 2.630 ;
        RECT 7.980 2.440 8.150 2.770 ;
        RECT 4.175 2.385 4.185 2.629 ;
        RECT 4.185 2.395 4.195 2.629 ;
        RECT 4.195 2.405 4.205 2.629 ;
        RECT 4.205 2.415 4.215 2.629 ;
        RECT 4.215 2.425 4.225 2.629 ;
        RECT 4.225 2.435 4.235 2.629 ;
        RECT 4.235 2.445 4.245 2.629 ;
        RECT 4.245 2.455 4.255 2.629 ;
        RECT 4.255 2.460 4.261 2.630 ;
        RECT 4.065 2.275 4.075 2.519 ;
        RECT 4.075 2.285 4.085 2.529 ;
        RECT 4.085 2.295 4.095 2.539 ;
        RECT 4.095 2.305 4.105 2.549 ;
        RECT 4.105 2.315 4.115 2.559 ;
        RECT 4.115 2.325 4.125 2.569 ;
        RECT 4.125 2.335 4.135 2.579 ;
        RECT 4.135 2.345 4.145 2.589 ;
        RECT 4.145 2.355 4.155 2.599 ;
        RECT 4.155 2.365 4.165 2.609 ;
        RECT 4.165 2.375 4.175 2.619 ;
        RECT 3.905 2.190 3.915 2.360 ;
        RECT 3.915 2.190 3.925 2.370 ;
        RECT 3.925 2.190 3.935 2.380 ;
        RECT 3.935 2.190 3.945 2.390 ;
        RECT 3.945 2.190 3.955 2.400 ;
        RECT 3.955 2.190 3.965 2.410 ;
        RECT 3.965 2.190 3.975 2.420 ;
        RECT 3.975 2.190 3.985 2.430 ;
        RECT 3.985 2.190 3.995 2.440 ;
        RECT 3.995 2.190 4.005 2.450 ;
        RECT 4.005 2.190 4.015 2.460 ;
        RECT 4.015 2.190 4.025 2.470 ;
        RECT 4.025 2.190 4.035 2.480 ;
        RECT 4.035 2.190 4.045 2.490 ;
        RECT 4.045 2.190 4.055 2.500 ;
        RECT 4.055 2.190 4.065 2.510 ;
        RECT 8.405 1.310 9.385 1.480 ;
        RECT 9.180 0.875 9.350 1.480 ;
        RECT 9.215 1.310 9.385 2.215 ;
        RECT 9.085 2.045 9.385 2.215 ;
        RECT 9.215 1.650 9.735 1.820 ;
        RECT 7.770 0.875 7.940 2.215 ;
        RECT 7.695 2.045 8.905 2.215 ;
        RECT 8.735 2.045 8.905 2.565 ;
        RECT 8.970 2.395 9.140 2.780 ;
        RECT 10.380 1.520 10.550 2.565 ;
        RECT 8.735 2.395 10.550 2.565 ;
        RECT 10.380 1.520 10.570 1.820 ;
  END 
END FFSDNHDMXHT

MACRO FFSDNHDLXHT
  CLASS  CORE ;
  FOREIGN FFSDNHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.070 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 3.670 1.525 4.160 2.010 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.730 1.060 10.970 1.360 ;
        RECT 10.760 1.060 10.970 2.280 ;
        RECT 10.730 1.980 10.970 2.280 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.750 1.060 9.920 1.470 ;
        RECT 9.750 1.290 10.150 1.470 ;
        RECT 9.940 1.290 10.150 2.215 ;
        RECT 9.685 2.045 10.150 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.110 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.435 -0.300 2.735 0.595 ;
        RECT 3.385 -0.300 3.685 0.595 ;
        RECT 5.875 -0.300 6.175 0.595 ;
        RECT 6.815 -0.300 7.115 0.565 ;
        RECT 8.715 -0.300 9.015 0.560 ;
        RECT 10.115 -0.300 10.415 0.745 ;
        RECT 0.000 -0.300 11.070 0.300 ;
    END
  END GND
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.385 2.575 2.685 3.990 ;
        RECT 3.310 2.890 3.480 3.990 ;
        RECT 6.055 3.160 7.035 3.990 ;
        RECT 8.660 2.745 8.830 3.990 ;
        RECT 10.115 2.745 10.415 3.990 ;
        RECT 0.000 3.390 11.070 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.500 1.350 2.630 ;
        RECT 1.180 0.500 1.555 0.670 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.010 ;
        RECT 1.530 0.885 1.700 2.280 ;
        RECT 1.530 0.885 1.720 1.210 ;
        RECT 2.010 0.775 2.180 1.055 ;
        RECT 1.530 0.885 2.180 1.055 ;
        RECT 2.010 0.775 4.530 0.945 ;
        RECT 4.295 0.505 4.530 0.945 ;
        RECT 4.370 1.890 4.570 1.949 ;
        RECT 4.380 1.890 4.570 1.959 ;
        RECT 4.390 1.890 4.570 1.969 ;
        RECT 4.360 0.505 4.530 1.939 ;
        RECT 4.360 1.860 4.540 1.939 ;
        RECT 4.360 1.870 4.550 1.939 ;
        RECT 4.360 1.880 4.560 1.939 ;
        RECT 4.400 1.890 4.570 2.280 ;
        RECT 5.080 0.900 5.250 1.554 ;
        RECT 5.090 1.475 5.270 1.564 ;
        RECT 5.100 0.900 5.250 2.280 ;
        RECT 5.080 1.465 5.260 1.554 ;
        RECT 5.100 1.475 5.270 2.279 ;
        RECT 6.215 1.675 6.515 1.865 ;
        RECT 5.100 1.695 6.515 1.865 ;
        RECT 5.725 1.325 6.025 1.515 ;
        RECT 6.490 0.900 6.660 1.495 ;
        RECT 5.725 1.325 7.225 1.495 ;
        RECT 7.055 1.325 7.225 2.215 ;
        RECT 6.415 2.045 7.225 2.215 ;
        RECT 2.805 1.985 3.070 2.285 ;
        RECT 2.805 1.125 2.975 2.285 ;
        RECT 2.900 1.985 3.070 2.710 ;
        RECT 2.805 1.125 3.125 1.295 ;
        RECT 2.900 2.540 3.870 2.710 ;
        RECT 3.700 2.540 3.870 2.980 ;
        RECT 3.700 2.810 7.685 2.980 ;
        RECT 3.190 1.525 3.485 1.825 ;
        RECT 3.315 1.125 3.485 2.360 ;
        RECT 3.315 2.190 4.220 2.360 ;
        RECT 3.315 1.125 4.165 1.295 ;
        RECT 4.050 2.190 4.220 2.630 ;
        RECT 4.720 1.710 4.920 1.769 ;
        RECT 4.730 1.710 4.920 1.779 ;
        RECT 4.740 1.710 4.920 1.789 ;
        RECT 4.710 0.535 4.880 1.759 ;
        RECT 4.710 1.680 4.890 1.759 ;
        RECT 4.710 1.690 4.900 1.759 ;
        RECT 4.710 1.700 4.910 1.759 ;
        RECT 4.750 1.710 4.920 2.630 ;
        RECT 4.710 0.535 5.525 0.705 ;
        RECT 7.405 0.500 7.575 2.630 ;
        RECT 7.405 0.500 7.805 0.670 ;
        RECT 4.050 2.460 8.275 2.630 ;
        RECT 8.465 1.400 9.455 1.570 ;
        RECT 9.240 0.875 9.410 1.570 ;
        RECT 9.285 1.400 9.455 2.215 ;
        RECT 9.145 2.045 9.455 2.215 ;
        RECT 9.285 1.650 9.760 1.820 ;
        RECT 7.830 0.875 8.000 2.215 ;
        RECT 7.755 2.045 8.965 2.215 ;
        RECT 8.795 2.045 8.965 2.565 ;
        RECT 9.030 2.395 9.200 2.770 ;
        RECT 10.380 1.520 10.550 2.565 ;
        RECT 8.795 2.395 10.550 2.565 ;
        RECT 10.380 1.520 10.580 1.820 ;
  END 
END FFSDNHDLXHT

MACRO FFSDNHD2XHT
  CLASS  CORE ;
  FOREIGN FFSDNHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.300 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 3.650 1.525 4.140 2.010 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.440 0.720 11.610 2.960 ;
        RECT 11.440 1.640 11.790 2.015 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.350 0.720 10.570 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.460 0.410 3.180 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.470 1.325 1.555 1.845 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.415 -0.300 2.715 0.595 ;
        RECT 3.365 -0.300 3.665 0.595 ;
        RECT 5.805 -0.300 6.105 0.595 ;
        RECT 6.820 -0.300 7.120 0.715 ;
        RECT 8.565 -0.300 8.735 0.780 ;
        RECT 9.920 -0.300 10.090 1.190 ;
        RECT 9.880 0.890 10.090 1.190 ;
        RECT 10.855 -0.300 11.155 1.055 ;
        RECT 11.895 -0.300 12.195 1.055 ;
        RECT 0.000 -0.300 12.300 0.300 ;
    END
  END GND
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.270 2.600 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.610 2.650 0.780 3.990 ;
        RECT 2.415 2.945 2.715 3.990 ;
        RECT 3.310 2.890 3.480 3.990 ;
        RECT 5.950 3.160 6.250 3.990 ;
        RECT 6.790 3.095 7.090 3.990 ;
        RECT 8.685 2.805 8.855 3.990 ;
        RECT 9.815 2.975 10.115 3.990 ;
        RECT 10.855 2.975 11.155 3.990 ;
        RECT 11.895 2.295 12.195 3.990 ;
        RECT 0.000 3.390 12.300 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 0.275 2.215 ;
        RECT 0.105 2.045 1.245 2.215 ;
        RECT 1.075 2.045 1.245 3.105 ;
        RECT 1.085 0.480 1.255 1.145 ;
        RECT 0.105 0.975 1.255 1.145 ;
        RECT 1.085 0.480 1.555 0.650 ;
        RECT 1.075 2.935 2.025 3.105 ;
        RECT 1.530 2.045 1.700 2.620 ;
        RECT 1.750 0.775 1.925 1.120 ;
        RECT 1.465 0.950 1.925 1.120 ;
        RECT 1.755 0.775 1.925 2.215 ;
        RECT 1.465 2.045 1.925 2.215 ;
        RECT 1.750 0.775 4.540 0.945 ;
        RECT 4.370 0.775 4.540 2.280 ;
        RECT 5.070 0.910 5.240 2.280 ;
        RECT 6.175 1.675 6.475 1.865 ;
        RECT 5.070 1.695 6.475 1.865 ;
        RECT 5.665 1.325 5.965 1.515 ;
        RECT 6.420 0.910 6.590 1.495 ;
        RECT 5.665 1.325 7.210 1.495 ;
        RECT 7.040 1.325 7.210 2.215 ;
        RECT 6.390 2.045 7.210 2.215 ;
        RECT 2.795 1.980 3.050 2.280 ;
        RECT 2.795 1.125 2.990 2.280 ;
        RECT 2.880 1.980 3.050 2.710 ;
        RECT 2.795 1.125 3.115 1.295 ;
        RECT 2.880 2.540 3.840 2.710 ;
        RECT 3.670 2.540 3.840 3.035 ;
        RECT 3.670 2.865 5.565 3.035 ;
        RECT 5.805 2.745 7.475 2.915 ;
        RECT 7.305 2.745 7.475 3.210 ;
        RECT 7.305 3.040 8.290 3.210 ;
        RECT 5.685 2.745 5.695 3.025 ;
        RECT 5.695 2.745 5.705 3.015 ;
        RECT 5.705 2.745 5.715 3.005 ;
        RECT 5.715 2.745 5.725 2.995 ;
        RECT 5.725 2.745 5.735 2.985 ;
        RECT 5.735 2.745 5.745 2.975 ;
        RECT 5.745 2.745 5.755 2.965 ;
        RECT 5.755 2.745 5.765 2.955 ;
        RECT 5.765 2.745 5.775 2.945 ;
        RECT 5.775 2.745 5.785 2.935 ;
        RECT 5.785 2.745 5.795 2.925 ;
        RECT 5.795 2.745 5.805 2.915 ;
        RECT 5.565 2.865 5.575 3.035 ;
        RECT 5.575 2.855 5.585 3.035 ;
        RECT 5.585 2.845 5.595 3.035 ;
        RECT 5.595 2.835 5.605 3.035 ;
        RECT 5.605 2.825 5.615 3.035 ;
        RECT 5.615 2.815 5.625 3.035 ;
        RECT 5.625 2.805 5.635 3.035 ;
        RECT 5.635 2.795 5.645 3.035 ;
        RECT 5.645 2.785 5.655 3.035 ;
        RECT 5.655 2.775 5.665 3.035 ;
        RECT 5.665 2.765 5.675 3.035 ;
        RECT 5.675 2.755 5.685 3.035 ;
        RECT 3.170 1.525 3.465 1.825 ;
        RECT 3.295 1.125 3.465 2.360 ;
        RECT 3.295 2.190 4.190 2.360 ;
        RECT 3.295 1.125 4.095 1.295 ;
        RECT 4.020 2.190 4.190 2.685 ;
        RECT 4.720 0.535 4.890 2.685 ;
        RECT 4.020 2.515 5.305 2.685 ;
        RECT 4.720 0.535 5.485 0.705 ;
        RECT 7.390 0.710 7.560 2.565 ;
        RECT 5.545 2.395 7.575 2.565 ;
        RECT 7.635 2.395 7.650 2.625 ;
        RECT 7.710 2.455 8.225 2.625 ;
        RECT 7.390 0.710 8.330 0.880 ;
        RECT 8.055 2.455 8.225 2.795 ;
        RECT 8.160 0.710 8.330 1.140 ;
        RECT 8.915 0.480 9.085 1.140 ;
        RECT 8.160 0.970 9.085 1.140 ;
        RECT 8.915 0.480 9.740 0.650 ;
        RECT 7.650 2.405 7.660 2.625 ;
        RECT 7.660 2.415 7.670 2.625 ;
        RECT 7.670 2.425 7.680 2.625 ;
        RECT 7.680 2.435 7.690 2.625 ;
        RECT 7.690 2.445 7.700 2.625 ;
        RECT 7.700 2.455 7.710 2.625 ;
        RECT 7.575 2.395 7.585 2.565 ;
        RECT 7.585 2.395 7.595 2.575 ;
        RECT 7.595 2.395 7.605 2.585 ;
        RECT 7.605 2.395 7.615 2.595 ;
        RECT 7.615 2.395 7.625 2.605 ;
        RECT 7.625 2.395 7.635 2.615 ;
        RECT 5.425 2.395 5.435 2.675 ;
        RECT 5.435 2.395 5.445 2.665 ;
        RECT 5.445 2.395 5.455 2.655 ;
        RECT 5.455 2.395 5.465 2.645 ;
        RECT 5.465 2.395 5.475 2.635 ;
        RECT 5.475 2.395 5.485 2.625 ;
        RECT 5.485 2.395 5.495 2.615 ;
        RECT 5.495 2.395 5.505 2.605 ;
        RECT 5.505 2.395 5.515 2.595 ;
        RECT 5.515 2.395 5.525 2.585 ;
        RECT 5.525 2.395 5.535 2.575 ;
        RECT 5.535 2.395 5.545 2.565 ;
        RECT 5.305 2.515 5.315 2.685 ;
        RECT 5.315 2.505 5.325 2.685 ;
        RECT 5.325 2.495 5.335 2.685 ;
        RECT 5.335 2.485 5.345 2.685 ;
        RECT 5.345 2.475 5.355 2.685 ;
        RECT 5.355 2.465 5.365 2.685 ;
        RECT 5.365 2.455 5.375 2.685 ;
        RECT 5.375 2.445 5.385 2.685 ;
        RECT 5.385 2.435 5.395 2.685 ;
        RECT 5.395 2.425 5.405 2.685 ;
        RECT 5.405 2.415 5.415 2.685 ;
        RECT 5.415 2.405 5.425 2.685 ;
        RECT 9.265 1.060 9.435 2.280 ;
        RECT 8.480 1.675 10.170 1.845 ;
        RECT 7.805 1.060 7.975 2.230 ;
        RECT 7.740 2.060 9.085 2.230 ;
        RECT 8.915 2.060 9.085 2.630 ;
        RECT 9.055 2.460 9.225 3.190 ;
        RECT 11.090 1.610 11.260 2.630 ;
        RECT 8.915 2.460 11.260 2.630 ;
  END 
END FFSDNHD2XHT

MACRO FFSDNHD1XHT
  CLASS  CORE ;
  FOREIGN FFSDNHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.070 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 3.650 1.525 4.140 2.010 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.730 0.720 10.970 1.360 ;
        RECT 10.760 0.720 10.970 2.960 ;
        RECT 10.730 1.980 10.970 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.690 0.720 9.860 1.470 ;
        RECT 9.690 1.290 10.150 1.470 ;
        RECT 9.940 1.290 10.150 2.215 ;
        RECT 9.625 2.045 10.150 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.460 0.410 3.180 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.470 1.325 1.555 1.845 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.415 -0.300 2.715 0.595 ;
        RECT 3.365 -0.300 3.665 0.595 ;
        RECT 5.845 -0.300 6.145 0.595 ;
        RECT 6.785 -0.300 7.085 0.565 ;
        RECT 8.675 -0.300 8.975 0.630 ;
        RECT 10.145 -0.300 10.445 1.055 ;
        RECT 0.000 -0.300 11.070 0.300 ;
    END
  END GND
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.105 1.270 2.600 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.610 2.880 0.780 3.990 ;
        RECT 2.395 2.580 2.695 3.990 ;
        RECT 3.310 2.890 3.480 3.990 ;
        RECT 6.025 3.160 7.005 3.990 ;
        RECT 8.600 2.745 8.770 3.990 ;
        RECT 10.145 2.975 10.445 3.990 ;
        RECT 0.000 3.390 11.070 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 0.275 2.215 ;
        RECT 0.105 2.045 1.250 2.215 ;
        RECT 1.080 2.045 1.250 3.210 ;
        RECT 1.085 0.480 1.255 1.145 ;
        RECT 0.105 0.975 1.255 1.145 ;
        RECT 1.085 0.480 1.555 0.650 ;
        RECT 1.080 3.040 1.985 3.210 ;
        RECT 1.540 2.045 1.710 2.620 ;
        RECT 1.750 0.775 1.925 1.120 ;
        RECT 1.465 0.950 1.925 1.120 ;
        RECT 1.755 0.775 1.925 2.215 ;
        RECT 1.475 2.045 1.925 2.215 ;
        RECT 1.750 0.775 4.540 0.945 ;
        RECT 4.370 0.775 4.540 2.280 ;
        RECT 5.070 0.900 5.240 2.280 ;
        RECT 6.215 1.675 6.525 1.865 ;
        RECT 5.070 1.695 6.525 1.865 ;
        RECT 5.715 1.325 6.015 1.515 ;
        RECT 6.460 0.910 6.630 1.495 ;
        RECT 5.715 1.325 7.195 1.495 ;
        RECT 7.025 1.325 7.195 2.215 ;
        RECT 6.395 2.045 7.195 2.215 ;
        RECT 2.810 1.980 3.050 2.280 ;
        RECT 2.810 1.125 2.990 2.280 ;
        RECT 2.880 1.980 3.050 2.710 ;
        RECT 2.810 1.125 3.115 1.295 ;
        RECT 2.880 2.540 3.840 2.710 ;
        RECT 3.670 2.540 3.840 2.980 ;
        RECT 3.670 2.810 7.775 2.980 ;
        RECT 3.170 1.525 3.465 1.825 ;
        RECT 3.295 1.125 3.465 2.360 ;
        RECT 3.295 2.190 4.190 2.360 ;
        RECT 3.295 1.125 4.095 1.295 ;
        RECT 4.020 2.190 4.190 2.630 ;
        RECT 4.720 0.535 4.890 2.630 ;
        RECT 4.720 0.535 5.515 0.705 ;
        RECT 7.375 0.500 7.545 2.630 ;
        RECT 7.375 0.500 7.775 0.670 ;
        RECT 7.375 2.440 8.220 2.630 ;
        RECT 4.020 2.460 8.220 2.630 ;
        RECT 8.050 2.440 8.220 2.995 ;
        RECT 8.415 1.400 9.390 1.570 ;
        RECT 9.180 0.945 9.350 1.570 ;
        RECT 9.220 1.400 9.390 2.215 ;
        RECT 9.085 2.045 9.390 2.215 ;
        RECT 9.220 1.650 9.735 1.820 ;
        RECT 7.790 0.945 7.960 2.215 ;
        RECT 7.725 2.045 8.905 2.215 ;
        RECT 8.735 2.045 8.905 2.565 ;
        RECT 8.970 2.395 9.140 2.780 ;
        RECT 10.380 1.520 10.550 2.565 ;
        RECT 8.735 2.395 10.550 2.565 ;
        RECT 10.380 1.520 10.570 1.820 ;
  END 
END FFSDNHD1XHT

MACRO FFSDHQHDMXHT
  CLASS  CORE ;
  FOREIGN FFSDHQHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.300 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.760 1.060 12.200 1.360 ;
        RECT 11.950 1.060 12.200 2.455 ;
        RECT 11.760 1.980 12.200 2.455 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.240 1.165 1.775 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.575 0.380 2.020 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.870 ;
        RECT 2.545 -0.300 2.845 0.595 ;
        RECT 3.525 -0.300 3.825 0.595 ;
        RECT 4.495 -0.300 4.795 0.595 ;
        RECT 7.350 -0.300 7.650 0.595 ;
        RECT 8.430 -0.300 8.730 0.595 ;
        RECT 10.585 -0.300 10.755 0.805 ;
        RECT 11.185 -0.300 11.485 0.945 ;
        RECT 0.000 -0.300 12.300 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 4.495 1.560 5.010 2.020 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.365 1.530 2.805 2.020 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.655 0.955 3.990 ;
        RECT 2.555 2.470 2.730 3.990 ;
        RECT 3.555 2.745 3.855 3.990 ;
        RECT 4.460 2.745 4.760 3.990 ;
        RECT 7.410 2.885 7.710 3.990 ;
        RECT 8.465 2.885 8.765 3.990 ;
        RECT 10.415 2.610 10.585 3.990 ;
        RECT 11.250 2.650 11.420 3.990 ;
        RECT 0.000 3.390 12.300 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.075 0.730 1.245 ;
        RECT 0.560 1.075 0.730 2.405 ;
        RECT 0.105 2.235 0.730 2.405 ;
        RECT 1.355 1.510 1.525 2.125 ;
        RECT 0.560 1.955 1.525 2.125 ;
        RECT 1.355 1.510 1.630 1.810 ;
        RECT 3.390 1.605 3.560 1.905 ;
        RECT 3.390 1.605 4.285 1.775 ;
        RECT 3.985 1.125 4.285 2.215 ;
        RECT 5.080 1.125 5.735 1.295 ;
        RECT 5.565 1.125 5.735 2.215 ;
        RECT 5.350 2.045 5.735 2.215 ;
        RECT 1.640 1.070 1.980 1.260 ;
        RECT 1.640 0.960 1.810 1.260 ;
        RECT 1.640 2.330 1.810 2.970 ;
        RECT 1.810 1.070 1.980 2.515 ;
        RECT 1.640 2.330 1.980 2.515 ;
        RECT 2.485 0.775 2.655 1.240 ;
        RECT 1.640 1.070 2.655 1.240 ;
        RECT 2.485 0.775 6.095 0.945 ;
        RECT 5.925 0.775 6.095 2.320 ;
        RECT 6.625 1.060 6.795 2.320 ;
        RECT 7.690 1.585 7.860 2.210 ;
        RECT 6.625 2.040 7.860 2.210 ;
        RECT 7.690 1.585 8.070 1.755 ;
        RECT 7.335 1.125 7.505 1.820 ;
        RECT 8.050 1.970 8.220 2.280 ;
        RECT 7.335 1.125 8.695 1.295 ;
        RECT 8.525 1.125 8.695 2.140 ;
        RECT 8.050 1.970 8.695 2.140 ;
        RECT 3.005 1.125 3.185 2.565 ;
        RECT 3.005 2.105 3.240 2.565 ;
        RECT 3.005 1.125 3.305 1.370 ;
        RECT 5.170 2.395 5.470 2.670 ;
        RECT 3.005 2.395 5.470 2.565 ;
        RECT 6.275 0.650 6.445 2.670 ;
        RECT 5.170 2.500 6.445 2.670 ;
        RECT 6.975 0.650 7.145 0.945 ;
        RECT 6.275 0.650 7.145 0.820 ;
        RECT 6.975 0.775 9.045 0.945 ;
        RECT 8.875 0.775 9.045 1.610 ;
        RECT 8.875 1.310 9.440 1.610 ;
        RECT 8.945 1.925 9.115 2.705 ;
        RECT 6.740 2.535 9.115 2.705 ;
        RECT 9.655 0.985 9.825 2.095 ;
        RECT 8.945 1.925 9.825 2.095 ;
        RECT 9.655 0.985 9.945 1.285 ;
        RECT 10.005 1.550 10.175 2.605 ;
        RECT 9.385 2.435 10.175 2.605 ;
        RECT 9.420 0.570 10.365 0.740 ;
        RECT 10.195 0.570 10.365 1.720 ;
        RECT 10.005 1.550 11.190 1.720 ;
        RECT 10.380 1.925 10.550 2.295 ;
        RECT 10.635 1.125 11.560 1.295 ;
        RECT 11.370 1.125 11.560 2.295 ;
        RECT 10.380 2.125 11.560 2.295 ;
  END 
END FFSDHQHDMXHT

MACRO FFSDHQHD3XHT
  CLASS  CORE ;
  FOREIGN FFSDHQHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.760 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.285 0.480 13.455 1.130 ;
        RECT 13.285 2.400 13.455 3.040 ;
        RECT 13.285 0.960 14.670 1.130 ;
        RECT 13.285 2.400 14.670 2.625 ;
        RECT 14.325 0.720 14.670 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.240 1.165 1.775 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.545 0.380 2.020 ;
        RECT 0.225 0.755 0.525 0.945 ;
        RECT 1.215 0.485 1.385 0.945 ;
        RECT 0.225 0.775 1.385 0.945 ;
        RECT 1.215 0.485 2.155 0.655 ;
        RECT 0.300 2.580 0.485 2.820 ;
        RECT 0.185 2.650 0.485 2.820 ;
        RECT 0.300 2.580 1.340 2.750 ;
        RECT 0.185 2.650 1.340 2.750 ;
        RECT 1.170 2.580 1.340 3.190 ;
        RECT 1.170 3.020 2.245 3.190 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.595 ;
        RECT 2.550 -0.300 2.850 0.595 ;
        RECT 3.475 -0.300 3.775 0.595 ;
        RECT 4.430 -0.300 4.730 0.595 ;
        RECT 5.530 -0.300 5.830 0.595 ;
        RECT 7.490 -0.300 7.790 0.595 ;
        RECT 9.870 -0.300 10.170 0.665 ;
        RECT 11.990 -0.300 12.160 0.850 ;
        RECT 12.765 -0.300 12.935 0.780 ;
        RECT 13.805 -0.300 13.975 0.780 ;
        RECT 0.000 -0.300 14.760 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 4.535 1.570 5.080 2.020 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.530 2.505 2.020 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.975 0.955 3.990 ;
        RECT 2.560 2.830 2.730 3.990 ;
        RECT 3.670 2.830 3.840 3.990 ;
        RECT 4.420 2.850 4.720 3.990 ;
        RECT 7.465 2.910 7.635 3.990 ;
        RECT 9.840 2.975 10.140 3.990 ;
        RECT 11.695 2.400 11.995 3.990 ;
        RECT 12.765 2.910 12.935 3.990 ;
        RECT 13.805 2.910 13.975 3.990 ;
        RECT 0.000 3.390 14.760 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.100 1.125 0.730 1.295 ;
        RECT 0.560 1.125 0.730 2.400 ;
        RECT 0.105 2.230 0.730 2.400 ;
        RECT 1.345 1.460 1.515 2.160 ;
        RECT 0.560 1.990 1.515 2.160 ;
        RECT 1.345 1.460 1.965 1.760 ;
        RECT 3.430 1.605 3.600 1.905 ;
        RECT 3.430 1.605 4.325 1.780 ;
        RECT 4.025 1.125 4.325 2.215 ;
        RECT 4.980 1.125 5.775 1.295 ;
        RECT 5.605 1.125 5.775 2.370 ;
        RECT 5.350 2.200 5.775 2.370 ;
        RECT 1.575 2.330 1.875 2.840 ;
        RECT 1.575 1.070 2.855 1.250 ;
        RECT 2.685 0.775 2.855 2.500 ;
        RECT 1.575 2.330 2.855 2.500 ;
        RECT 2.685 0.775 6.155 0.945 ;
        RECT 5.985 0.775 6.155 2.720 ;
        RECT 6.685 1.060 6.855 2.400 ;
        RECT 7.815 1.520 7.985 2.210 ;
        RECT 6.685 2.040 7.985 2.210 ;
        RECT 7.815 1.520 8.070 1.820 ;
        RECT 7.395 1.170 7.565 1.820 ;
        RECT 8.045 1.125 8.420 1.340 ;
        RECT 7.395 1.170 8.420 1.340 ;
        RECT 8.165 2.065 8.335 2.705 ;
        RECT 8.250 1.125 8.420 2.235 ;
        RECT 8.165 2.065 8.420 2.235 ;
        RECT 8.250 1.550 10.145 1.720 ;
        RECT 3.045 1.125 3.225 2.680 ;
        RECT 3.045 2.040 3.280 2.680 ;
        RECT 3.045 1.125 3.345 1.295 ;
        RECT 3.045 2.440 5.095 2.610 ;
        RECT 4.925 2.440 5.095 3.135 ;
        RECT 4.925 2.870 5.470 3.135 ;
        RECT 6.335 0.555 6.505 3.135 ;
        RECT 4.925 2.965 6.505 3.135 ;
        RECT 6.335 0.555 7.195 0.725 ;
        RECT 7.025 0.555 7.195 0.945 ;
        RECT 7.025 0.775 8.575 0.945 ;
        RECT 8.890 0.980 9.155 1.150 ;
        RECT 8.985 0.980 9.155 1.365 ;
        RECT 8.985 1.195 10.815 1.365 ;
        RECT 10.645 1.195 10.815 1.680 ;
        RECT 8.780 0.880 8.790 1.150 ;
        RECT 8.790 0.890 8.800 1.150 ;
        RECT 8.800 0.900 8.810 1.150 ;
        RECT 8.810 0.910 8.820 1.150 ;
        RECT 8.820 0.920 8.830 1.150 ;
        RECT 8.830 0.930 8.840 1.150 ;
        RECT 8.840 0.940 8.850 1.150 ;
        RECT 8.850 0.950 8.860 1.150 ;
        RECT 8.860 0.960 8.870 1.150 ;
        RECT 8.870 0.970 8.880 1.150 ;
        RECT 8.880 0.980 8.890 1.150 ;
        RECT 8.770 0.870 8.780 1.140 ;
        RECT 8.600 0.525 8.610 0.969 ;
        RECT 8.610 0.525 8.620 0.979 ;
        RECT 8.620 0.525 8.630 0.989 ;
        RECT 8.630 0.525 8.640 0.999 ;
        RECT 8.640 0.525 8.650 1.009 ;
        RECT 8.650 0.525 8.660 1.019 ;
        RECT 8.660 0.525 8.670 1.029 ;
        RECT 8.670 0.525 8.680 1.039 ;
        RECT 8.680 0.525 8.690 1.049 ;
        RECT 8.690 0.525 8.700 1.059 ;
        RECT 8.700 0.525 8.710 1.069 ;
        RECT 8.710 0.525 8.720 1.079 ;
        RECT 8.720 0.525 8.730 1.089 ;
        RECT 8.730 0.525 8.740 1.099 ;
        RECT 8.740 0.525 8.750 1.109 ;
        RECT 8.750 0.525 8.760 1.119 ;
        RECT 8.760 0.525 8.770 1.129 ;
        RECT 8.575 0.775 8.585 0.945 ;
        RECT 8.585 0.775 8.595 0.955 ;
        RECT 8.595 0.775 8.601 0.965 ;
        RECT 7.025 2.475 7.195 3.060 ;
        RECT 7.025 2.475 7.985 2.645 ;
        RECT 7.815 2.475 7.985 3.130 ;
        RECT 8.600 1.900 8.770 3.130 ;
        RECT 9.430 2.600 9.600 3.130 ;
        RECT 7.815 2.960 9.600 3.130 ;
        RECT 9.430 2.600 10.510 2.770 ;
        RECT 10.340 2.600 10.510 3.175 ;
        RECT 10.995 0.985 11.165 2.070 ;
        RECT 8.600 1.900 11.165 2.070 ;
        RECT 10.995 0.985 11.400 1.285 ;
        RECT 10.340 3.005 11.400 3.175 ;
        RECT 8.950 2.250 9.250 2.760 ;
        RECT 8.950 0.590 9.565 0.760 ;
        RECT 9.395 0.590 9.565 1.015 ;
        RECT 10.580 0.615 10.750 1.015 ;
        RECT 9.395 0.845 10.750 1.015 ;
        RECT 10.730 2.250 11.030 2.825 ;
        RECT 11.345 1.475 11.515 2.420 ;
        RECT 8.950 2.250 11.515 2.420 ;
        RECT 10.580 0.615 11.770 0.785 ;
        RECT 11.600 0.615 11.770 1.645 ;
        RECT 11.345 1.475 12.540 1.645 ;
        RECT 12.340 1.475 12.540 1.830 ;
        RECT 12.340 1.660 13.560 1.830 ;
        RECT 11.740 1.830 12.040 2.220 ;
        RECT 12.225 1.125 12.960 1.295 ;
        RECT 12.790 1.125 12.960 1.480 ;
        RECT 12.790 1.310 13.955 1.480 ;
        RECT 13.785 1.310 13.955 2.220 ;
        RECT 11.740 2.050 13.955 2.220 ;
  END 
END FFSDHQHD3XHT

MACRO FFSDHQHD2XHT
  CLASS  CORE ;
  FOREIGN FFSDHQHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.940 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.080 0.595 13.250 3.075 ;
        RECT 13.080 0.595 13.315 2.015 ;
        RECT 13.080 1.360 13.430 2.015 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 1.240 1.165 1.775 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.545 0.380 2.020 ;
        RECT 0.370 2.580 0.585 2.840 ;
        RECT 0.285 2.670 0.585 2.840 ;
        RECT 0.370 2.580 1.375 2.750 ;
        RECT 0.285 2.670 1.375 2.750 ;
        RECT 1.205 2.580 1.375 3.190 ;
        RECT 1.205 3.020 2.310 3.190 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.905 ;
        RECT 2.545 -0.300 2.845 0.595 ;
        RECT 3.535 -0.300 3.835 0.595 ;
        RECT 4.535 -0.300 4.835 0.595 ;
        RECT 7.435 -0.300 7.735 0.595 ;
        RECT 9.745 -0.300 10.045 0.665 ;
        RECT 11.865 -0.300 12.035 0.850 ;
        RECT 12.560 -0.300 12.730 0.780 ;
        RECT 13.600 -0.300 13.770 1.120 ;
        RECT 0.000 -0.300 13.940 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 4.535 1.605 5.100 2.020 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.610 2.505 2.020 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 3.060 0.955 3.990 ;
        RECT 2.555 2.830 2.730 3.990 ;
        RECT 3.575 2.770 3.875 3.990 ;
        RECT 4.445 2.770 4.745 3.990 ;
        RECT 7.450 2.870 7.750 3.990 ;
        RECT 9.740 2.880 10.040 3.990 ;
        RECT 11.695 2.590 11.865 3.990 ;
        RECT 12.560 2.910 12.730 3.990 ;
        RECT 13.600 2.230 13.770 3.990 ;
        RECT 0.000 3.390 13.940 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.085 0.730 1.255 ;
        RECT 0.560 1.085 0.730 2.400 ;
        RECT 0.105 2.230 0.730 2.400 ;
        RECT 1.355 1.460 1.525 2.125 ;
        RECT 0.560 1.955 1.525 2.125 ;
        RECT 1.355 1.460 1.965 1.760 ;
        RECT 3.400 1.605 3.570 1.905 ;
        RECT 3.400 1.605 4.295 1.790 ;
        RECT 3.995 1.125 4.295 2.215 ;
        RECT 5.085 1.125 5.755 1.295 ;
        RECT 5.585 1.125 5.755 2.215 ;
        RECT 5.320 2.045 5.755 2.215 ;
        RECT 1.575 2.330 1.875 2.840 ;
        RECT 1.575 0.825 2.460 1.005 ;
        RECT 1.575 2.330 2.685 2.500 ;
        RECT 2.630 0.775 6.115 0.945 ;
        RECT 5.945 0.775 6.115 2.320 ;
        RECT 2.685 1.285 2.695 2.499 ;
        RECT 2.695 1.295 2.705 2.499 ;
        RECT 2.705 1.305 2.715 2.499 ;
        RECT 2.715 1.315 2.725 2.499 ;
        RECT 2.725 1.325 2.735 2.499 ;
        RECT 2.735 1.335 2.745 2.499 ;
        RECT 2.745 1.345 2.755 2.499 ;
        RECT 2.755 1.355 2.765 2.499 ;
        RECT 2.765 1.365 2.775 2.499 ;
        RECT 2.775 1.375 2.785 2.499 ;
        RECT 2.785 1.385 2.795 2.499 ;
        RECT 2.795 1.395 2.805 2.499 ;
        RECT 2.805 1.405 2.815 2.499 ;
        RECT 2.815 1.415 2.825 2.499 ;
        RECT 2.825 1.425 2.835 2.499 ;
        RECT 2.835 1.435 2.845 2.499 ;
        RECT 2.845 1.445 2.855 2.499 ;
        RECT 2.630 1.230 2.640 1.464 ;
        RECT 2.640 1.240 2.650 1.474 ;
        RECT 2.650 1.250 2.660 1.484 ;
        RECT 2.660 1.260 2.670 1.494 ;
        RECT 2.670 1.270 2.680 1.504 ;
        RECT 2.680 1.275 2.686 1.515 ;
        RECT 2.460 0.775 2.470 1.295 ;
        RECT 2.470 0.775 2.480 1.305 ;
        RECT 2.480 0.775 2.490 1.315 ;
        RECT 2.490 0.775 2.500 1.325 ;
        RECT 2.500 0.775 2.510 1.335 ;
        RECT 2.510 0.775 2.520 1.345 ;
        RECT 2.520 0.775 2.530 1.355 ;
        RECT 2.530 0.775 2.540 1.365 ;
        RECT 2.540 0.775 2.550 1.375 ;
        RECT 2.550 0.775 2.560 1.385 ;
        RECT 2.560 0.775 2.570 1.395 ;
        RECT 2.570 0.775 2.580 1.405 ;
        RECT 2.580 0.775 2.590 1.415 ;
        RECT 2.590 0.775 2.600 1.425 ;
        RECT 2.600 0.775 2.610 1.435 ;
        RECT 2.610 0.775 2.620 1.445 ;
        RECT 2.620 0.775 2.630 1.455 ;
        RECT 6.645 1.060 6.815 2.340 ;
        RECT 7.730 1.520 7.900 2.210 ;
        RECT 6.645 2.040 7.900 2.210 ;
        RECT 7.730 1.520 8.005 1.820 ;
        RECT 7.355 1.170 7.525 1.820 ;
        RECT 8.025 1.125 8.355 1.340 ;
        RECT 7.355 1.170 8.355 1.340 ;
        RECT 8.090 2.040 8.260 2.340 ;
        RECT 8.185 1.125 8.355 2.210 ;
        RECT 8.090 2.040 8.355 2.210 ;
        RECT 8.185 1.570 10.175 1.740 ;
        RECT 3.050 1.125 3.220 2.735 ;
        RECT 3.050 2.095 3.250 2.735 ;
        RECT 3.015 1.125 3.315 1.295 ;
        RECT 3.050 2.400 5.375 2.590 ;
        RECT 5.205 2.400 5.375 2.900 ;
        RECT 6.295 0.550 6.465 2.900 ;
        RECT 5.205 2.730 6.465 2.900 ;
        RECT 6.295 0.550 7.155 0.730 ;
        RECT 6.985 0.550 7.155 0.945 ;
        RECT 6.985 0.775 8.435 0.945 ;
        RECT 8.715 0.970 9.110 1.140 ;
        RECT 8.940 0.970 9.110 1.365 ;
        RECT 8.940 1.195 10.720 1.365 ;
        RECT 10.550 1.195 10.720 1.675 ;
        RECT 8.630 0.895 8.640 1.139 ;
        RECT 8.640 0.905 8.650 1.139 ;
        RECT 8.650 0.915 8.660 1.139 ;
        RECT 8.660 0.925 8.670 1.139 ;
        RECT 8.670 0.935 8.680 1.139 ;
        RECT 8.680 0.945 8.690 1.139 ;
        RECT 8.690 0.955 8.700 1.139 ;
        RECT 8.700 0.965 8.710 1.139 ;
        RECT 8.710 0.970 8.716 1.140 ;
        RECT 8.520 0.785 8.530 1.029 ;
        RECT 8.530 0.795 8.540 1.039 ;
        RECT 8.540 0.805 8.550 1.049 ;
        RECT 8.550 0.815 8.560 1.059 ;
        RECT 8.560 0.825 8.570 1.069 ;
        RECT 8.570 0.835 8.580 1.079 ;
        RECT 8.580 0.845 8.590 1.089 ;
        RECT 8.590 0.855 8.600 1.099 ;
        RECT 8.600 0.865 8.610 1.109 ;
        RECT 8.610 0.875 8.620 1.119 ;
        RECT 8.620 0.885 8.630 1.129 ;
        RECT 8.435 0.775 8.445 0.945 ;
        RECT 8.445 0.775 8.455 0.955 ;
        RECT 8.455 0.775 8.465 0.965 ;
        RECT 8.465 0.775 8.475 0.975 ;
        RECT 8.475 0.775 8.485 0.985 ;
        RECT 8.485 0.775 8.495 0.995 ;
        RECT 8.495 0.775 8.505 1.005 ;
        RECT 8.505 0.775 8.515 1.015 ;
        RECT 8.515 0.775 8.521 1.025 ;
        RECT 6.760 2.520 7.060 2.835 ;
        RECT 8.540 1.990 8.710 2.690 ;
        RECT 6.760 2.520 8.710 2.690 ;
        RECT 10.925 0.985 11.095 2.160 ;
        RECT 8.540 1.990 11.095 2.160 ;
        RECT 10.925 0.985 11.275 1.285 ;
        RECT 8.890 2.475 9.060 3.115 ;
        RECT 8.795 0.590 9.560 0.760 ;
        RECT 9.390 0.590 9.560 1.015 ;
        RECT 10.550 0.615 10.720 1.015 ;
        RECT 9.390 0.845 10.720 1.015 ;
        RECT 10.700 2.475 10.870 3.115 ;
        RECT 11.275 1.550 11.445 2.645 ;
        RECT 8.890 2.475 11.445 2.645 ;
        RECT 10.550 0.615 11.645 0.785 ;
        RECT 11.475 0.615 11.645 1.720 ;
        RECT 11.275 1.550 12.485 1.720 ;
        RECT 11.660 1.925 11.830 2.225 ;
        RECT 12.020 1.125 12.860 1.295 ;
        RECT 12.670 1.125 12.860 2.225 ;
        RECT 11.660 2.055 12.860 2.225 ;
  END 
END FFSDHQHD2XHT

MACRO FFSDHDMXHT
  CLASS  CORE ;
  FOREIGN FFSDHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.070 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.730 1.060 10.970 1.360 ;
        RECT 10.760 1.060 10.970 2.280 ;
        RECT 10.730 1.980 10.970 2.280 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.625 1.125 10.150 1.295 ;
        RECT 9.940 1.125 10.150 2.215 ;
        RECT 9.625 2.045 10.150 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.415 -0.300 2.715 0.595 ;
        RECT 3.325 -0.300 3.625 0.595 ;
        RECT 5.815 -0.300 6.115 0.595 ;
        RECT 6.755 -0.300 7.055 0.595 ;
        RECT 8.655 -0.300 8.955 0.560 ;
        RECT 10.145 -0.300 10.445 0.595 ;
        RECT 0.000 -0.300 11.070 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.740 1.525 3.230 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.585 2.740 3.225 3.990 ;
        RECT 5.995 3.160 6.975 3.990 ;
        RECT 8.600 2.745 8.770 3.990 ;
        RECT 10.145 2.925 10.445 3.990 ;
        RECT 0.000 3.390 11.070 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.555 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.070 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.990 0.775 2.160 1.035 ;
        RECT 1.530 0.865 2.160 1.035 ;
        RECT 1.990 0.775 4.510 0.945 ;
        RECT 4.275 0.480 4.510 0.945 ;
        RECT 4.350 1.890 4.540 1.960 ;
        RECT 4.360 1.890 4.540 1.970 ;
        RECT 4.340 0.480 4.510 1.950 ;
        RECT 4.340 1.870 4.520 1.950 ;
        RECT 4.340 1.880 4.530 1.950 ;
        RECT 4.370 1.890 4.540 2.280 ;
        RECT 5.050 1.230 5.240 1.294 ;
        RECT 5.060 1.230 5.240 1.304 ;
        RECT 5.040 0.900 5.210 1.284 ;
        RECT 5.040 1.210 5.220 1.284 ;
        RECT 5.040 1.220 5.230 1.284 ;
        RECT 5.070 1.230 5.240 2.280 ;
        RECT 6.185 1.675 6.495 1.865 ;
        RECT 5.070 1.695 6.495 1.865 ;
        RECT 5.685 1.325 5.985 1.515 ;
        RECT 6.430 0.900 6.600 1.495 ;
        RECT 5.685 1.325 7.165 1.495 ;
        RECT 6.995 1.325 7.165 2.215 ;
        RECT 6.365 2.045 7.165 2.215 ;
        RECT 2.805 1.125 3.585 1.295 ;
        RECT 2.785 2.190 3.585 2.360 ;
        RECT 3.415 1.125 3.585 2.980 ;
        RECT 3.415 1.525 3.795 1.825 ;
        RECT 3.415 2.810 7.635 2.980 ;
        RECT 3.845 1.125 4.145 1.295 ;
        RECT 3.975 1.125 4.145 2.630 ;
        RECT 3.830 2.125 4.145 2.630 ;
        RECT 4.690 0.535 4.860 1.765 ;
        RECT 4.700 1.705 4.890 1.775 ;
        RECT 4.710 1.705 4.890 1.785 ;
        RECT 3.830 2.460 4.860 2.630 ;
        RECT 4.690 1.685 4.870 1.765 ;
        RECT 4.690 1.695 4.880 1.765 ;
        RECT 4.720 1.705 4.890 2.629 ;
        RECT 4.690 0.535 5.485 0.705 ;
        RECT 7.345 0.500 7.515 2.630 ;
        RECT 7.345 0.500 7.745 0.670 ;
        RECT 7.345 2.440 8.150 2.630 ;
        RECT 4.890 2.460 8.150 2.630 ;
        RECT 7.980 2.440 8.150 2.770 ;
        RECT 8.405 1.310 9.385 1.480 ;
        RECT 9.180 0.875 9.350 1.480 ;
        RECT 9.215 1.310 9.385 2.215 ;
        RECT 9.085 2.045 9.385 2.215 ;
        RECT 9.215 1.595 9.735 1.765 ;
        RECT 7.770 0.875 7.940 2.215 ;
        RECT 7.695 2.045 8.905 2.215 ;
        RECT 8.735 2.045 8.905 2.565 ;
        RECT 8.970 2.395 9.140 2.780 ;
        RECT 10.380 1.520 10.550 2.565 ;
        RECT 8.735 2.395 10.550 2.565 ;
        RECT 10.380 1.520 10.570 1.820 ;
  END 
END FFSDHDMXHT

MACRO FFSDHDLXHT
  CLASS  CORE ;
  FOREIGN FFSDHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.070 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.730 1.060 10.970 1.360 ;
        RECT 10.800 1.060 10.970 2.460 ;
        RECT 10.730 1.980 10.970 2.460 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.685 1.125 10.150 1.295 ;
        RECT 9.940 1.125 10.150 2.215 ;
        RECT 9.685 2.045 10.150 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.925 1.415 2.980 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.935 2.810 1.115 3.095 ;
        RECT 0.100 2.810 1.115 2.980 ;
        RECT 0.935 2.925 1.415 3.095 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.435 -0.300 2.735 0.595 ;
        RECT 3.405 -0.300 3.705 0.595 ;
        RECT 5.845 -0.300 6.145 0.635 ;
        RECT 6.815 -0.300 7.115 0.565 ;
        RECT 8.715 -0.300 9.015 0.560 ;
        RECT 10.115 -0.300 10.415 0.745 ;
        RECT 0.000 -0.300 11.070 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.790 1.525 3.280 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.455 3.160 0.755 3.990 ;
        RECT 2.645 2.710 3.285 3.990 ;
        RECT 6.050 3.160 7.030 3.990 ;
        RECT 8.660 2.745 8.830 3.990 ;
        RECT 10.115 2.745 10.415 3.990 ;
        RECT 0.000 3.390 11.070 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.045 0.975 2.215 ;
        RECT 0.105 0.975 1.180 1.145 ;
        RECT 1.350 0.480 1.575 0.650 ;
        RECT 1.370 2.555 1.870 2.725 ;
        RECT 1.700 2.555 1.870 2.855 ;
        RECT 1.285 2.480 1.295 2.724 ;
        RECT 1.295 2.490 1.305 2.724 ;
        RECT 1.305 2.500 1.315 2.724 ;
        RECT 1.315 2.510 1.325 2.724 ;
        RECT 1.325 2.520 1.335 2.724 ;
        RECT 1.335 2.530 1.345 2.724 ;
        RECT 1.345 2.540 1.355 2.724 ;
        RECT 1.355 2.550 1.365 2.724 ;
        RECT 1.365 2.555 1.371 2.725 ;
        RECT 1.275 0.480 1.285 2.020 ;
        RECT 1.285 0.480 1.295 2.010 ;
        RECT 1.295 0.480 1.305 2.000 ;
        RECT 1.305 0.480 1.315 1.990 ;
        RECT 1.315 0.480 1.325 1.980 ;
        RECT 1.325 0.480 1.335 1.970 ;
        RECT 1.335 0.480 1.345 1.960 ;
        RECT 1.345 0.480 1.351 1.954 ;
        RECT 1.275 2.470 1.285 2.714 ;
        RECT 1.180 0.480 1.190 2.620 ;
        RECT 1.190 0.480 1.200 2.630 ;
        RECT 1.200 0.480 1.210 2.640 ;
        RECT 1.210 0.480 1.220 2.650 ;
        RECT 1.220 0.480 1.230 2.660 ;
        RECT 1.230 0.480 1.240 2.670 ;
        RECT 1.240 0.480 1.250 2.680 ;
        RECT 1.250 0.480 1.260 2.690 ;
        RECT 1.260 0.480 1.270 2.700 ;
        RECT 1.270 0.480 1.276 2.710 ;
        RECT 1.105 1.915 1.115 2.545 ;
        RECT 1.115 1.905 1.125 2.555 ;
        RECT 1.125 1.895 1.135 2.565 ;
        RECT 1.135 1.885 1.145 2.575 ;
        RECT 1.145 1.875 1.155 2.585 ;
        RECT 1.155 1.865 1.165 2.595 ;
        RECT 1.165 1.855 1.175 2.605 ;
        RECT 1.175 1.845 1.181 2.615 ;
        RECT 0.975 2.045 0.985 2.215 ;
        RECT 0.985 2.035 0.995 2.215 ;
        RECT 0.995 2.025 1.005 2.215 ;
        RECT 1.005 2.015 1.015 2.215 ;
        RECT 1.015 2.005 1.025 2.215 ;
        RECT 1.025 1.995 1.035 2.215 ;
        RECT 1.035 1.985 1.045 2.215 ;
        RECT 1.045 1.975 1.055 2.215 ;
        RECT 1.055 1.965 1.065 2.215 ;
        RECT 1.065 1.955 1.075 2.215 ;
        RECT 1.075 1.945 1.085 2.215 ;
        RECT 1.085 1.935 1.095 2.215 ;
        RECT 1.095 1.925 1.105 2.215 ;
        RECT 1.550 0.865 1.720 2.340 ;
        RECT 1.520 2.040 1.720 2.340 ;
        RECT 2.000 0.775 2.170 1.035 ;
        RECT 1.550 0.865 2.170 1.035 ;
        RECT 2.000 0.775 4.550 0.945 ;
        RECT 4.375 0.500 4.550 0.945 ;
        RECT 4.380 0.500 4.550 2.280 ;
        RECT 5.080 0.900 5.250 2.280 ;
        RECT 6.215 1.675 6.515 1.865 ;
        RECT 5.080 1.695 6.515 1.865 ;
        RECT 5.735 1.325 6.035 1.515 ;
        RECT 6.490 0.900 6.660 1.495 ;
        RECT 5.735 1.325 6.905 1.495 ;
        RECT 6.735 1.325 6.905 2.215 ;
        RECT 6.415 2.045 6.905 2.215 ;
        RECT 6.735 1.410 7.225 1.580 ;
        RECT 2.825 1.125 3.635 1.295 ;
        RECT 2.765 2.190 3.635 2.360 ;
        RECT 3.465 1.125 3.635 2.980 ;
        RECT 3.465 1.525 3.760 1.825 ;
        RECT 3.465 2.810 7.685 2.980 ;
        RECT 3.940 1.125 4.135 2.630 ;
        RECT 3.835 2.125 4.135 2.630 ;
        RECT 3.865 1.125 4.165 1.295 ;
        RECT 4.730 0.535 4.900 2.630 ;
        RECT 4.730 0.535 5.525 0.705 ;
        RECT 7.405 1.425 7.575 2.630 ;
        RECT 7.470 0.500 7.640 1.595 ;
        RECT 7.405 1.425 7.640 1.595 ;
        RECT 7.470 0.500 7.805 0.670 ;
        RECT 7.405 2.440 8.210 2.630 ;
        RECT 3.835 2.460 8.210 2.630 ;
        RECT 8.040 2.440 8.210 2.770 ;
        RECT 8.465 1.415 9.445 1.585 ;
        RECT 9.240 0.875 9.410 1.585 ;
        RECT 9.275 1.415 9.445 2.215 ;
        RECT 9.145 2.045 9.445 2.215 ;
        RECT 9.275 1.650 9.760 1.820 ;
        RECT 7.830 0.875 8.000 2.215 ;
        RECT 7.755 2.045 8.965 2.215 ;
        RECT 8.795 2.045 8.965 2.565 ;
        RECT 9.030 2.395 9.200 2.695 ;
        RECT 10.380 1.520 10.550 2.565 ;
        RECT 8.795 2.395 10.550 2.565 ;
        RECT 10.380 1.520 10.580 1.820 ;
  END 
END FFSDHDLXHT

MACRO FFSDHD1XHT
  CLASS  CORE ;
  FOREIGN FFSDHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.070 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.730 0.720 10.970 1.360 ;
        RECT 10.760 0.720 10.970 2.960 ;
        RECT 10.730 1.980 10.970 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.690 0.720 9.860 1.405 ;
        RECT 9.690 1.235 10.150 1.405 ;
        RECT 9.940 1.235 10.150 2.235 ;
        RECT 9.625 2.065 10.150 2.235 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.500 0.595 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.385 -0.300 2.685 0.595 ;
        RECT 3.335 -0.300 3.635 0.595 ;
        RECT 5.815 -0.300 6.115 0.595 ;
        RECT 6.755 -0.300 7.055 0.595 ;
        RECT 8.710 -0.300 8.880 0.535 ;
        RECT 10.145 -0.300 10.445 1.055 ;
        RECT 0.000 -0.300 11.070 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.740 1.525 3.230 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.385 2.700 2.685 3.990 ;
        RECT 3.125 2.675 3.295 3.990 ;
        RECT 6.010 3.160 6.990 3.990 ;
        RECT 8.600 2.765 8.770 3.990 ;
        RECT 10.145 2.975 10.445 3.990 ;
        RECT 0.000 3.390 11.070 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.555 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.150 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.985 0.775 2.155 1.035 ;
        RECT 1.530 0.865 2.155 1.035 ;
        RECT 1.985 0.775 4.510 0.945 ;
        RECT 4.340 0.775 4.510 2.280 ;
        RECT 5.040 0.900 5.210 2.280 ;
        RECT 6.185 1.675 6.495 1.865 ;
        RECT 5.040 1.695 6.495 1.865 ;
        RECT 5.685 1.325 5.985 1.515 ;
        RECT 6.430 0.910 6.600 1.495 ;
        RECT 5.685 1.325 7.165 1.495 ;
        RECT 6.995 1.325 7.165 2.215 ;
        RECT 6.365 2.045 7.165 2.215 ;
        RECT 2.785 1.125 3.585 1.295 ;
        RECT 2.785 2.190 3.645 2.360 ;
        RECT 3.415 1.125 3.585 2.360 ;
        RECT 3.475 1.525 3.645 2.980 ;
        RECT 3.415 1.525 3.710 1.825 ;
        RECT 3.475 2.810 7.745 2.980 ;
        RECT 3.765 1.125 4.085 1.295 ;
        RECT 3.830 1.980 4.085 2.280 ;
        RECT 3.915 1.125 4.085 2.630 ;
        RECT 4.690 0.535 4.860 2.630 ;
        RECT 4.690 0.535 5.485 0.705 ;
        RECT 7.345 0.500 7.515 2.630 ;
        RECT 7.345 0.500 7.745 0.670 ;
        RECT 7.345 2.440 8.125 2.630 ;
        RECT 7.955 2.440 8.125 2.705 ;
        RECT 3.915 2.460 8.125 2.630 ;
        RECT 7.955 2.535 8.255 2.705 ;
        RECT 8.405 1.220 9.385 1.390 ;
        RECT 9.180 0.785 9.350 1.390 ;
        RECT 9.215 1.220 9.385 2.215 ;
        RECT 9.085 2.045 9.385 2.215 ;
        RECT 9.215 1.585 9.760 1.885 ;
        RECT 7.760 0.875 7.930 2.215 ;
        RECT 7.695 2.045 8.905 2.215 ;
        RECT 8.735 2.045 8.905 2.585 ;
        RECT 8.970 2.415 9.140 2.780 ;
        RECT 10.380 1.520 10.550 2.585 ;
        RECT 8.735 2.415 10.550 2.585 ;
        RECT 10.380 1.520 10.570 1.820 ;
  END 
END FFSDHD1XHT

MACRO FFSDHD2XHT
  CLASS  CORE ;
  FOREIGN FFSDHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.300 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.440 0.720 11.610 2.960 ;
        RECT 11.440 1.645 11.790 2.015 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.350 0.720 10.570 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.265 -0.300 2.565 0.595 ;
        RECT 3.325 -0.300 3.625 0.595 ;
        RECT 5.765 -0.300 6.065 0.595 ;
        RECT 6.780 -0.300 7.080 0.715 ;
        RECT 8.525 -0.300 8.695 0.780 ;
        RECT 9.880 -0.300 10.050 1.120 ;
        RECT 10.920 -0.300 11.090 1.120 ;
        RECT 11.960 -0.300 12.130 1.120 ;
        RECT 0.000 -0.300 12.300 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.730 1.525 3.220 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.520 2.360 2.435 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.555 2.700 3.195 3.990 ;
        RECT 5.910 3.160 6.210 3.990 ;
        RECT 6.750 3.095 7.050 3.990 ;
        RECT 8.645 2.805 8.815 3.990 ;
        RECT 9.815 2.975 10.115 3.990 ;
        RECT 10.855 2.975 11.155 3.990 ;
        RECT 11.895 2.295 12.195 3.990 ;
        RECT 0.000 3.390 12.300 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.555 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.150 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.970 0.775 2.140 1.035 ;
        RECT 1.530 0.865 2.140 1.035 ;
        RECT 1.970 0.775 4.500 0.945 ;
        RECT 4.330 0.775 4.500 2.280 ;
        RECT 5.030 0.910 5.200 2.280 ;
        RECT 6.135 1.675 6.435 1.865 ;
        RECT 5.030 1.695 6.435 1.865 ;
        RECT 5.625 1.325 5.925 1.515 ;
        RECT 6.380 0.910 6.550 1.495 ;
        RECT 5.625 1.325 7.170 1.495 ;
        RECT 7.000 1.325 7.170 2.215 ;
        RECT 6.350 2.045 7.170 2.215 ;
        RECT 2.775 1.125 3.575 1.295 ;
        RECT 2.775 2.190 3.575 2.360 ;
        RECT 3.405 1.125 3.575 3.035 ;
        RECT 3.405 1.525 3.700 1.825 ;
        RECT 3.405 2.865 5.525 3.035 ;
        RECT 5.765 2.745 7.265 2.915 ;
        RECT 7.650 3.040 8.250 3.210 ;
        RECT 7.560 2.960 7.570 3.210 ;
        RECT 7.570 2.970 7.580 3.210 ;
        RECT 7.580 2.980 7.590 3.210 ;
        RECT 7.590 2.990 7.600 3.210 ;
        RECT 7.600 3.000 7.610 3.210 ;
        RECT 7.610 3.010 7.620 3.210 ;
        RECT 7.620 3.020 7.630 3.210 ;
        RECT 7.630 3.030 7.640 3.210 ;
        RECT 7.640 3.040 7.650 3.210 ;
        RECT 7.355 2.755 7.365 3.005 ;
        RECT 7.365 2.765 7.375 3.015 ;
        RECT 7.375 2.775 7.385 3.025 ;
        RECT 7.385 2.785 7.395 3.035 ;
        RECT 7.395 2.795 7.405 3.045 ;
        RECT 7.405 2.805 7.415 3.055 ;
        RECT 7.415 2.815 7.425 3.065 ;
        RECT 7.425 2.825 7.435 3.075 ;
        RECT 7.435 2.835 7.445 3.085 ;
        RECT 7.445 2.845 7.455 3.095 ;
        RECT 7.455 2.855 7.465 3.105 ;
        RECT 7.465 2.865 7.475 3.115 ;
        RECT 7.475 2.875 7.485 3.125 ;
        RECT 7.485 2.885 7.495 3.135 ;
        RECT 7.495 2.895 7.505 3.145 ;
        RECT 7.505 2.905 7.515 3.155 ;
        RECT 7.515 2.915 7.525 3.165 ;
        RECT 7.525 2.925 7.535 3.175 ;
        RECT 7.535 2.935 7.545 3.185 ;
        RECT 7.545 2.945 7.555 3.195 ;
        RECT 7.555 2.950 7.561 3.204 ;
        RECT 7.265 2.745 7.275 2.915 ;
        RECT 7.275 2.745 7.285 2.925 ;
        RECT 7.285 2.745 7.295 2.935 ;
        RECT 7.295 2.745 7.305 2.945 ;
        RECT 7.305 2.745 7.315 2.955 ;
        RECT 7.315 2.745 7.325 2.965 ;
        RECT 7.325 2.745 7.335 2.975 ;
        RECT 7.335 2.745 7.345 2.985 ;
        RECT 7.345 2.745 7.355 2.995 ;
        RECT 5.645 2.745 5.655 3.025 ;
        RECT 5.655 2.745 5.665 3.015 ;
        RECT 5.665 2.745 5.675 3.005 ;
        RECT 5.675 2.745 5.685 2.995 ;
        RECT 5.685 2.745 5.695 2.985 ;
        RECT 5.695 2.745 5.705 2.975 ;
        RECT 5.705 2.745 5.715 2.965 ;
        RECT 5.715 2.745 5.725 2.955 ;
        RECT 5.725 2.745 5.735 2.945 ;
        RECT 5.735 2.745 5.745 2.935 ;
        RECT 5.745 2.745 5.755 2.925 ;
        RECT 5.755 2.745 5.765 2.915 ;
        RECT 5.525 2.865 5.535 3.035 ;
        RECT 5.535 2.855 5.545 3.035 ;
        RECT 5.545 2.845 5.555 3.035 ;
        RECT 5.555 2.835 5.565 3.035 ;
        RECT 5.565 2.825 5.575 3.035 ;
        RECT 5.575 2.815 5.585 3.035 ;
        RECT 5.585 2.805 5.595 3.035 ;
        RECT 5.595 2.795 5.605 3.035 ;
        RECT 5.605 2.785 5.615 3.035 ;
        RECT 5.615 2.775 5.625 3.035 ;
        RECT 5.625 2.765 5.635 3.035 ;
        RECT 5.635 2.755 5.645 3.035 ;
        RECT 3.755 1.125 4.075 1.295 ;
        RECT 3.905 1.125 4.075 2.685 ;
        RECT 3.820 1.980 4.075 2.685 ;
        RECT 4.680 0.535 4.850 2.685 ;
        RECT 3.820 2.515 5.225 2.685 ;
        RECT 5.345 2.395 5.385 2.685 ;
        RECT 4.680 0.535 5.445 0.705 ;
        RECT 7.350 0.710 7.435 2.565 ;
        RECT 5.505 2.395 7.435 2.565 ;
        RECT 7.520 0.710 8.290 0.880 ;
        RECT 7.685 2.560 8.250 2.730 ;
        RECT 8.120 0.710 8.290 1.140 ;
        RECT 8.875 0.480 9.045 1.140 ;
        RECT 8.120 0.970 9.045 1.140 ;
        RECT 8.875 0.480 9.700 0.650 ;
        RECT 7.600 2.485 7.610 2.729 ;
        RECT 7.610 2.495 7.620 2.729 ;
        RECT 7.620 2.505 7.630 2.729 ;
        RECT 7.630 2.515 7.640 2.729 ;
        RECT 7.640 2.525 7.650 2.729 ;
        RECT 7.650 2.535 7.660 2.729 ;
        RECT 7.660 2.545 7.670 2.729 ;
        RECT 7.670 2.555 7.680 2.729 ;
        RECT 7.680 2.560 7.686 2.730 ;
        RECT 7.520 2.405 7.530 2.649 ;
        RECT 7.530 2.415 7.540 2.659 ;
        RECT 7.540 2.425 7.550 2.669 ;
        RECT 7.550 2.435 7.560 2.679 ;
        RECT 7.560 2.445 7.570 2.689 ;
        RECT 7.570 2.455 7.580 2.699 ;
        RECT 7.580 2.465 7.590 2.709 ;
        RECT 7.590 2.475 7.600 2.719 ;
        RECT 7.435 0.710 7.445 2.564 ;
        RECT 7.445 0.710 7.455 2.574 ;
        RECT 7.455 0.710 7.465 2.584 ;
        RECT 7.465 0.710 7.475 2.594 ;
        RECT 7.475 0.710 7.485 2.604 ;
        RECT 7.485 0.710 7.495 2.614 ;
        RECT 7.495 0.710 7.505 2.624 ;
        RECT 7.505 0.710 7.515 2.634 ;
        RECT 7.515 0.710 7.521 2.644 ;
        RECT 5.385 2.395 5.395 2.675 ;
        RECT 5.395 2.395 5.405 2.665 ;
        RECT 5.405 2.395 5.415 2.655 ;
        RECT 5.415 2.395 5.425 2.645 ;
        RECT 5.425 2.395 5.435 2.635 ;
        RECT 5.435 2.395 5.445 2.625 ;
        RECT 5.445 2.395 5.455 2.615 ;
        RECT 5.455 2.395 5.465 2.605 ;
        RECT 5.465 2.395 5.475 2.595 ;
        RECT 5.475 2.395 5.485 2.585 ;
        RECT 5.485 2.395 5.495 2.575 ;
        RECT 5.495 2.395 5.505 2.565 ;
        RECT 5.225 2.515 5.235 2.685 ;
        RECT 5.235 2.505 5.245 2.685 ;
        RECT 5.245 2.495 5.255 2.685 ;
        RECT 5.255 2.485 5.265 2.685 ;
        RECT 5.265 2.475 5.275 2.685 ;
        RECT 5.275 2.465 5.285 2.685 ;
        RECT 5.285 2.455 5.295 2.685 ;
        RECT 5.295 2.445 5.305 2.685 ;
        RECT 5.305 2.435 5.315 2.685 ;
        RECT 5.315 2.425 5.325 2.685 ;
        RECT 5.325 2.415 5.335 2.685 ;
        RECT 5.335 2.405 5.345 2.685 ;
        RECT 9.225 1.060 9.395 2.280 ;
        RECT 8.440 1.675 10.170 1.845 ;
        RECT 7.765 1.060 7.935 2.230 ;
        RECT 7.700 2.060 9.045 2.230 ;
        RECT 8.875 2.060 9.045 2.630 ;
        RECT 9.015 2.460 9.185 3.190 ;
        RECT 11.090 1.610 11.260 2.630 ;
        RECT 8.875 2.460 11.260 2.630 ;
  END 
END FFSDHD2XHT

MACRO FFSDHD1XSPGHT
  CLASS  CORE ;
  FOREIGN FFSDHD1XSPGHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.070 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 10.185 0.300 10.725 3.075 ;
      LAYER V7 ;
        RECT 10.275 2.075 10.635 2.435 ;
      LAYER M7 ;
        RECT 9.985 2.065 10.865 2.445 ;
      LAYER V6 ;
        RECT 10.360 2.160 10.550 2.350 ;
      LAYER M4 ;
        RECT 10.355 1.785 10.555 2.585 ;
      LAYER V3 ;
        RECT 10.360 2.160 10.550 2.350 ;
      LAYER M3 ;
        RECT 10.240 2.155 10.965 2.355 ;
        RECT 10.765 2.090 10.965 2.425 ;
      LAYER V2 ;
        RECT 10.770 2.160 10.960 2.350 ;
      LAYER M2 ;
        RECT 10.765 1.745 10.965 2.515 ;
      LAYER V1 ;
        RECT 10.770 2.160 10.960 2.350 ;
      LAYER M1 ;
        RECT 10.730 0.720 10.970 1.360 ;
        RECT 10.760 0.720 10.970 2.960 ;
        RECT 10.730 1.980 10.970 2.960 ;
      LAYER M6 ;
        RECT 10.355 1.030 10.555 3.075 ;
      LAYER V5 ;
        RECT 10.360 2.160 10.550 2.350 ;
      LAYER M5 ;
        RECT 9.985 2.155 10.865 2.355 ;
      LAYER V4 ;
        RECT 10.360 2.160 10.550 2.350 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 8.955 0.300 9.495 3.075 ;
      LAYER V7 ;
        RECT 9.045 1.255 9.405 1.615 ;
      LAYER M7 ;
        RECT 8.575 1.245 9.825 1.625 ;
      LAYER V6 ;
        RECT 9.130 1.340 9.320 1.530 ;
      LAYER M4 ;
        RECT 9.125 0.915 9.325 1.840 ;
      LAYER V3 ;
        RECT 9.130 1.340 9.320 1.530 ;
      LAYER M3 ;
        RECT 8.985 1.335 10.235 1.535 ;
      LAYER V2 ;
        RECT 9.950 1.340 10.140 1.530 ;
      LAYER M2 ;
        RECT 9.945 1.030 10.145 1.840 ;
      LAYER V1 ;
        RECT 9.950 1.340 10.140 1.530 ;
      LAYER M1 ;
        RECT 9.690 0.720 9.860 1.405 ;
        RECT 9.690 1.235 10.150 1.405 ;
        RECT 9.940 1.235 10.150 2.235 ;
        RECT 9.625 2.065 10.150 2.235 ;
      LAYER M6 ;
        RECT 9.125 1.030 9.325 3.075 ;
      LAYER V5 ;
        RECT 9.130 1.340 9.320 1.530 ;
      LAYER M5 ;
        RECT 8.575 1.335 9.825 1.535 ;
      LAYER V4 ;
        RECT 9.130 1.340 9.320 1.530 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 1.575 0.300 2.115 3.075 ;
      LAYER V7 ;
        RECT 1.665 1.255 2.025 1.615 ;
      LAYER M7 ;
        RECT 1.100 1.245 2.115 1.625 ;
      LAYER V6 ;
        RECT 1.750 1.340 1.940 1.530 ;
      LAYER M4 ;
        RECT 1.745 0.810 1.945 1.735 ;
      LAYER V3 ;
        RECT 1.750 1.340 1.940 1.530 ;
      LAYER M3 ;
        RECT 0.395 1.335 2.065 1.535 ;
      LAYER V2 ;
        RECT 0.520 1.340 0.710 1.530 ;
      LAYER M2 ;
        RECT 0.515 0.915 0.715 1.735 ;
      LAYER V1 ;
        RECT 0.520 1.340 0.710 1.530 ;
      LAYER M1 ;
        RECT 0.450 1.330 1.000 1.735 ;
      LAYER M6 ;
        RECT 1.745 1.030 1.945 3.075 ;
      LAYER V5 ;
        RECT 1.750 1.340 1.940 1.530 ;
      LAYER M5 ;
        RECT 1.100 1.335 2.115 1.535 ;
      LAYER V4 ;
        RECT 1.750 1.340 1.940 1.530 ;
    END
  END D
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 0.345 0.300 0.885 3.075 ;
      LAYER V7 ;
        RECT 0.435 2.485 0.795 2.845 ;
      LAYER M7 ;
        RECT 0.175 2.475 1.160 2.855 ;
      LAYER V6 ;
        RECT 0.520 2.570 0.710 2.760 ;
      LAYER M4 ;
        RECT 0.515 2.255 0.715 2.980 ;
      LAYER V3 ;
        RECT 0.520 2.570 0.710 2.760 ;
      LAYER M3 ;
        RECT 0.105 2.500 0.305 2.830 ;
        RECT 0.105 2.565 0.955 2.765 ;
      LAYER V2 ;
        RECT 0.110 2.570 0.300 2.760 ;
      LAYER M2 ;
        RECT 0.105 2.255 0.305 2.980 ;
      LAYER V1 ;
        RECT 0.110 2.570 0.300 2.760 ;
      LAYER M1 ;
        RECT 0.100 2.500 0.595 2.980 ;
        RECT 0.100 2.810 1.460 2.980 ;
        RECT 1.290 2.810 1.460 3.160 ;
      LAYER M6 ;
        RECT 0.515 1.030 0.715 3.075 ;
      LAYER V5 ;
        RECT 0.520 2.570 0.710 2.760 ;
      LAYER M5 ;
        RECT 0.175 2.565 1.160 2.765 ;
      LAYER V4 ;
        RECT 0.520 2.570 0.710 2.760 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.595 ;
        RECT 2.385 -0.300 2.685 0.595 ;
        RECT 3.335 -0.300 3.635 0.595 ;
        RECT 5.815 -0.300 6.115 0.595 ;
        RECT 6.755 -0.300 7.055 0.595 ;
        RECT 8.710 -0.300 8.880 0.535 ;
        RECT 10.145 -0.300 10.445 1.055 ;
        RECT 0.000 -0.300 11.070 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M8 ;
        RECT 4.035 0.300 4.575 3.070 ;
      LAYER V7 ;
        RECT 4.125 1.665 4.485 2.025 ;
      LAYER M7 ;
        RECT 3.800 1.655 4.795 2.035 ;
      LAYER V6 ;
        RECT 4.210 1.750 4.400 1.940 ;
      LAYER M4 ;
        RECT 4.205 1.530 4.405 2.290 ;
      LAYER V3 ;
        RECT 4.210 1.750 4.400 1.940 ;
      LAYER M3 ;
        RECT 2.890 1.745 4.575 1.945 ;
      LAYER V2 ;
        RECT 2.980 1.750 3.170 1.940 ;
      LAYER M2 ;
        RECT 2.975 1.455 3.175 2.210 ;
      LAYER V1 ;
        RECT 2.980 1.750 3.170 1.940 ;
      LAYER M1 ;
        RECT 2.740 1.525 3.230 2.010 ;
      LAYER M6 ;
        RECT 4.205 1.030 4.405 3.075 ;
      LAYER V5 ;
        RECT 4.210 1.750 4.400 1.940 ;
      LAYER M5 ;
        RECT 3.800 1.745 4.780 1.945 ;
      LAYER V4 ;
        RECT 4.210 1.750 4.400 1.940 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 2.805 0.300 3.345 3.070 ;
      LAYER V7 ;
        RECT 2.895 2.075 3.255 2.435 ;
      LAYER M7 ;
        RECT 2.425 2.065 3.345 2.445 ;
      LAYER V6 ;
        RECT 2.980 2.160 3.170 2.350 ;
      LAYER M4 ;
        RECT 2.975 1.970 3.175 2.820 ;
      LAYER V3 ;
        RECT 2.980 2.160 3.170 2.350 ;
      LAYER M3 ;
        RECT 2.040 2.155 3.290 2.355 ;
      LAYER V2 ;
        RECT 2.160 2.160 2.350 2.350 ;
      LAYER M2 ;
        RECT 2.155 1.430 2.355 2.485 ;
      LAYER V1 ;
        RECT 2.160 1.520 2.350 1.710 ;
      LAYER M1 ;
        RECT 2.030 1.290 2.440 1.800 ;
      LAYER M6 ;
        RECT 2.975 1.030 3.175 3.075 ;
      LAYER V5 ;
        RECT 2.980 2.160 3.170 2.350 ;
      LAYER M5 ;
        RECT 2.425 2.155 3.345 2.355 ;
      LAYER V4 ;
        RECT 2.980 2.160 3.170 2.350 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.160 0.835 3.990 ;
        RECT 2.385 2.700 2.685 3.990 ;
        RECT 3.125 2.675 3.295 3.990 ;
        RECT 6.010 3.160 6.990 3.990 ;
        RECT 8.600 2.765 8.770 3.990 ;
        RECT 10.145 2.975 10.445 3.990 ;
        RECT 0.000 3.390 11.070 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.975 1.350 1.145 ;
        RECT 0.105 2.045 1.350 2.215 ;
        RECT 1.180 0.480 1.350 2.630 ;
        RECT 1.180 0.480 1.555 0.650 ;
        RECT 1.180 2.460 1.940 2.630 ;
        RECT 1.770 2.460 1.940 3.150 ;
        RECT 1.530 0.865 1.700 2.280 ;
        RECT 1.985 0.775 2.155 1.035 ;
        RECT 1.530 0.865 2.155 1.035 ;
        RECT 1.985 0.775 4.510 0.945 ;
        RECT 4.340 0.775 4.510 2.280 ;
        RECT 5.040 0.900 5.210 2.280 ;
        RECT 6.185 1.675 6.495 1.865 ;
        RECT 5.040 1.695 6.495 1.865 ;
        RECT 5.685 1.325 5.985 1.515 ;
        RECT 6.430 0.910 6.600 1.495 ;
        RECT 5.685 1.325 7.165 1.495 ;
        RECT 6.995 1.325 7.165 2.215 ;
        RECT 6.365 2.045 7.165 2.215 ;
        RECT 2.785 1.125 3.585 1.295 ;
        RECT 2.785 2.190 3.645 2.360 ;
        RECT 3.415 1.125 3.585 2.360 ;
        RECT 3.475 1.525 3.645 2.980 ;
        RECT 3.415 1.525 3.710 1.825 ;
        RECT 3.475 2.810 7.745 2.980 ;
        RECT 3.765 1.125 4.085 1.295 ;
        RECT 3.830 1.980 4.085 2.280 ;
        RECT 3.915 1.125 4.085 2.630 ;
        RECT 4.690 0.535 4.860 2.630 ;
        RECT 4.690 0.535 5.485 0.705 ;
        RECT 7.345 0.500 7.515 2.630 ;
        RECT 7.345 0.500 7.745 0.670 ;
        RECT 7.345 2.440 8.125 2.630 ;
        RECT 7.955 2.440 8.125 2.705 ;
        RECT 3.915 2.460 8.125 2.630 ;
        RECT 7.955 2.535 8.255 2.705 ;
        RECT 8.405 1.220 9.385 1.390 ;
        RECT 9.180 0.785 9.350 1.390 ;
        RECT 9.215 1.220 9.385 2.215 ;
        RECT 9.085 2.045 9.385 2.215 ;
        RECT 9.215 1.585 9.760 1.885 ;
        RECT 7.760 0.875 7.930 2.215 ;
        RECT 7.695 2.045 8.905 2.215 ;
        RECT 8.735 2.045 8.905 2.585 ;
        RECT 8.970 2.415 9.140 2.780 ;
        RECT 10.380 1.520 10.550 2.585 ;
        RECT 8.735 2.415 10.550 2.585 ;
        RECT 10.380 1.520 10.570 1.820 ;
  END 
END FFSDHD1XSPGHT

MACRO FFSDCRHDMXHT
  CLASS  CORE ;
  FOREIGN FFSDCRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.890 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.550 1.060 11.790 1.360 ;
        RECT 11.580 1.060 11.790 2.435 ;
        RECT 11.550 1.980 11.790 2.435 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.510 1.060 10.680 1.470 ;
        RECT 10.510 2.000 10.680 2.300 ;
        RECT 10.510 1.290 10.970 1.470 ;
        RECT 10.760 1.290 10.970 2.235 ;
        RECT 10.510 2.000 10.970 2.235 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.935 2.485 2.390 2.950 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.455 1.625 3.075 1.950 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.960 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 -0.300 0.890 0.800 ;
        RECT 2.865 -0.300 3.165 0.595 ;
        RECT 4.020 -0.300 4.320 0.595 ;
        RECT 6.635 -0.300 6.935 0.595 ;
        RECT 7.575 -0.300 7.875 0.645 ;
        RECT 9.465 -0.300 9.765 0.560 ;
        RECT 10.965 -0.300 11.265 0.595 ;
        RECT 0.000 -0.300 11.890 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 3.560 1.525 4.050 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.780 1.330 1.190 1.820 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 2.650 0.890 3.990 ;
        RECT 2.590 2.845 2.760 3.990 ;
        RECT 3.945 2.675 4.115 3.990 ;
        RECT 6.825 3.160 7.805 3.990 ;
        RECT 9.420 2.830 9.590 3.990 ;
        RECT 10.965 2.925 11.265 3.990 ;
        RECT 0.000 3.390 11.890 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.980 0.340 2.280 ;
        RECT 0.170 2.110 1.275 2.280 ;
        RECT 1.105 0.555 1.275 1.150 ;
        RECT 0.170 0.980 1.275 1.150 ;
        RECT 1.105 2.110 1.275 2.885 ;
        RECT 1.105 2.715 1.575 2.885 ;
        RECT 1.105 0.555 2.055 0.725 ;
        RECT 1.975 2.130 3.255 2.300 ;
        RECT 1.520 1.060 1.690 2.280 ;
        RECT 2.455 0.775 2.625 1.230 ;
        RECT 1.520 1.060 2.625 1.230 ;
        RECT 2.455 0.775 5.330 0.945 ;
        RECT 5.160 0.775 5.330 2.280 ;
        RECT 5.860 0.900 6.030 2.280 ;
        RECT 7.005 1.675 7.315 1.865 ;
        RECT 5.860 1.695 7.315 1.865 ;
        RECT 6.505 1.325 6.805 1.515 ;
        RECT 7.250 0.900 7.420 1.495 ;
        RECT 6.505 1.325 7.985 1.495 ;
        RECT 7.815 1.325 7.985 2.215 ;
        RECT 7.185 2.045 7.985 2.215 ;
        RECT 3.455 1.125 4.405 1.295 ;
        RECT 3.485 2.190 4.465 2.360 ;
        RECT 4.235 1.125 4.405 2.360 ;
        RECT 4.295 1.525 4.465 2.980 ;
        RECT 4.235 1.525 4.530 1.825 ;
        RECT 4.295 2.810 8.465 2.980 ;
        RECT 4.585 1.125 4.905 1.295 ;
        RECT 4.650 1.980 4.905 2.280 ;
        RECT 4.735 1.125 4.905 2.630 ;
        RECT 5.510 0.535 5.680 2.630 ;
        RECT 5.510 0.535 6.305 0.705 ;
        RECT 8.165 1.425 8.335 2.630 ;
        RECT 8.230 0.500 8.400 1.595 ;
        RECT 8.165 1.425 8.400 1.595 ;
        RECT 8.230 0.500 8.565 0.670 ;
        RECT 8.165 2.440 8.970 2.630 ;
        RECT 4.735 2.460 8.970 2.630 ;
        RECT 8.800 2.440 8.970 2.770 ;
        RECT 9.225 1.430 10.330 1.600 ;
        RECT 10.000 0.875 10.170 1.600 ;
        RECT 10.160 1.430 10.330 2.215 ;
        RECT 9.905 2.045 10.330 2.215 ;
        RECT 10.160 1.650 10.555 1.820 ;
        RECT 8.590 0.875 8.760 2.215 ;
        RECT 8.515 2.045 9.595 2.215 ;
        RECT 9.425 2.045 9.595 2.650 ;
        RECT 9.790 2.480 9.960 2.780 ;
        RECT 11.200 1.520 11.370 2.650 ;
        RECT 9.425 2.480 11.370 2.650 ;
        RECT 11.200 1.520 11.390 1.820 ;
  END 
END FFSDCRHDMXHT

MACRO FFSDCRHDLXHT
  CLASS  CORE ;
  FOREIGN FFSDCRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.480 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.140 1.060 11.380 1.360 ;
        RECT 11.170 1.060 11.380 2.450 ;
        RECT 11.140 1.980 11.380 2.450 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.160 1.060 10.330 1.470 ;
        RECT 10.160 2.000 10.330 2.300 ;
        RECT 10.160 1.290 10.560 1.470 ;
        RECT 10.350 1.290 10.560 2.235 ;
        RECT 10.160 2.000 10.560 2.235 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 2.485 2.270 3.000 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.455 1.605 3.075 1.950 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.960 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 -0.300 0.890 0.800 ;
        RECT 2.825 -0.300 3.125 0.595 ;
        RECT 3.795 -0.300 4.095 0.595 ;
        RECT 6.285 -0.300 6.585 0.595 ;
        RECT 7.400 -0.300 7.700 0.565 ;
        RECT 9.125 -0.300 9.425 0.560 ;
        RECT 10.525 -0.300 10.825 0.745 ;
        RECT 0.000 -0.300 11.480 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 3.255 1.475 3.690 1.950 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.780 1.330 1.190 1.820 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 2.540 0.890 3.990 ;
        RECT 2.470 2.620 2.640 3.990 ;
        RECT 3.585 2.830 3.755 3.990 ;
        RECT 6.470 3.160 7.450 3.990 ;
        RECT 9.005 2.895 9.305 3.990 ;
        RECT 10.525 2.830 10.825 3.990 ;
        RECT 0.000 3.390 11.480 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.980 0.340 2.280 ;
        RECT 0.170 2.110 1.275 2.280 ;
        RECT 1.105 0.710 1.275 1.150 ;
        RECT 0.170 0.980 1.275 1.150 ;
        RECT 1.105 2.110 1.275 2.645 ;
        RECT 1.105 2.475 1.510 2.645 ;
        RECT 1.340 2.475 1.510 2.775 ;
        RECT 1.105 0.710 2.015 0.880 ;
        RECT 2.040 1.980 2.210 2.300 ;
        RECT 2.040 2.130 3.255 2.300 ;
        RECT 1.550 1.060 1.720 2.280 ;
        RECT 1.520 1.980 1.720 2.280 ;
        RECT 2.410 0.775 2.580 1.230 ;
        RECT 1.550 1.060 2.580 1.230 ;
        RECT 2.410 0.775 4.980 0.945 ;
        RECT 4.810 0.670 4.980 2.280 ;
        RECT 5.510 0.900 5.680 2.280 ;
        RECT 6.655 1.675 6.965 1.865 ;
        RECT 5.510 1.695 6.965 1.865 ;
        RECT 6.165 1.325 6.465 1.515 ;
        RECT 6.920 0.610 7.200 1.495 ;
        RECT 6.165 1.325 7.635 1.495 ;
        RECT 7.465 1.325 7.635 2.215 ;
        RECT 6.825 2.045 7.635 2.215 ;
        RECT 3.005 2.480 3.175 3.130 ;
        RECT 3.215 1.125 4.045 1.295 ;
        RECT 3.005 2.480 4.105 2.650 ;
        RECT 3.875 1.125 4.045 2.650 ;
        RECT 3.935 1.525 4.105 2.980 ;
        RECT 3.875 1.525 4.170 1.825 ;
        RECT 3.935 2.810 8.105 2.980 ;
        RECT 4.255 1.125 4.555 1.295 ;
        RECT 4.290 1.980 4.555 2.280 ;
        RECT 4.385 1.125 4.555 2.630 ;
        RECT 5.160 0.535 5.330 2.630 ;
        RECT 5.160 0.535 5.955 0.705 ;
        RECT 7.815 1.425 7.985 2.630 ;
        RECT 7.880 0.500 8.050 1.595 ;
        RECT 7.815 1.425 8.050 1.595 ;
        RECT 7.880 0.500 8.265 0.670 ;
        RECT 4.385 2.460 8.685 2.630 ;
        RECT 8.875 1.450 9.820 1.620 ;
        RECT 9.620 1.450 9.790 2.280 ;
        RECT 9.650 0.875 9.820 1.820 ;
        RECT 9.620 1.450 9.820 1.820 ;
        RECT 9.620 1.650 10.170 1.820 ;
        RECT 8.240 0.875 8.410 2.215 ;
        RECT 8.175 2.045 9.235 2.215 ;
        RECT 9.065 2.045 9.235 2.650 ;
        RECT 10.790 1.520 10.960 2.650 ;
        RECT 9.065 2.480 10.960 2.650 ;
        RECT 10.790 1.520 10.990 1.820 ;
  END 
END FFSDCRHDLXHT

MACRO FFSDCRHD2XHT
  CLASS  CORE ;
  FOREIGN FFSDCRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.120 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 12.260 0.720 12.430 2.960 ;
        RECT 12.260 1.270 12.610 1.640 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.170 0.720 11.380 2.280 ;
        RECT 11.170 0.720 11.390 1.360 ;
        RECT 11.170 1.980 11.390 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.935 2.485 2.390 2.950 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.455 1.590 3.075 1.950 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.960 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 -0.300 0.890 0.800 ;
        RECT 2.865 -0.300 3.165 0.595 ;
        RECT 4.025 -0.300 4.325 0.595 ;
        RECT 6.585 -0.300 6.885 0.595 ;
        RECT 7.600 -0.300 7.900 0.715 ;
        RECT 9.345 -0.300 9.515 0.780 ;
        RECT 10.700 -0.300 10.870 1.120 ;
        RECT 11.675 -0.300 11.975 1.055 ;
        RECT 12.715 -0.300 13.015 1.055 ;
        RECT 0.000 -0.300 13.120 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 3.550 1.525 4.040 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.780 1.330 1.190 1.820 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 2.650 0.890 3.990 ;
        RECT 2.590 2.845 2.760 3.990 ;
        RECT 3.935 2.675 4.105 3.990 ;
        RECT 6.730 3.160 7.030 3.990 ;
        RECT 7.570 3.095 7.870 3.990 ;
        RECT 9.465 2.805 9.635 3.990 ;
        RECT 10.635 2.975 10.935 3.990 ;
        RECT 11.675 2.975 11.975 3.990 ;
        RECT 12.715 2.295 13.015 3.990 ;
        RECT 0.000 3.390 13.120 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.980 0.340 2.280 ;
        RECT 0.170 2.110 1.275 2.280 ;
        RECT 1.105 0.555 1.275 1.150 ;
        RECT 0.170 0.980 1.275 1.150 ;
        RECT 1.105 2.110 1.275 2.885 ;
        RECT 1.105 2.715 1.575 2.885 ;
        RECT 1.105 0.555 2.055 0.725 ;
        RECT 1.975 2.130 3.255 2.300 ;
        RECT 1.520 1.060 1.690 2.280 ;
        RECT 2.455 0.775 2.625 1.230 ;
        RECT 1.520 1.060 2.625 1.230 ;
        RECT 2.455 0.775 5.320 0.945 ;
        RECT 5.150 0.775 5.320 2.280 ;
        RECT 5.850 0.910 6.020 2.280 ;
        RECT 6.955 1.675 7.255 1.865 ;
        RECT 5.850 1.695 7.255 1.865 ;
        RECT 6.445 1.325 6.745 1.515 ;
        RECT 7.200 0.910 7.370 1.495 ;
        RECT 6.445 1.325 8.015 1.495 ;
        RECT 7.845 1.325 8.015 2.215 ;
        RECT 7.170 2.045 8.015 2.215 ;
        RECT 3.475 1.125 4.395 1.295 ;
        RECT 3.475 2.190 4.455 2.360 ;
        RECT 4.225 1.125 4.395 2.360 ;
        RECT 4.285 1.525 4.455 3.050 ;
        RECT 4.225 1.525 4.520 1.825 ;
        RECT 4.285 2.880 6.330 3.050 ;
        RECT 6.555 2.745 7.965 2.915 ;
        RECT 8.025 2.745 8.055 2.975 ;
        RECT 8.115 2.805 8.555 2.975 ;
        RECT 8.385 2.805 8.555 3.210 ;
        RECT 8.385 3.040 9.070 3.210 ;
        RECT 8.055 2.755 8.065 2.975 ;
        RECT 8.065 2.765 8.075 2.975 ;
        RECT 8.075 2.775 8.085 2.975 ;
        RECT 8.085 2.785 8.095 2.975 ;
        RECT 8.095 2.795 8.105 2.975 ;
        RECT 8.105 2.805 8.115 2.975 ;
        RECT 7.965 2.745 7.975 2.915 ;
        RECT 7.975 2.745 7.985 2.925 ;
        RECT 7.985 2.745 7.995 2.935 ;
        RECT 7.995 2.745 8.005 2.945 ;
        RECT 8.005 2.745 8.015 2.955 ;
        RECT 8.015 2.745 8.025 2.965 ;
        RECT 6.465 2.745 6.475 2.995 ;
        RECT 6.475 2.745 6.485 2.985 ;
        RECT 6.485 2.745 6.495 2.975 ;
        RECT 6.495 2.745 6.505 2.965 ;
        RECT 6.505 2.745 6.515 2.955 ;
        RECT 6.515 2.745 6.525 2.945 ;
        RECT 6.525 2.745 6.535 2.935 ;
        RECT 6.535 2.745 6.545 2.925 ;
        RECT 6.545 2.745 6.555 2.915 ;
        RECT 6.420 2.790 6.430 3.040 ;
        RECT 6.430 2.780 6.440 3.030 ;
        RECT 6.440 2.770 6.450 3.020 ;
        RECT 6.450 2.760 6.460 3.010 ;
        RECT 6.460 2.750 6.466 3.004 ;
        RECT 6.330 2.880 6.340 3.050 ;
        RECT 6.340 2.870 6.350 3.050 ;
        RECT 6.350 2.860 6.360 3.050 ;
        RECT 6.360 2.850 6.370 3.050 ;
        RECT 6.370 2.840 6.380 3.050 ;
        RECT 6.380 2.830 6.390 3.050 ;
        RECT 6.390 2.820 6.400 3.050 ;
        RECT 6.400 2.810 6.410 3.050 ;
        RECT 6.410 2.800 6.420 3.050 ;
        RECT 4.575 1.125 4.895 1.295 ;
        RECT 4.725 1.125 4.895 2.635 ;
        RECT 4.640 1.980 4.895 2.635 ;
        RECT 5.500 0.535 5.670 2.700 ;
        RECT 5.415 2.465 5.715 2.700 ;
        RECT 6.165 2.435 6.255 2.635 ;
        RECT 6.155 2.445 9.005 2.565 ;
        RECT 6.175 2.425 6.255 2.635 ;
        RECT 6.145 2.455 9.005 2.565 ;
        RECT 4.640 2.465 6.255 2.635 ;
        RECT 5.500 0.535 6.265 0.705 ;
        RECT 4.640 2.465 6.265 2.625 ;
        RECT 4.640 2.465 6.275 2.615 ;
        RECT 4.640 2.465 6.285 2.605 ;
        RECT 4.640 2.465 6.295 2.595 ;
        RECT 4.640 2.465 6.305 2.585 ;
        RECT 4.640 2.465 6.315 2.575 ;
        RECT 6.205 2.395 8.395 2.565 ;
        RECT 6.195 2.405 8.395 2.565 ;
        RECT 8.225 0.710 8.395 2.590 ;
        RECT 6.185 2.415 8.395 2.565 ;
        RECT 8.225 2.420 9.005 2.590 ;
        RECT 8.225 0.710 9.110 0.880 ;
        RECT 8.835 2.420 9.005 2.795 ;
        RECT 8.940 0.710 9.110 1.140 ;
        RECT 9.695 0.480 9.865 1.140 ;
        RECT 8.940 0.970 9.865 1.140 ;
        RECT 9.695 0.480 10.520 0.650 ;
        RECT 9.260 1.675 10.215 1.845 ;
        RECT 10.045 1.060 10.215 2.280 ;
        RECT 10.045 1.625 10.990 1.795 ;
        RECT 8.585 1.060 8.755 2.240 ;
        RECT 8.575 2.070 9.865 2.240 ;
        RECT 9.695 2.070 9.865 2.630 ;
        RECT 9.835 2.460 10.005 3.190 ;
        RECT 11.910 1.570 12.080 2.630 ;
        RECT 9.695 2.460 12.080 2.630 ;
  END 
END FFSDCRHD2XHT

MACRO FFSDCRHD1XHT
  CLASS  CORE ;
  FOREIGN FFSDCRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.890 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.550 0.720 11.790 1.360 ;
        RECT 11.620 0.720 11.790 2.960 ;
        RECT 11.550 1.980 11.790 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.510 0.720 10.680 1.445 ;
        RECT 10.510 2.000 10.680 2.300 ;
        RECT 10.510 1.265 10.970 1.445 ;
        RECT 10.760 1.265 10.970 2.235 ;
        RECT 10.510 2.000 10.970 2.235 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.935 2.485 2.390 2.950 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.455 1.590 3.075 1.950 ;
    END
  END RN
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.960 ;
    END
  END TE
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 -0.300 0.890 0.800 ;
        RECT 2.865 -0.300 3.165 0.595 ;
        RECT 4.035 -0.300 4.335 0.595 ;
        RECT 6.635 -0.300 6.935 0.595 ;
        RECT 7.575 -0.300 7.875 0.615 ;
        RECT 9.465 -0.300 9.765 0.630 ;
        RECT 10.965 -0.300 11.265 1.055 ;
        RECT 0.000 -0.300 11.890 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 3.560 1.525 4.050 2.010 ;
    END
  END CK
  PIN TI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.780 1.330 1.190 1.820 ;
    END
  END TI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 2.680 0.890 3.990 ;
        RECT 2.590 2.845 2.760 3.990 ;
        RECT 3.945 2.675 4.115 3.990 ;
        RECT 6.810 3.160 7.790 3.990 ;
        RECT 9.420 2.850 9.590 3.990 ;
        RECT 10.965 2.975 11.265 3.990 ;
        RECT 0.000 3.390 11.890 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.980 0.340 2.280 ;
        RECT 0.170 2.110 1.275 2.280 ;
        RECT 1.105 0.555 1.275 1.150 ;
        RECT 0.170 0.980 1.275 1.150 ;
        RECT 1.105 2.110 1.275 2.885 ;
        RECT 1.105 2.715 1.575 2.885 ;
        RECT 1.105 0.555 2.055 0.725 ;
        RECT 1.975 2.130 3.255 2.300 ;
        RECT 1.520 1.060 1.690 2.280 ;
        RECT 2.455 0.775 2.625 1.230 ;
        RECT 1.520 1.060 2.625 1.230 ;
        RECT 2.455 0.775 5.330 0.945 ;
        RECT 5.160 0.775 5.330 2.280 ;
        RECT 5.860 0.900 6.030 2.280 ;
        RECT 7.005 1.675 7.315 1.865 ;
        RECT 5.860 1.695 7.315 1.865 ;
        RECT 6.505 1.325 6.805 1.515 ;
        RECT 7.250 0.910 7.420 1.495 ;
        RECT 6.505 1.325 8.020 1.495 ;
        RECT 7.850 1.325 8.020 2.215 ;
        RECT 7.185 2.045 8.020 2.215 ;
        RECT 3.485 1.125 4.405 1.295 ;
        RECT 3.465 2.190 4.465 2.360 ;
        RECT 4.235 1.125 4.405 2.360 ;
        RECT 4.295 1.525 4.465 2.980 ;
        RECT 4.235 1.525 4.530 1.825 ;
        RECT 4.295 2.810 8.565 2.980 ;
        RECT 4.585 1.125 4.905 1.295 ;
        RECT 4.650 1.980 4.905 2.280 ;
        RECT 4.735 1.125 4.905 2.630 ;
        RECT 5.510 0.535 5.680 2.630 ;
        RECT 5.510 0.535 6.305 0.705 ;
        RECT 8.200 0.480 8.370 2.630 ;
        RECT 8.200 0.480 8.565 0.650 ;
        RECT 8.200 2.440 9.010 2.630 ;
        RECT 4.735 2.460 9.010 2.630 ;
        RECT 8.840 2.440 9.010 2.770 ;
        RECT 9.225 1.570 10.330 1.740 ;
        RECT 10.000 0.945 10.170 1.740 ;
        RECT 10.160 1.570 10.330 2.215 ;
        RECT 9.905 2.045 10.330 2.215 ;
        RECT 10.160 1.650 10.555 1.820 ;
        RECT 8.610 0.945 8.780 2.215 ;
        RECT 8.555 2.045 9.725 2.215 ;
        RECT 9.555 2.045 9.725 2.650 ;
        RECT 9.790 2.480 9.960 2.780 ;
        RECT 11.200 1.520 11.370 2.650 ;
        RECT 9.555 2.480 11.370 2.650 ;
        RECT 11.200 1.520 11.390 1.820 ;
  END 
END FFSDCRHD1XHT

MACRO FFEDQHDMXHT
  CLASS  CORE ;
  FOREIGN FFEDQHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.320 1.060 10.560 1.360 ;
        RECT 10.350 1.060 10.560 2.445 ;
        RECT 10.320 1.980 10.560 2.445 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 1.325 1.220 2.005 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.595 0.620 2.015 ;
        RECT 0.385 2.665 2.215 2.835 ;
        RECT 1.915 2.665 2.215 2.900 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.755 -0.300 1.055 0.795 ;
        RECT 2.610 -0.300 3.590 0.520 ;
        RECT 6.105 -0.300 6.405 0.525 ;
        RECT 7.065 -0.300 7.365 0.565 ;
        RECT 8.885 -0.300 9.185 0.470 ;
        RECT 9.705 -0.300 10.005 0.470 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.970 1.525 3.485 2.015 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.735 3.035 1.035 3.990 ;
        RECT 2.685 2.905 3.665 3.990 ;
        RECT 6.050 3.160 7.030 3.990 ;
        RECT 8.690 2.920 8.990 3.990 ;
        RECT 9.705 2.920 10.005 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.205 0.975 1.590 1.145 ;
        RECT 1.420 0.975 1.590 2.430 ;
        RECT 0.205 2.260 1.590 2.430 ;
        RECT 1.420 1.705 1.700 2.005 ;
        RECT 3.015 1.125 3.845 1.295 ;
        RECT 3.665 1.125 3.845 2.365 ;
        RECT 3.045 2.195 3.845 2.365 ;
        RECT 3.665 1.525 4.000 1.825 ;
        RECT 4.055 1.065 4.355 1.235 ;
        RECT 4.180 1.065 4.350 2.280 ;
        RECT 4.170 1.980 4.350 2.280 ;
        RECT 4.180 1.065 4.355 1.840 ;
        RECT 4.180 1.540 4.480 1.840 ;
        RECT 1.770 0.945 2.110 1.245 ;
        RECT 1.940 0.945 2.110 2.485 ;
        RECT 1.780 2.185 2.110 2.485 ;
        RECT 1.780 2.305 2.800 2.485 ;
        RECT 2.630 2.305 2.800 2.725 ;
        RECT 4.660 1.065 4.830 2.725 ;
        RECT 2.630 2.545 4.830 2.725 ;
        RECT 4.575 1.065 4.875 1.235 ;
        RECT 5.165 1.060 5.335 2.280 ;
        RECT 5.165 1.060 5.360 1.930 ;
        RECT 5.155 1.060 5.455 1.230 ;
        RECT 6.355 1.675 6.655 1.930 ;
        RECT 5.165 1.760 6.655 1.930 ;
        RECT 5.875 1.325 6.175 1.540 ;
        RECT 6.565 1.125 6.865 1.495 ;
        RECT 5.875 1.325 7.320 1.495 ;
        RECT 7.150 1.325 7.320 2.280 ;
        RECT 6.480 2.110 7.320 2.280 ;
        RECT 5.535 2.810 5.705 3.145 ;
        RECT 3.925 2.975 5.705 3.145 ;
        RECT 5.535 2.810 7.240 2.980 ;
        RECT 7.485 2.975 7.850 3.145 ;
        RECT 7.405 2.905 7.415 3.145 ;
        RECT 7.415 2.915 7.425 3.145 ;
        RECT 7.425 2.925 7.435 3.145 ;
        RECT 7.435 2.935 7.445 3.145 ;
        RECT 7.445 2.945 7.455 3.145 ;
        RECT 7.455 2.955 7.465 3.145 ;
        RECT 7.465 2.965 7.475 3.145 ;
        RECT 7.475 2.975 7.485 3.145 ;
        RECT 7.320 2.820 7.330 3.060 ;
        RECT 7.330 2.830 7.340 3.070 ;
        RECT 7.340 2.840 7.350 3.080 ;
        RECT 7.350 2.850 7.360 3.090 ;
        RECT 7.360 2.860 7.370 3.100 ;
        RECT 7.370 2.870 7.380 3.110 ;
        RECT 7.380 2.880 7.390 3.120 ;
        RECT 7.390 2.890 7.400 3.130 ;
        RECT 7.400 2.895 7.406 3.139 ;
        RECT 7.240 2.810 7.250 2.980 ;
        RECT 7.250 2.810 7.260 2.990 ;
        RECT 7.260 2.810 7.270 3.000 ;
        RECT 7.270 2.810 7.280 3.010 ;
        RECT 7.280 2.810 7.290 3.020 ;
        RECT 7.290 2.810 7.300 3.030 ;
        RECT 7.300 2.810 7.310 3.040 ;
        RECT 7.310 2.810 7.320 3.050 ;
        RECT 5.035 2.460 5.205 2.770 ;
        RECT 7.500 1.310 7.540 2.630 ;
        RECT 5.035 2.460 7.540 2.630 ;
        RECT 7.650 1.310 7.670 2.740 ;
        RECT 7.650 1.310 7.900 1.480 ;
        RECT 7.780 2.570 8.305 2.740 ;
        RECT 8.135 2.570 8.305 2.870 ;
        RECT 7.670 2.470 7.680 2.740 ;
        RECT 7.680 2.480 7.690 2.740 ;
        RECT 7.690 2.490 7.700 2.740 ;
        RECT 7.700 2.500 7.710 2.740 ;
        RECT 7.710 2.510 7.720 2.740 ;
        RECT 7.720 2.520 7.730 2.740 ;
        RECT 7.730 2.530 7.740 2.740 ;
        RECT 7.740 2.540 7.750 2.740 ;
        RECT 7.750 2.550 7.760 2.740 ;
        RECT 7.760 2.560 7.770 2.740 ;
        RECT 7.770 2.570 7.780 2.740 ;
        RECT 7.540 1.310 7.550 2.630 ;
        RECT 7.550 1.310 7.560 2.640 ;
        RECT 7.560 1.310 7.570 2.650 ;
        RECT 7.570 1.310 7.580 2.660 ;
        RECT 7.580 1.310 7.590 2.670 ;
        RECT 7.590 1.310 7.600 2.680 ;
        RECT 7.600 1.310 7.610 2.690 ;
        RECT 7.610 1.310 7.620 2.700 ;
        RECT 7.620 1.310 7.630 2.710 ;
        RECT 7.630 1.310 7.640 2.720 ;
        RECT 7.640 1.310 7.650 2.730 ;
        RECT 2.510 0.700 2.680 1.825 ;
        RECT 2.510 0.700 3.205 0.890 ;
        RECT 4.405 0.590 4.585 0.885 ;
        RECT 2.510 0.700 4.585 0.885 ;
        RECT 4.405 0.590 5.765 0.760 ;
        RECT 5.595 0.590 5.765 0.945 ;
        RECT 7.650 0.480 7.820 0.945 ;
        RECT 5.595 0.765 7.820 0.945 ;
        RECT 7.650 0.480 8.560 0.665 ;
        RECT 8.655 1.355 8.785 1.525 ;
        RECT 8.810 0.650 8.955 1.525 ;
        RECT 8.810 0.650 9.670 0.820 ;
        RECT 9.380 0.650 9.670 1.175 ;
        RECT 9.500 0.650 9.670 2.390 ;
        RECT 9.240 2.220 9.670 2.390 ;
        RECT 8.785 0.635 8.795 1.525 ;
        RECT 8.795 0.645 8.805 1.525 ;
        RECT 8.805 0.650 8.811 1.524 ;
        RECT 8.715 0.565 8.725 0.819 ;
        RECT 8.725 0.575 8.735 0.819 ;
        RECT 8.735 0.585 8.745 0.819 ;
        RECT 8.745 0.595 8.755 0.819 ;
        RECT 8.755 0.605 8.765 0.819 ;
        RECT 8.765 0.615 8.775 0.819 ;
        RECT 8.775 0.625 8.785 0.819 ;
        RECT 8.640 0.490 8.650 0.744 ;
        RECT 8.650 0.500 8.660 0.754 ;
        RECT 8.660 0.510 8.670 0.764 ;
        RECT 8.670 0.520 8.680 0.774 ;
        RECT 8.680 0.530 8.690 0.784 ;
        RECT 8.690 0.540 8.700 0.794 ;
        RECT 8.700 0.550 8.710 0.804 ;
        RECT 8.710 0.555 8.716 0.815 ;
        RECT 8.560 0.480 8.570 0.664 ;
        RECT 8.570 0.480 8.580 0.674 ;
        RECT 8.580 0.480 8.590 0.684 ;
        RECT 8.590 0.480 8.600 0.694 ;
        RECT 8.600 0.480 8.610 0.704 ;
        RECT 8.610 0.480 8.620 0.714 ;
        RECT 8.620 0.480 8.630 0.724 ;
        RECT 8.630 0.480 8.640 0.734 ;
        RECT 8.000 0.845 8.265 1.145 ;
        RECT 8.095 0.845 8.265 2.390 ;
        RECT 7.890 2.220 8.265 2.390 ;
        RECT 8.095 1.740 9.295 1.910 ;
        RECT 8.890 1.740 9.060 2.740 ;
        RECT 8.890 1.740 9.295 2.040 ;
        RECT 9.970 1.520 10.140 2.740 ;
        RECT 8.890 2.570 10.140 2.740 ;
        RECT 9.970 1.520 10.160 1.820 ;
  END 
END FFEDQHDMXHT

MACRO FFEDQHDLXHT
  CLASS  CORE ;
  FOREIGN FFEDQHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.000 1.040 10.560 1.340 ;
        RECT 10.350 1.040 10.560 2.460 ;
        RECT 10.320 2.100 10.560 2.460 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 1.325 1.195 2.005 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.550 0.565 2.015 ;
        RECT 0.330 2.665 2.160 2.835 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 -0.300 1.020 0.795 ;
        RECT 2.510 -0.300 2.810 0.520 ;
        RECT 3.480 -0.300 3.780 0.520 ;
        RECT 6.010 -0.300 6.310 0.585 ;
        RECT 6.980 -0.300 7.280 0.565 ;
        RECT 8.880 -0.300 9.180 0.470 ;
        RECT 9.935 -0.300 10.235 0.755 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.970 1.525 3.555 2.015 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 3.015 1.020 3.990 ;
        RECT 2.705 2.905 3.685 3.990 ;
        RECT 6.215 3.160 7.195 3.990 ;
        RECT 8.880 2.745 9.180 3.990 ;
        RECT 9.705 2.745 10.005 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.150 2.205 0.450 2.430 ;
        RECT 0.150 0.975 1.545 1.145 ;
        RECT 1.375 0.975 1.545 2.375 ;
        RECT 0.150 2.205 1.545 2.375 ;
        RECT 1.375 1.705 1.710 1.955 ;
        RECT 3.020 1.125 3.905 1.295 ;
        RECT 3.735 1.125 3.905 2.365 ;
        RECT 2.990 2.195 3.905 2.365 ;
        RECT 3.735 1.525 3.970 1.825 ;
        RECT 4.085 1.125 4.385 1.295 ;
        RECT 4.150 1.125 4.320 2.280 ;
        RECT 4.150 1.125 4.385 1.850 ;
        RECT 4.150 1.550 4.450 1.850 ;
        RECT 1.745 1.045 2.060 1.345 ;
        RECT 1.890 1.045 2.060 2.485 ;
        RECT 1.725 2.135 2.060 2.485 ;
        RECT 1.725 2.305 2.775 2.485 ;
        RECT 2.605 2.305 2.775 2.725 ;
        RECT 4.665 1.060 4.845 2.725 ;
        RECT 2.605 2.545 4.845 2.725 ;
        RECT 4.595 1.060 4.895 1.230 ;
        RECT 5.245 1.060 5.415 2.280 ;
        RECT 5.180 1.060 5.480 1.230 ;
        RECT 6.380 1.675 6.680 1.930 ;
        RECT 5.245 1.760 6.680 1.930 ;
        RECT 5.900 1.325 6.200 1.540 ;
        RECT 6.590 1.125 6.890 1.495 ;
        RECT 5.900 1.325 7.400 1.495 ;
        RECT 7.230 1.325 7.400 2.280 ;
        RECT 6.590 2.110 7.400 2.280 ;
        RECT 5.615 2.810 5.785 3.145 ;
        RECT 3.875 2.975 5.785 3.145 ;
        RECT 5.615 2.810 7.860 2.980 ;
        RECT 5.035 2.460 5.205 2.770 ;
        RECT 7.580 1.310 7.750 2.630 ;
        RECT 7.580 1.310 7.980 1.480 ;
        RECT 5.035 2.460 8.375 2.630 ;
        RECT 8.205 2.460 8.375 2.865 ;
        RECT 2.455 0.700 2.625 1.825 ;
        RECT 5.660 0.700 5.830 0.945 ;
        RECT 2.455 0.700 5.830 0.880 ;
        RECT 7.500 0.575 7.670 0.945 ;
        RECT 5.660 0.765 7.670 0.945 ;
        RECT 7.500 0.575 8.730 0.760 ;
        RECT 8.560 0.575 8.730 1.480 ;
        RECT 8.560 1.310 9.745 1.480 ;
        RECT 9.415 0.875 9.585 1.480 ;
        RECT 9.575 1.310 9.745 2.215 ;
        RECT 9.310 2.045 9.745 2.215 ;
        RECT 7.930 0.940 8.330 1.110 ;
        RECT 8.160 0.940 8.330 2.215 ;
        RECT 7.930 2.045 8.330 2.215 ;
        RECT 8.960 1.675 9.130 2.565 ;
        RECT 8.160 1.675 9.395 1.845 ;
        RECT 9.970 1.610 10.140 2.565 ;
        RECT 8.960 2.395 10.140 2.565 ;
        RECT 9.970 1.610 10.160 1.910 ;
  END 
END FFEDQHDLXHT

MACRO FFEDQHD2XHT
  CLASS  CORE ;
  FOREIGN FFEDQHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.480 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.620 0.720 10.790 2.960 ;
        RECT 10.620 2.050 10.975 2.425 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.875 1.265 1.130 2.015 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.600 0.605 2.015 ;
        RECT 0.285 2.665 2.115 2.835 ;
        RECT 1.815 2.665 2.115 3.180 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.675 -0.300 0.975 0.710 ;
        RECT 2.435 -0.300 2.735 0.520 ;
        RECT 3.495 -0.300 3.795 0.520 ;
        RECT 5.860 -0.300 6.160 0.525 ;
        RECT 6.850 -0.300 7.150 0.565 ;
        RECT 9.020 -0.300 9.320 0.445 ;
        RECT 10.100 -0.300 10.270 1.120 ;
        RECT 11.075 -0.300 11.375 1.055 ;
        RECT 0.000 -0.300 11.480 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.870 1.525 3.425 1.950 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.635 3.035 0.935 3.990 ;
        RECT 2.585 2.840 3.565 3.990 ;
        RECT 5.980 3.160 6.280 3.990 ;
        RECT 6.750 3.160 7.050 3.990 ;
        RECT 8.975 2.780 9.275 3.990 ;
        RECT 10.035 2.975 10.335 3.990 ;
        RECT 11.075 2.635 11.375 3.990 ;
        RECT 0.000 3.390 11.480 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.915 0.405 1.145 ;
        RECT 0.105 2.205 0.405 2.430 ;
        RECT 0.105 0.915 1.500 1.085 ;
        RECT 1.330 0.915 1.500 2.375 ;
        RECT 0.105 2.205 1.500 2.375 ;
        RECT 1.330 1.705 1.600 2.005 ;
        RECT 2.945 1.125 3.775 1.295 ;
        RECT 3.605 1.125 3.775 2.300 ;
        RECT 2.945 2.130 3.775 2.300 ;
        RECT 3.605 1.525 3.840 1.825 ;
        RECT 3.955 1.065 4.255 1.235 ;
        RECT 4.020 1.065 4.190 2.280 ;
        RECT 4.020 1.065 4.255 1.850 ;
        RECT 4.020 1.550 4.320 1.850 ;
        RECT 1.680 0.945 2.010 1.245 ;
        RECT 1.840 0.945 2.010 2.485 ;
        RECT 1.680 2.185 2.010 2.485 ;
        RECT 2.520 2.305 2.690 2.660 ;
        RECT 1.680 2.305 2.690 2.485 ;
        RECT 4.535 1.980 4.705 2.660 ;
        RECT 2.520 2.480 4.705 2.660 ;
        RECT 4.545 1.060 4.715 2.380 ;
        RECT 4.535 1.980 4.715 2.380 ;
        RECT 4.465 1.060 4.765 1.230 ;
        RECT 5.095 1.060 5.265 2.280 ;
        RECT 5.030 1.060 5.330 1.230 ;
        RECT 6.230 1.675 6.530 1.930 ;
        RECT 5.095 1.760 6.530 1.930 ;
        RECT 5.750 1.325 6.050 1.540 ;
        RECT 6.440 1.125 6.740 1.495 ;
        RECT 5.750 1.325 7.285 1.495 ;
        RECT 7.115 1.325 7.285 2.280 ;
        RECT 6.410 2.110 7.285 2.280 ;
        RECT 4.885 2.460 5.055 2.770 ;
        RECT 4.885 2.460 8.295 2.630 ;
        RECT 8.125 2.460 8.295 2.795 ;
        RECT 3.745 2.950 4.045 3.185 ;
        RECT 5.465 2.810 5.635 3.120 ;
        RECT 3.745 2.950 5.635 3.120 ;
        RECT 5.465 2.810 7.850 2.980 ;
        RECT 7.680 2.810 7.850 3.210 ;
        RECT 8.220 1.350 8.665 1.520 ;
        RECT 8.485 1.350 8.665 3.210 ;
        RECT 7.680 3.040 8.665 3.210 ;
        RECT 2.410 0.700 2.580 1.825 ;
        RECT 2.410 0.700 5.650 0.880 ;
        RECT 5.715 0.700 5.775 0.945 ;
        RECT 5.840 0.765 7.280 0.945 ;
        RECT 8.540 0.580 8.840 0.820 ;
        RECT 7.480 0.635 8.840 0.820 ;
        RECT 7.480 0.650 9.695 0.820 ;
        RECT 9.525 0.650 9.695 1.295 ;
        RECT 9.525 1.125 9.920 1.295 ;
        RECT 9.750 1.125 9.920 2.240 ;
        RECT 9.525 2.070 9.920 2.240 ;
        RECT 7.410 0.635 7.420 0.879 ;
        RECT 7.420 0.635 7.430 0.869 ;
        RECT 7.430 0.635 7.440 0.859 ;
        RECT 7.440 0.635 7.450 0.849 ;
        RECT 7.450 0.635 7.460 0.839 ;
        RECT 7.460 0.635 7.470 0.829 ;
        RECT 7.470 0.635 7.480 0.819 ;
        RECT 7.355 0.690 7.365 0.934 ;
        RECT 7.365 0.680 7.375 0.924 ;
        RECT 7.375 0.670 7.385 0.914 ;
        RECT 7.385 0.660 7.395 0.904 ;
        RECT 7.395 0.650 7.405 0.894 ;
        RECT 7.405 0.640 7.411 0.890 ;
        RECT 7.280 0.765 7.290 0.945 ;
        RECT 7.290 0.755 7.300 0.945 ;
        RECT 7.300 0.745 7.310 0.945 ;
        RECT 7.310 0.735 7.320 0.945 ;
        RECT 7.320 0.725 7.330 0.945 ;
        RECT 7.330 0.715 7.340 0.945 ;
        RECT 7.340 0.705 7.350 0.945 ;
        RECT 7.350 0.695 7.356 0.945 ;
        RECT 5.775 0.710 5.785 0.944 ;
        RECT 5.785 0.720 5.795 0.944 ;
        RECT 5.795 0.730 5.805 0.944 ;
        RECT 5.805 0.740 5.815 0.944 ;
        RECT 5.815 0.750 5.825 0.944 ;
        RECT 5.825 0.760 5.835 0.944 ;
        RECT 5.835 0.765 5.841 0.945 ;
        RECT 5.650 0.700 5.660 0.880 ;
        RECT 5.660 0.700 5.670 0.890 ;
        RECT 5.670 0.700 5.680 0.900 ;
        RECT 5.680 0.700 5.690 0.910 ;
        RECT 5.690 0.700 5.700 0.920 ;
        RECT 5.700 0.700 5.710 0.930 ;
        RECT 5.710 0.700 5.716 0.940 ;
        RECT 7.555 1.000 7.735 2.240 ;
        RECT 7.555 2.070 8.020 2.240 ;
        RECT 7.555 1.000 9.250 1.170 ;
        RECT 9.080 1.000 9.250 2.600 ;
        RECT 9.080 1.590 9.570 1.760 ;
        RECT 10.100 1.540 10.270 2.600 ;
        RECT 9.080 2.430 10.270 2.600 ;
        RECT 10.100 1.540 10.440 1.840 ;
  END 
END FFEDQHD2XHT

MACRO FFDSHQHD3XHT
  CLASS  CORE ;
  FOREIGN FFDSHQHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.530 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.540 0.720 11.840 1.495 ;
        RECT 11.705 2.070 11.875 3.210 ;
        RECT 11.585 2.230 11.875 3.210 ;
        RECT 11.705 2.070 12.880 2.390 ;
        RECT 11.585 2.230 12.880 2.390 ;
        RECT 12.580 0.720 12.880 1.495 ;
        RECT 11.540 1.255 12.880 1.495 ;
        RECT 12.640 0.720 12.880 2.960 ;
        RECT 12.580 2.070 12.880 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.645 1.600 3.180 2.020 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 0.965 ;
        RECT 1.145 -0.300 1.445 0.965 ;
        RECT 2.715 -0.300 3.015 1.230 ;
        RECT 4.545 -0.300 4.780 1.130 ;
        RECT 6.555 -0.300 6.855 0.435 ;
        RECT 7.655 -0.300 7.955 0.435 ;
        RECT 10.110 -0.300 10.410 0.790 ;
        RECT 12.060 -0.300 12.360 1.055 ;
        RECT 13.100 -0.300 13.400 1.055 ;
        RECT 0.000 -0.300 13.530 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 1.090 1.230 1.665 1.700 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.975 0.615 9.865 0.650 ;
        RECT 4.975 0.615 8.265 0.715 ;
        RECT 4.975 1.250 5.380 1.260 ;
        RECT 5.145 0.545 5.315 1.415 ;
        RECT 5.145 1.250 5.380 1.415 ;
        RECT 5.210 0.545 5.315 1.665 ;
        RECT 4.975 0.545 5.315 1.260 ;
        RECT 5.210 1.250 5.380 1.665 ;
        RECT 5.210 1.495 6.000 1.665 ;
        RECT 6.175 0.545 6.345 0.785 ;
        RECT 4.975 0.545 6.345 0.715 ;
        RECT 8.115 0.530 8.265 0.785 ;
        RECT 8.115 0.530 9.865 0.650 ;
        RECT 8.245 0.480 8.265 0.785 ;
        RECT 6.175 0.615 8.265 0.785 ;
        RECT 8.245 0.480 8.370 0.700 ;
        RECT 4.975 0.615 8.370 0.700 ;
        RECT 9.165 0.480 9.245 0.670 ;
        RECT 8.245 0.480 9.245 0.650 ;
        RECT 9.165 0.500 9.865 0.670 ;
        RECT 9.695 0.500 9.865 1.140 ;
        RECT 10.590 0.655 10.760 1.140 ;
        RECT 9.695 0.970 10.760 1.140 ;
        RECT 10.590 0.655 11.110 0.825 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.280 0.860 3.990 ;
        RECT 1.675 2.965 1.975 3.990 ;
        RECT 2.685 2.965 2.985 3.990 ;
        RECT 4.625 3.095 4.925 3.990 ;
        RECT 5.815 3.095 6.455 3.990 ;
        RECT 7.345 3.155 7.645 3.990 ;
        RECT 10.110 2.845 10.410 3.990 ;
        RECT 11.030 2.745 11.330 3.990 ;
        RECT 12.115 2.570 12.360 3.990 ;
        RECT 13.100 2.295 13.400 3.990 ;
        RECT 0.000 3.390 13.530 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 2.280 0.340 3.175 ;
        RECT 0.105 3.005 0.405 3.175 ;
        RECT 1.665 0.795 2.020 1.050 ;
        RECT 1.850 0.795 2.020 1.700 ;
        RECT 1.850 1.400 2.080 1.700 ;
        RECT 3.720 2.145 3.825 2.445 ;
        RECT 4.055 1.445 4.810 1.615 ;
        RECT 4.860 1.445 4.910 1.865 ;
        RECT 4.910 1.455 4.920 1.865 ;
        RECT 4.920 1.465 4.930 1.865 ;
        RECT 4.930 1.475 4.940 1.865 ;
        RECT 4.940 1.485 4.950 1.865 ;
        RECT 4.950 1.495 4.960 1.865 ;
        RECT 4.960 1.505 4.970 1.865 ;
        RECT 4.970 1.515 4.980 1.865 ;
        RECT 4.980 1.525 4.990 1.865 ;
        RECT 4.990 1.535 5.000 1.865 ;
        RECT 5.000 1.545 5.010 1.865 ;
        RECT 5.010 1.555 5.020 1.865 ;
        RECT 5.020 1.565 5.030 1.865 ;
        RECT 4.810 1.445 4.820 1.615 ;
        RECT 4.820 1.445 4.830 1.625 ;
        RECT 4.830 1.445 4.840 1.635 ;
        RECT 4.840 1.445 4.850 1.645 ;
        RECT 4.850 1.445 4.860 1.655 ;
        RECT 4.025 1.425 4.035 1.615 ;
        RECT 4.035 1.435 4.045 1.615 ;
        RECT 4.045 1.445 4.055 1.615 ;
        RECT 3.890 1.290 3.900 2.434 ;
        RECT 3.900 1.300 3.910 2.424 ;
        RECT 3.910 1.310 3.920 2.414 ;
        RECT 3.920 1.320 3.930 2.404 ;
        RECT 3.930 1.330 3.940 2.394 ;
        RECT 3.940 1.340 3.950 2.384 ;
        RECT 3.950 1.350 3.960 2.374 ;
        RECT 3.960 1.360 3.970 2.364 ;
        RECT 3.970 1.370 3.980 2.354 ;
        RECT 3.980 1.380 3.990 2.344 ;
        RECT 3.990 1.390 4.000 2.334 ;
        RECT 4.000 1.400 4.010 2.324 ;
        RECT 4.010 1.410 4.020 2.314 ;
        RECT 4.020 1.415 4.026 2.309 ;
        RECT 3.855 1.255 3.865 2.445 ;
        RECT 3.865 1.265 3.875 2.445 ;
        RECT 3.875 1.275 3.885 2.445 ;
        RECT 3.885 1.280 3.891 2.444 ;
        RECT 3.840 1.240 3.850 1.480 ;
        RECT 3.850 1.245 3.856 1.489 ;
        RECT 3.825 2.145 3.835 2.445 ;
        RECT 3.835 2.135 3.845 2.445 ;
        RECT 3.845 2.125 3.855 2.445 ;
        RECT 3.670 0.995 3.680 1.309 ;
        RECT 3.680 0.995 3.690 1.319 ;
        RECT 3.690 0.995 3.700 1.329 ;
        RECT 3.700 0.995 3.710 1.339 ;
        RECT 3.710 0.995 3.720 1.349 ;
        RECT 3.720 0.995 3.730 1.359 ;
        RECT 3.730 0.995 3.740 1.369 ;
        RECT 3.740 0.995 3.750 1.379 ;
        RECT 3.750 0.995 3.760 1.389 ;
        RECT 3.760 0.995 3.770 1.399 ;
        RECT 3.770 0.995 3.780 1.409 ;
        RECT 3.780 0.995 3.790 1.419 ;
        RECT 3.790 0.995 3.800 1.429 ;
        RECT 3.800 0.995 3.810 1.439 ;
        RECT 3.810 0.995 3.820 1.449 ;
        RECT 3.820 0.995 3.830 1.459 ;
        RECT 3.830 0.995 3.840 1.469 ;
        RECT 4.315 1.795 4.615 2.215 ;
        RECT 5.810 1.845 5.980 2.215 ;
        RECT 4.315 2.045 5.980 2.215 ;
        RECT 5.810 1.845 6.130 2.015 ;
        RECT 5.525 0.965 6.220 1.135 ;
        RECT 6.390 1.495 7.400 1.665 ;
        RECT 6.220 0.965 6.230 1.995 ;
        RECT 6.230 0.965 6.240 1.985 ;
        RECT 6.240 0.965 6.250 1.975 ;
        RECT 6.250 0.965 6.260 1.965 ;
        RECT 6.260 0.965 6.270 1.955 ;
        RECT 6.270 0.965 6.280 1.945 ;
        RECT 6.280 0.965 6.290 1.935 ;
        RECT 6.290 0.965 6.300 1.925 ;
        RECT 6.300 0.965 6.310 1.915 ;
        RECT 6.310 0.965 6.320 1.905 ;
        RECT 6.320 0.965 6.330 1.895 ;
        RECT 6.330 0.965 6.340 1.885 ;
        RECT 6.340 0.965 6.350 1.875 ;
        RECT 6.350 0.965 6.360 1.865 ;
        RECT 6.360 0.965 6.370 1.855 ;
        RECT 6.370 0.965 6.380 1.845 ;
        RECT 6.380 0.965 6.390 1.835 ;
        RECT 6.210 1.765 6.220 2.005 ;
        RECT 6.130 1.845 6.140 2.015 ;
        RECT 6.140 1.835 6.150 2.015 ;
        RECT 6.150 1.825 6.160 2.015 ;
        RECT 6.160 1.815 6.170 2.015 ;
        RECT 6.170 1.805 6.180 2.015 ;
        RECT 6.180 1.795 6.190 2.015 ;
        RECT 6.190 1.785 6.200 2.015 ;
        RECT 6.200 1.775 6.210 2.015 ;
        RECT 0.690 1.030 0.860 2.100 ;
        RECT 0.690 1.930 1.335 2.100 ;
        RECT 1.165 1.930 1.335 2.625 ;
        RECT 1.645 2.455 1.815 2.785 ;
        RECT 1.165 2.455 1.815 2.625 ;
        RECT 1.645 2.615 3.060 2.785 ;
        RECT 3.355 2.975 4.160 3.145 ;
        RECT 4.465 2.745 6.570 2.915 ;
        RECT 6.630 2.745 6.655 2.975 ;
        RECT 6.715 2.805 8.110 2.975 ;
        RECT 6.655 2.755 6.665 2.975 ;
        RECT 6.665 2.765 6.675 2.975 ;
        RECT 6.675 2.775 6.685 2.975 ;
        RECT 6.685 2.785 6.695 2.975 ;
        RECT 6.695 2.795 6.705 2.975 ;
        RECT 6.705 2.805 6.715 2.975 ;
        RECT 6.570 2.745 6.580 2.915 ;
        RECT 6.580 2.745 6.590 2.925 ;
        RECT 6.590 2.745 6.600 2.935 ;
        RECT 6.600 2.745 6.610 2.945 ;
        RECT 6.610 2.745 6.620 2.955 ;
        RECT 6.620 2.745 6.630 2.965 ;
        RECT 4.390 2.745 4.400 2.979 ;
        RECT 4.400 2.745 4.410 2.969 ;
        RECT 4.410 2.745 4.420 2.959 ;
        RECT 4.420 2.745 4.430 2.949 ;
        RECT 4.430 2.745 4.440 2.939 ;
        RECT 4.440 2.745 4.450 2.929 ;
        RECT 4.450 2.745 4.460 2.919 ;
        RECT 4.460 2.745 4.466 2.915 ;
        RECT 4.235 2.900 4.245 3.134 ;
        RECT 4.245 2.890 4.255 3.124 ;
        RECT 4.255 2.880 4.265 3.114 ;
        RECT 4.265 2.870 4.275 3.104 ;
        RECT 4.275 2.860 4.285 3.094 ;
        RECT 4.285 2.850 4.295 3.084 ;
        RECT 4.295 2.840 4.305 3.074 ;
        RECT 4.305 2.830 4.315 3.064 ;
        RECT 4.315 2.820 4.325 3.054 ;
        RECT 4.325 2.810 4.335 3.044 ;
        RECT 4.335 2.800 4.345 3.034 ;
        RECT 4.345 2.790 4.355 3.024 ;
        RECT 4.355 2.780 4.365 3.014 ;
        RECT 4.365 2.770 4.375 3.004 ;
        RECT 4.375 2.760 4.385 2.994 ;
        RECT 4.385 2.750 4.391 2.990 ;
        RECT 4.160 2.975 4.170 3.145 ;
        RECT 4.170 2.965 4.180 3.145 ;
        RECT 4.180 2.955 4.190 3.145 ;
        RECT 4.190 2.945 4.200 3.145 ;
        RECT 4.200 2.935 4.210 3.145 ;
        RECT 4.210 2.925 4.220 3.145 ;
        RECT 4.220 2.915 4.230 3.145 ;
        RECT 4.230 2.905 4.236 3.145 ;
        RECT 3.185 2.675 3.195 3.145 ;
        RECT 3.195 2.685 3.205 3.145 ;
        RECT 3.205 2.695 3.215 3.145 ;
        RECT 3.215 2.705 3.225 3.145 ;
        RECT 3.225 2.715 3.235 3.145 ;
        RECT 3.235 2.725 3.245 3.145 ;
        RECT 3.245 2.735 3.255 3.145 ;
        RECT 3.255 2.745 3.265 3.145 ;
        RECT 3.265 2.755 3.275 3.145 ;
        RECT 3.275 2.765 3.285 3.145 ;
        RECT 3.285 2.775 3.295 3.145 ;
        RECT 3.295 2.785 3.305 3.145 ;
        RECT 3.305 2.795 3.315 3.145 ;
        RECT 3.315 2.805 3.325 3.145 ;
        RECT 3.325 2.815 3.335 3.145 ;
        RECT 3.335 2.825 3.345 3.145 ;
        RECT 3.345 2.835 3.355 3.145 ;
        RECT 3.135 2.625 3.145 2.859 ;
        RECT 3.145 2.635 3.155 2.869 ;
        RECT 3.155 2.645 3.165 2.879 ;
        RECT 3.165 2.655 3.175 2.889 ;
        RECT 3.175 2.665 3.185 2.899 ;
        RECT 3.060 2.615 3.070 2.785 ;
        RECT 3.070 2.615 3.080 2.795 ;
        RECT 3.080 2.615 3.090 2.805 ;
        RECT 3.090 2.615 3.100 2.815 ;
        RECT 3.100 2.615 3.110 2.825 ;
        RECT 3.110 2.615 3.120 2.835 ;
        RECT 3.120 2.615 3.130 2.845 ;
        RECT 3.130 2.615 3.136 2.855 ;
        RECT 7.710 2.395 7.880 2.625 ;
        RECT 6.750 2.395 7.880 2.565 ;
        RECT 7.710 2.455 8.845 2.625 ;
        RECT 8.610 2.455 8.845 3.095 ;
        RECT 7.105 1.125 7.880 1.295 ;
        RECT 7.710 1.125 7.880 1.485 ;
        RECT 8.640 1.185 8.810 1.485 ;
        RECT 7.710 1.315 8.810 1.485 ;
        RECT 8.640 1.185 8.940 1.355 ;
        RECT 1.795 1.945 2.430 2.115 ;
        RECT 2.260 0.995 2.430 2.400 ;
        RECT 2.165 1.945 2.430 2.400 ;
        RECT 2.165 2.230 3.305 2.400 ;
        RECT 3.530 1.795 3.675 1.965 ;
        RECT 3.645 2.625 3.965 2.795 ;
        RECT 3.475 0.525 4.185 0.695 ;
        RECT 4.270 2.395 6.330 2.565 ;
        RECT 7.710 1.675 7.880 2.215 ;
        RECT 6.625 2.045 7.880 2.215 ;
        RECT 7.710 1.675 9.065 1.845 ;
        RECT 9.650 2.115 9.710 2.285 ;
        RECT 9.410 1.885 9.420 2.285 ;
        RECT 9.420 1.895 9.430 2.285 ;
        RECT 9.430 1.905 9.440 2.285 ;
        RECT 9.440 1.915 9.450 2.285 ;
        RECT 9.450 1.925 9.460 2.285 ;
        RECT 9.460 1.935 9.470 2.285 ;
        RECT 9.470 1.945 9.480 2.285 ;
        RECT 9.480 1.955 9.490 2.285 ;
        RECT 9.490 1.965 9.500 2.285 ;
        RECT 9.500 1.975 9.510 2.285 ;
        RECT 9.510 1.985 9.520 2.285 ;
        RECT 9.520 1.995 9.530 2.285 ;
        RECT 9.530 2.005 9.540 2.285 ;
        RECT 9.540 2.015 9.550 2.285 ;
        RECT 9.550 2.025 9.560 2.285 ;
        RECT 9.560 2.035 9.570 2.285 ;
        RECT 9.570 2.045 9.580 2.285 ;
        RECT 9.580 2.055 9.590 2.285 ;
        RECT 9.590 2.065 9.600 2.285 ;
        RECT 9.600 2.075 9.610 2.285 ;
        RECT 9.610 2.085 9.620 2.285 ;
        RECT 9.620 2.095 9.630 2.285 ;
        RECT 9.630 2.105 9.640 2.285 ;
        RECT 9.640 2.115 9.650 2.285 ;
        RECT 9.210 1.685 9.220 1.989 ;
        RECT 9.220 1.695 9.230 1.999 ;
        RECT 9.230 1.705 9.240 2.009 ;
        RECT 9.240 1.715 9.250 2.019 ;
        RECT 9.250 1.725 9.260 2.029 ;
        RECT 9.260 1.735 9.270 2.039 ;
        RECT 9.270 1.745 9.280 2.049 ;
        RECT 9.280 1.755 9.290 2.059 ;
        RECT 9.290 1.765 9.300 2.069 ;
        RECT 9.300 1.775 9.310 2.079 ;
        RECT 9.310 1.785 9.320 2.089 ;
        RECT 9.320 1.795 9.330 2.099 ;
        RECT 9.330 1.805 9.340 2.109 ;
        RECT 9.340 1.815 9.350 2.119 ;
        RECT 9.350 1.825 9.360 2.129 ;
        RECT 9.360 1.835 9.370 2.139 ;
        RECT 9.370 1.845 9.380 2.149 ;
        RECT 9.380 1.855 9.390 2.159 ;
        RECT 9.390 1.865 9.400 2.169 ;
        RECT 9.400 1.875 9.410 2.179 ;
        RECT 9.065 1.675 9.075 1.845 ;
        RECT 9.075 1.675 9.085 1.855 ;
        RECT 9.085 1.675 9.095 1.865 ;
        RECT 9.095 1.675 9.105 1.875 ;
        RECT 9.105 1.675 9.115 1.885 ;
        RECT 9.115 1.675 9.125 1.895 ;
        RECT 9.125 1.675 9.135 1.905 ;
        RECT 9.135 1.675 9.145 1.915 ;
        RECT 9.145 1.675 9.155 1.925 ;
        RECT 9.155 1.675 9.165 1.935 ;
        RECT 9.165 1.675 9.175 1.945 ;
        RECT 9.175 1.675 9.185 1.955 ;
        RECT 9.185 1.675 9.195 1.965 ;
        RECT 9.195 1.675 9.205 1.975 ;
        RECT 9.205 1.675 9.211 1.985 ;
        RECT 6.535 2.045 6.545 2.295 ;
        RECT 6.545 2.045 6.555 2.285 ;
        RECT 6.555 2.045 6.565 2.275 ;
        RECT 6.565 2.045 6.575 2.265 ;
        RECT 6.575 2.045 6.585 2.255 ;
        RECT 6.585 2.045 6.595 2.245 ;
        RECT 6.595 2.045 6.605 2.235 ;
        RECT 6.605 2.045 6.615 2.225 ;
        RECT 6.615 2.045 6.625 2.215 ;
        RECT 6.500 2.080 6.510 2.330 ;
        RECT 6.510 2.070 6.520 2.320 ;
        RECT 6.520 2.060 6.530 2.310 ;
        RECT 6.530 2.050 6.536 2.304 ;
        RECT 6.330 2.250 6.340 2.564 ;
        RECT 6.340 2.240 6.350 2.564 ;
        RECT 6.350 2.230 6.360 2.564 ;
        RECT 6.360 2.220 6.370 2.564 ;
        RECT 6.370 2.210 6.380 2.564 ;
        RECT 6.380 2.200 6.390 2.564 ;
        RECT 6.390 2.190 6.400 2.564 ;
        RECT 6.400 2.180 6.410 2.564 ;
        RECT 6.410 2.170 6.420 2.564 ;
        RECT 6.420 2.160 6.430 2.564 ;
        RECT 6.430 2.150 6.440 2.564 ;
        RECT 6.440 2.140 6.450 2.564 ;
        RECT 6.450 2.130 6.460 2.564 ;
        RECT 6.460 2.120 6.470 2.564 ;
        RECT 6.470 2.110 6.480 2.564 ;
        RECT 6.480 2.100 6.490 2.564 ;
        RECT 6.490 2.090 6.500 2.564 ;
        RECT 4.195 2.395 4.205 2.629 ;
        RECT 4.205 2.395 4.215 2.619 ;
        RECT 4.215 2.395 4.225 2.609 ;
        RECT 4.225 2.395 4.235 2.599 ;
        RECT 4.235 2.395 4.245 2.589 ;
        RECT 4.245 2.395 4.255 2.579 ;
        RECT 4.255 2.395 4.265 2.569 ;
        RECT 4.265 2.395 4.271 2.565 ;
        RECT 4.040 2.550 4.050 2.784 ;
        RECT 4.050 2.540 4.060 2.774 ;
        RECT 4.060 2.530 4.070 2.764 ;
        RECT 4.070 2.520 4.080 2.754 ;
        RECT 4.080 2.510 4.090 2.744 ;
        RECT 4.090 2.500 4.100 2.734 ;
        RECT 4.100 2.490 4.110 2.724 ;
        RECT 4.110 2.480 4.120 2.714 ;
        RECT 4.120 2.470 4.130 2.704 ;
        RECT 4.130 2.460 4.140 2.694 ;
        RECT 4.140 2.450 4.150 2.684 ;
        RECT 4.150 2.440 4.160 2.674 ;
        RECT 4.160 2.430 4.170 2.664 ;
        RECT 4.170 2.420 4.180 2.654 ;
        RECT 4.180 2.410 4.190 2.644 ;
        RECT 4.190 2.400 4.196 2.640 ;
        RECT 3.965 2.625 3.975 2.795 ;
        RECT 3.975 2.615 3.985 2.795 ;
        RECT 3.985 2.605 3.995 2.795 ;
        RECT 3.995 2.595 4.005 2.795 ;
        RECT 4.005 2.585 4.015 2.795 ;
        RECT 4.015 2.575 4.025 2.795 ;
        RECT 4.025 2.565 4.035 2.795 ;
        RECT 4.035 2.555 4.041 2.795 ;
        RECT 3.570 2.560 3.580 2.794 ;
        RECT 3.580 2.570 3.590 2.794 ;
        RECT 3.590 2.580 3.600 2.794 ;
        RECT 3.600 2.590 3.610 2.794 ;
        RECT 3.610 2.600 3.620 2.794 ;
        RECT 3.620 2.610 3.630 2.794 ;
        RECT 3.630 2.620 3.640 2.794 ;
        RECT 3.640 2.625 3.646 2.795 ;
        RECT 3.530 2.520 3.540 2.754 ;
        RECT 3.540 2.530 3.550 2.764 ;
        RECT 3.550 2.540 3.560 2.774 ;
        RECT 3.560 2.550 3.570 2.784 ;
        RECT 3.475 1.405 3.485 2.699 ;
        RECT 3.485 1.415 3.495 2.709 ;
        RECT 3.495 1.425 3.505 2.719 ;
        RECT 3.505 1.435 3.515 2.729 ;
        RECT 3.515 1.445 3.525 2.739 ;
        RECT 3.525 1.450 3.531 2.750 ;
        RECT 3.360 0.525 3.370 2.585 ;
        RECT 3.370 0.525 3.380 2.595 ;
        RECT 3.380 0.525 3.390 2.605 ;
        RECT 3.390 0.525 3.400 2.615 ;
        RECT 3.400 0.525 3.410 2.625 ;
        RECT 3.410 0.525 3.420 2.635 ;
        RECT 3.420 0.525 3.430 2.645 ;
        RECT 3.430 0.525 3.440 2.655 ;
        RECT 3.440 0.525 3.450 2.665 ;
        RECT 3.450 0.525 3.460 2.675 ;
        RECT 3.460 0.525 3.470 2.685 ;
        RECT 3.470 0.525 3.476 2.695 ;
        RECT 3.305 0.525 3.315 1.469 ;
        RECT 3.315 0.525 3.325 1.479 ;
        RECT 3.325 0.525 3.335 1.489 ;
        RECT 3.335 0.525 3.345 1.499 ;
        RECT 3.345 0.525 3.355 1.509 ;
        RECT 3.355 0.525 3.361 1.519 ;
        RECT 3.305 2.230 3.315 2.530 ;
        RECT 3.315 2.230 3.325 2.540 ;
        RECT 3.325 2.230 3.335 2.550 ;
        RECT 3.335 2.230 3.345 2.560 ;
        RECT 3.345 2.230 3.355 2.570 ;
        RECT 3.355 2.230 3.361 2.580 ;
        RECT 10.885 1.400 11.055 2.215 ;
        RECT 10.600 2.045 11.055 2.215 ;
        RECT 10.940 1.025 11.110 1.570 ;
        RECT 10.000 1.400 11.110 1.570 ;
        RECT 10.940 1.025 11.330 1.195 ;
        RECT 8.120 0.965 8.360 1.135 ;
        RECT 8.090 2.025 8.390 2.275 ;
        RECT 8.090 2.025 8.845 2.195 ;
        RECT 8.565 0.835 9.015 1.005 ;
        RECT 9.190 0.895 9.380 1.415 ;
        RECT 9.230 2.465 9.430 3.015 ;
        RECT 9.455 0.895 9.490 1.490 ;
        RECT 9.580 1.320 9.640 1.490 ;
        RECT 9.230 2.465 9.890 2.645 ;
        RECT 10.060 2.465 10.655 2.645 ;
        RECT 10.725 2.395 10.780 2.645 ;
        RECT 11.235 1.860 11.405 2.565 ;
        RECT 10.860 2.395 11.405 2.565 ;
        RECT 11.355 1.675 11.525 2.030 ;
        RECT 11.235 1.860 11.525 2.030 ;
        RECT 11.355 1.675 12.460 1.845 ;
        RECT 10.780 2.395 10.790 2.635 ;
        RECT 10.790 2.395 10.800 2.625 ;
        RECT 10.800 2.395 10.810 2.615 ;
        RECT 10.810 2.395 10.820 2.605 ;
        RECT 10.820 2.395 10.830 2.595 ;
        RECT 10.830 2.395 10.840 2.585 ;
        RECT 10.840 2.395 10.850 2.575 ;
        RECT 10.850 2.395 10.860 2.565 ;
        RECT 10.655 2.465 10.665 2.645 ;
        RECT 10.665 2.455 10.675 2.645 ;
        RECT 10.675 2.445 10.685 2.645 ;
        RECT 10.685 2.435 10.695 2.645 ;
        RECT 10.695 2.425 10.705 2.645 ;
        RECT 10.705 2.415 10.715 2.645 ;
        RECT 10.715 2.405 10.725 2.645 ;
        RECT 9.890 1.805 9.900 2.645 ;
        RECT 9.900 1.815 9.910 2.645 ;
        RECT 9.910 1.825 9.920 2.645 ;
        RECT 9.920 1.835 9.930 2.645 ;
        RECT 9.930 1.845 9.940 2.645 ;
        RECT 9.940 1.855 9.950 2.645 ;
        RECT 9.950 1.865 9.960 2.645 ;
        RECT 9.960 1.875 9.970 2.645 ;
        RECT 9.970 1.885 9.980 2.645 ;
        RECT 9.980 1.895 9.990 2.645 ;
        RECT 9.990 1.905 10.000 2.645 ;
        RECT 10.000 1.915 10.010 2.645 ;
        RECT 10.010 1.925 10.020 2.645 ;
        RECT 10.020 1.935 10.030 2.645 ;
        RECT 10.030 1.945 10.040 2.645 ;
        RECT 10.040 1.955 10.050 2.645 ;
        RECT 10.050 1.965 10.060 2.645 ;
        RECT 9.810 1.725 9.820 1.959 ;
        RECT 9.820 1.735 9.830 1.969 ;
        RECT 9.830 1.745 9.840 1.979 ;
        RECT 9.840 1.755 9.850 1.989 ;
        RECT 9.850 1.765 9.860 1.999 ;
        RECT 9.860 1.775 9.870 2.009 ;
        RECT 9.870 1.785 9.880 2.019 ;
        RECT 9.880 1.795 9.890 2.029 ;
        RECT 9.640 1.320 9.650 1.790 ;
        RECT 9.650 1.320 9.660 1.800 ;
        RECT 9.660 1.320 9.670 1.810 ;
        RECT 9.670 1.320 9.680 1.820 ;
        RECT 9.680 1.320 9.690 1.830 ;
        RECT 9.690 1.320 9.700 1.840 ;
        RECT 9.700 1.320 9.710 1.850 ;
        RECT 9.710 1.320 9.720 1.860 ;
        RECT 9.720 1.320 9.730 1.870 ;
        RECT 9.730 1.320 9.740 1.880 ;
        RECT 9.740 1.320 9.750 1.890 ;
        RECT 9.750 1.320 9.760 1.900 ;
        RECT 9.760 1.320 9.770 1.910 ;
        RECT 9.770 1.320 9.780 1.920 ;
        RECT 9.780 1.320 9.790 1.930 ;
        RECT 9.790 1.320 9.800 1.940 ;
        RECT 9.800 1.320 9.810 1.950 ;
        RECT 9.490 1.240 9.500 1.490 ;
        RECT 9.500 1.250 9.510 1.490 ;
        RECT 9.510 1.260 9.520 1.490 ;
        RECT 9.520 1.270 9.530 1.490 ;
        RECT 9.530 1.280 9.540 1.490 ;
        RECT 9.540 1.290 9.550 1.490 ;
        RECT 9.550 1.300 9.560 1.490 ;
        RECT 9.560 1.310 9.570 1.490 ;
        RECT 9.570 1.320 9.580 1.490 ;
        RECT 9.380 0.895 9.390 1.415 ;
        RECT 9.390 0.895 9.400 1.425 ;
        RECT 9.400 0.895 9.410 1.435 ;
        RECT 9.410 0.895 9.420 1.445 ;
        RECT 9.420 0.895 9.430 1.455 ;
        RECT 9.430 0.895 9.440 1.465 ;
        RECT 9.440 0.895 9.450 1.475 ;
        RECT 9.450 0.895 9.456 1.485 ;
        RECT 9.060 2.170 9.070 3.014 ;
        RECT 9.070 2.180 9.080 3.014 ;
        RECT 9.080 2.190 9.090 3.014 ;
        RECT 9.090 2.200 9.100 3.014 ;
        RECT 9.100 2.210 9.110 3.014 ;
        RECT 9.110 2.220 9.120 3.014 ;
        RECT 9.120 2.230 9.130 3.014 ;
        RECT 9.130 2.240 9.140 3.014 ;
        RECT 9.140 2.250 9.150 3.014 ;
        RECT 9.150 2.260 9.160 3.014 ;
        RECT 9.160 2.270 9.170 3.014 ;
        RECT 9.170 2.280 9.180 3.014 ;
        RECT 9.180 2.290 9.190 3.014 ;
        RECT 9.190 2.300 9.200 3.014 ;
        RECT 9.200 2.310 9.210 3.014 ;
        RECT 9.210 2.320 9.220 3.014 ;
        RECT 9.220 2.330 9.230 3.014 ;
        RECT 9.150 0.895 9.160 1.139 ;
        RECT 9.160 0.895 9.170 1.149 ;
        RECT 9.170 0.895 9.180 1.159 ;
        RECT 9.180 0.895 9.190 1.169 ;
        RECT 9.090 0.845 9.100 1.079 ;
        RECT 9.100 0.855 9.110 1.089 ;
        RECT 9.110 0.865 9.120 1.099 ;
        RECT 9.120 0.875 9.130 1.109 ;
        RECT 9.130 0.885 9.140 1.119 ;
        RECT 9.140 0.895 9.150 1.129 ;
        RECT 9.015 0.835 9.025 1.005 ;
        RECT 9.025 0.835 9.035 1.015 ;
        RECT 9.035 0.835 9.045 1.025 ;
        RECT 9.045 0.835 9.055 1.035 ;
        RECT 9.055 0.835 9.065 1.045 ;
        RECT 9.065 0.835 9.075 1.055 ;
        RECT 9.075 0.835 9.085 1.065 ;
        RECT 9.085 0.835 9.091 1.075 ;
        RECT 8.925 2.035 8.935 2.275 ;
        RECT 8.935 2.045 8.945 2.285 ;
        RECT 8.945 2.055 8.955 2.295 ;
        RECT 8.955 2.065 8.965 2.305 ;
        RECT 8.965 2.075 8.975 2.315 ;
        RECT 8.975 2.085 8.985 2.325 ;
        RECT 8.985 2.095 8.995 2.335 ;
        RECT 8.995 2.105 9.005 2.345 ;
        RECT 9.005 2.115 9.015 2.355 ;
        RECT 9.015 2.125 9.025 2.365 ;
        RECT 9.025 2.135 9.035 2.375 ;
        RECT 9.035 2.145 9.045 2.385 ;
        RECT 9.045 2.155 9.055 2.395 ;
        RECT 9.055 2.160 9.061 2.404 ;
        RECT 8.845 2.025 8.855 2.195 ;
        RECT 8.855 2.025 8.865 2.205 ;
        RECT 8.865 2.025 8.875 2.215 ;
        RECT 8.875 2.025 8.885 2.225 ;
        RECT 8.885 2.025 8.895 2.235 ;
        RECT 8.895 2.025 8.905 2.245 ;
        RECT 8.905 2.025 8.915 2.255 ;
        RECT 8.915 2.025 8.925 2.265 ;
        RECT 8.490 0.835 8.500 1.069 ;
        RECT 8.500 0.835 8.510 1.059 ;
        RECT 8.510 0.835 8.520 1.049 ;
        RECT 8.520 0.835 8.530 1.039 ;
        RECT 8.530 0.835 8.540 1.029 ;
        RECT 8.540 0.835 8.550 1.019 ;
        RECT 8.550 0.835 8.560 1.009 ;
        RECT 8.560 0.835 8.566 1.005 ;
        RECT 8.435 0.890 8.445 1.124 ;
        RECT 8.445 0.880 8.455 1.114 ;
        RECT 8.455 0.870 8.465 1.104 ;
        RECT 8.465 0.860 8.475 1.094 ;
        RECT 8.475 0.850 8.485 1.084 ;
        RECT 8.485 0.840 8.491 1.080 ;
        RECT 8.360 0.965 8.370 1.135 ;
        RECT 8.370 0.955 8.380 1.135 ;
        RECT 8.380 0.945 8.390 1.135 ;
        RECT 8.390 0.935 8.400 1.135 ;
        RECT 8.400 0.925 8.410 1.135 ;
        RECT 8.410 0.915 8.420 1.135 ;
        RECT 8.420 0.905 8.430 1.135 ;
        RECT 8.430 0.895 8.436 1.135 ;
  END 
END FFDSHQHD3XHT

MACRO FFDSHQHD2XHT
  CLASS  CORE ;
  FOREIGN FFDSHQHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.890 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.325 0.720 10.660 1.495 ;
        RECT 10.325 2.230 10.660 3.210 ;
        RECT 10.325 1.320 11.665 1.495 ;
        RECT 10.325 2.230 11.665 2.430 ;
        RECT 11.365 0.720 11.665 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.500 2.560 2.205 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.995 ;
        RECT 2.175 -0.300 2.475 1.230 ;
        RECT 4.035 -0.300 4.335 1.115 ;
        RECT 5.345 -0.300 5.645 0.435 ;
        RECT 6.445 -0.300 6.745 0.435 ;
        RECT 8.895 -0.300 9.195 0.870 ;
        RECT 10.900 -0.300 11.145 1.120 ;
        RECT 0.000 -0.300 11.890 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.870 1.260 1.130 1.800 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.610 1.345 4.840 1.430 ;
        RECT 4.670 0.615 4.825 1.665 ;
        RECT 4.610 0.615 4.825 1.430 ;
        RECT 4.670 1.345 4.840 1.665 ;
        RECT 4.670 1.495 5.175 1.665 ;
        RECT 6.915 0.500 7.085 0.785 ;
        RECT 4.610 0.615 7.085 0.785 ;
        RECT 6.915 0.500 8.715 0.670 ;
        RECT 4.610 0.615 8.715 0.670 ;
        RECT 8.545 0.500 8.715 1.220 ;
        RECT 9.375 0.655 9.545 1.220 ;
        RECT 8.545 1.050 9.545 1.220 ;
        RECT 9.375 0.655 9.895 0.825 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 1.980 0.340 3.990 ;
        RECT 2.145 3.215 2.445 3.990 ;
        RECT 4.175 3.095 4.475 3.990 ;
        RECT 5.275 3.095 5.575 3.990 ;
        RECT 6.375 3.175 6.675 3.990 ;
        RECT 8.895 2.845 9.195 3.990 ;
        RECT 9.815 2.745 10.115 3.990 ;
        RECT 10.845 2.635 11.145 3.990 ;
        RECT 0.000 3.390 11.890 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.000 1.980 1.170 2.215 ;
        RECT 0.870 2.045 1.170 2.215 ;
        RECT 1.145 0.825 1.480 0.995 ;
        RECT 1.000 1.980 1.480 2.150 ;
        RECT 1.310 0.825 1.480 2.150 ;
        RECT 1.310 1.610 1.540 1.910 ;
        RECT 3.115 2.165 3.285 2.335 ;
        RECT 3.130 0.995 3.300 1.495 ;
        RECT 3.130 1.325 3.415 1.495 ;
        RECT 3.315 1.325 3.415 2.335 ;
        RECT 3.485 1.325 4.150 1.495 ;
        RECT 4.320 1.405 4.330 1.865 ;
        RECT 4.330 1.415 4.340 1.865 ;
        RECT 4.340 1.425 4.350 1.865 ;
        RECT 4.350 1.435 4.360 1.865 ;
        RECT 4.360 1.445 4.370 1.865 ;
        RECT 4.370 1.455 4.380 1.865 ;
        RECT 4.380 1.465 4.390 1.865 ;
        RECT 4.390 1.475 4.400 1.865 ;
        RECT 4.400 1.485 4.410 1.865 ;
        RECT 4.410 1.495 4.420 1.865 ;
        RECT 4.420 1.505 4.430 1.865 ;
        RECT 4.430 1.515 4.440 1.865 ;
        RECT 4.440 1.525 4.450 1.865 ;
        RECT 4.450 1.535 4.460 1.865 ;
        RECT 4.460 1.545 4.470 1.865 ;
        RECT 4.470 1.555 4.480 1.865 ;
        RECT 4.480 1.565 4.490 1.865 ;
        RECT 4.250 1.335 4.260 1.595 ;
        RECT 4.260 1.345 4.270 1.605 ;
        RECT 4.270 1.355 4.280 1.615 ;
        RECT 4.280 1.365 4.290 1.625 ;
        RECT 4.290 1.375 4.300 1.635 ;
        RECT 4.300 1.385 4.310 1.645 ;
        RECT 4.310 1.395 4.320 1.655 ;
        RECT 4.150 1.325 4.160 1.495 ;
        RECT 4.160 1.325 4.170 1.505 ;
        RECT 4.170 1.325 4.180 1.515 ;
        RECT 4.180 1.325 4.190 1.525 ;
        RECT 4.190 1.325 4.200 1.535 ;
        RECT 4.200 1.325 4.210 1.545 ;
        RECT 4.210 1.325 4.220 1.555 ;
        RECT 4.220 1.325 4.230 1.565 ;
        RECT 4.230 1.325 4.240 1.575 ;
        RECT 4.240 1.325 4.250 1.585 ;
        RECT 3.415 1.325 3.425 2.325 ;
        RECT 3.425 1.325 3.435 2.315 ;
        RECT 3.435 1.325 3.445 2.305 ;
        RECT 3.445 1.325 3.455 2.295 ;
        RECT 3.455 1.325 3.465 2.285 ;
        RECT 3.465 1.325 3.475 2.275 ;
        RECT 3.475 1.325 3.485 2.265 ;
        RECT 3.285 2.165 3.295 2.335 ;
        RECT 3.295 2.155 3.305 2.335 ;
        RECT 3.305 2.145 3.315 2.335 ;
        RECT 3.775 1.675 4.075 2.215 ;
        RECT 5.005 0.965 5.175 1.265 ;
        RECT 5.035 1.845 5.205 2.215 ;
        RECT 3.770 2.045 5.205 2.215 ;
        RECT 5.035 1.845 5.305 2.015 ;
        RECT 5.005 1.095 5.445 1.265 ;
        RECT 5.615 1.495 6.285 1.665 ;
        RECT 5.445 1.095 5.455 1.965 ;
        RECT 5.455 1.095 5.465 1.955 ;
        RECT 5.465 1.095 5.475 1.945 ;
        RECT 5.475 1.095 5.485 1.935 ;
        RECT 5.485 1.095 5.495 1.925 ;
        RECT 5.495 1.095 5.505 1.915 ;
        RECT 5.505 1.095 5.515 1.905 ;
        RECT 5.515 1.095 5.525 1.895 ;
        RECT 5.525 1.095 5.535 1.885 ;
        RECT 5.535 1.095 5.545 1.875 ;
        RECT 5.545 1.095 5.555 1.865 ;
        RECT 5.555 1.095 5.565 1.855 ;
        RECT 5.565 1.095 5.575 1.845 ;
        RECT 5.575 1.095 5.585 1.835 ;
        RECT 5.585 1.095 5.595 1.825 ;
        RECT 5.595 1.095 5.605 1.815 ;
        RECT 5.605 1.095 5.615 1.805 ;
        RECT 5.405 1.745 5.415 2.005 ;
        RECT 5.415 1.735 5.425 1.995 ;
        RECT 5.425 1.725 5.435 1.985 ;
        RECT 5.435 1.715 5.445 1.975 ;
        RECT 5.305 1.845 5.315 2.015 ;
        RECT 5.315 1.835 5.325 2.015 ;
        RECT 5.325 1.825 5.335 2.015 ;
        RECT 5.335 1.815 5.345 2.015 ;
        RECT 5.345 1.805 5.355 2.015 ;
        RECT 5.355 1.795 5.365 2.015 ;
        RECT 5.365 1.785 5.375 2.015 ;
        RECT 5.375 1.775 5.385 2.015 ;
        RECT 5.385 1.765 5.395 2.015 ;
        RECT 5.395 1.755 5.405 2.015 ;
        RECT 6.505 2.395 6.675 2.645 ;
        RECT 5.825 2.395 6.675 2.565 ;
        RECT 6.505 2.475 7.640 2.645 ;
        RECT 7.470 2.475 7.640 2.775 ;
        RECT 5.895 0.965 6.655 1.135 ;
        RECT 6.485 0.965 6.655 1.510 ;
        RECT 7.425 1.205 7.725 1.510 ;
        RECT 6.485 1.340 7.725 1.510 ;
        RECT 0.170 0.720 0.340 1.790 ;
        RECT 0.170 1.620 0.690 1.790 ;
        RECT 0.520 1.620 0.690 2.665 ;
        RECT 0.520 2.495 1.230 2.665 ;
        RECT 1.060 2.495 1.230 3.035 ;
        RECT 1.060 2.865 3.640 3.035 ;
        RECT 6.155 2.745 6.325 2.995 ;
        RECT 3.835 2.745 6.325 2.915 ;
        RECT 6.155 2.825 7.225 2.995 ;
        RECT 7.055 2.825 7.225 3.190 ;
        RECT 7.055 3.020 7.865 3.190 ;
        RECT 3.760 2.745 3.770 2.979 ;
        RECT 3.770 2.745 3.780 2.969 ;
        RECT 3.780 2.745 3.790 2.959 ;
        RECT 3.790 2.745 3.800 2.949 ;
        RECT 3.800 2.745 3.810 2.939 ;
        RECT 3.810 2.745 3.820 2.929 ;
        RECT 3.820 2.745 3.830 2.919 ;
        RECT 3.830 2.745 3.836 2.915 ;
        RECT 3.715 2.790 3.725 3.024 ;
        RECT 3.725 2.780 3.735 3.014 ;
        RECT 3.735 2.770 3.745 3.004 ;
        RECT 3.745 2.760 3.755 2.994 ;
        RECT 3.755 2.750 3.761 2.990 ;
        RECT 3.640 2.865 3.650 3.035 ;
        RECT 3.650 2.855 3.660 3.035 ;
        RECT 3.660 2.845 3.670 3.035 ;
        RECT 3.670 2.835 3.680 3.035 ;
        RECT 3.680 2.825 3.690 3.035 ;
        RECT 3.690 2.815 3.700 3.035 ;
        RECT 3.700 2.805 3.710 3.035 ;
        RECT 3.710 2.795 3.716 3.035 ;
        RECT 1.720 0.990 1.890 2.685 ;
        RECT 1.440 2.345 1.890 2.685 ;
        RECT 2.765 0.525 2.935 2.685 ;
        RECT 2.765 1.795 3.135 1.965 ;
        RECT 1.440 2.515 3.490 2.685 ;
        RECT 2.765 0.525 3.595 0.695 ;
        RECT 3.685 2.395 5.475 2.565 ;
        RECT 6.505 1.690 6.675 2.210 ;
        RECT 5.755 2.040 6.675 2.210 ;
        RECT 6.505 1.690 7.880 1.860 ;
        RECT 8.385 2.115 8.505 2.285 ;
        RECT 8.205 1.945 8.215 2.285 ;
        RECT 8.215 1.955 8.225 2.285 ;
        RECT 8.225 1.965 8.235 2.285 ;
        RECT 8.235 1.975 8.245 2.285 ;
        RECT 8.245 1.985 8.255 2.285 ;
        RECT 8.255 1.995 8.265 2.285 ;
        RECT 8.265 2.005 8.275 2.285 ;
        RECT 8.275 2.015 8.285 2.285 ;
        RECT 8.285 2.025 8.295 2.285 ;
        RECT 8.295 2.035 8.305 2.285 ;
        RECT 8.305 2.045 8.315 2.285 ;
        RECT 8.315 2.055 8.325 2.285 ;
        RECT 8.325 2.065 8.335 2.285 ;
        RECT 8.335 2.075 8.345 2.285 ;
        RECT 8.345 2.085 8.355 2.285 ;
        RECT 8.355 2.095 8.365 2.285 ;
        RECT 8.365 2.105 8.375 2.285 ;
        RECT 8.375 2.115 8.385 2.285 ;
        RECT 8.100 1.840 8.110 2.080 ;
        RECT 8.110 1.850 8.120 2.090 ;
        RECT 8.120 1.860 8.130 2.100 ;
        RECT 8.130 1.870 8.140 2.110 ;
        RECT 8.140 1.880 8.150 2.120 ;
        RECT 8.150 1.890 8.160 2.130 ;
        RECT 8.160 1.900 8.170 2.140 ;
        RECT 8.170 1.910 8.180 2.150 ;
        RECT 8.180 1.920 8.190 2.160 ;
        RECT 8.190 1.930 8.200 2.170 ;
        RECT 8.200 1.935 8.206 2.179 ;
        RECT 7.880 1.690 7.890 1.860 ;
        RECT 7.890 1.690 7.900 1.870 ;
        RECT 7.900 1.690 7.910 1.880 ;
        RECT 7.910 1.690 7.920 1.890 ;
        RECT 7.920 1.690 7.930 1.900 ;
        RECT 7.930 1.690 7.940 1.910 ;
        RECT 7.940 1.690 7.950 1.920 ;
        RECT 7.950 1.690 7.960 1.930 ;
        RECT 7.960 1.690 7.970 1.940 ;
        RECT 7.970 1.690 7.980 1.950 ;
        RECT 7.980 1.690 7.990 1.960 ;
        RECT 7.990 1.690 8.000 1.970 ;
        RECT 8.000 1.690 8.010 1.980 ;
        RECT 8.010 1.690 8.020 1.990 ;
        RECT 8.020 1.690 8.030 2.000 ;
        RECT 8.030 1.690 8.040 2.010 ;
        RECT 8.040 1.690 8.050 2.020 ;
        RECT 8.050 1.690 8.060 2.030 ;
        RECT 8.060 1.690 8.070 2.040 ;
        RECT 8.070 1.690 8.080 2.050 ;
        RECT 8.080 1.690 8.090 2.060 ;
        RECT 8.090 1.690 8.100 2.070 ;
        RECT 5.680 2.040 5.690 2.274 ;
        RECT 5.690 2.040 5.700 2.264 ;
        RECT 5.700 2.040 5.710 2.254 ;
        RECT 5.710 2.040 5.720 2.244 ;
        RECT 5.720 2.040 5.730 2.234 ;
        RECT 5.730 2.040 5.740 2.224 ;
        RECT 5.740 2.040 5.750 2.214 ;
        RECT 5.750 2.040 5.756 2.210 ;
        RECT 5.645 2.075 5.655 2.309 ;
        RECT 5.655 2.065 5.665 2.299 ;
        RECT 5.665 2.055 5.675 2.289 ;
        RECT 5.675 2.045 5.681 2.285 ;
        RECT 5.475 2.245 5.485 2.565 ;
        RECT 5.485 2.235 5.495 2.565 ;
        RECT 5.495 2.225 5.505 2.565 ;
        RECT 5.505 2.215 5.515 2.565 ;
        RECT 5.515 2.205 5.525 2.565 ;
        RECT 5.525 2.195 5.535 2.565 ;
        RECT 5.535 2.185 5.545 2.565 ;
        RECT 5.545 2.175 5.555 2.565 ;
        RECT 5.555 2.165 5.565 2.565 ;
        RECT 5.565 2.155 5.575 2.565 ;
        RECT 5.575 2.145 5.585 2.565 ;
        RECT 5.585 2.135 5.595 2.565 ;
        RECT 5.595 2.125 5.605 2.565 ;
        RECT 5.605 2.115 5.615 2.565 ;
        RECT 5.615 2.105 5.625 2.565 ;
        RECT 5.625 2.095 5.635 2.565 ;
        RECT 5.635 2.085 5.645 2.565 ;
        RECT 3.610 2.395 3.620 2.629 ;
        RECT 3.620 2.395 3.630 2.619 ;
        RECT 3.630 2.395 3.640 2.609 ;
        RECT 3.640 2.395 3.650 2.599 ;
        RECT 3.650 2.395 3.660 2.589 ;
        RECT 3.660 2.395 3.670 2.579 ;
        RECT 3.670 2.395 3.680 2.569 ;
        RECT 3.680 2.395 3.686 2.565 ;
        RECT 3.565 2.440 3.575 2.674 ;
        RECT 3.575 2.430 3.585 2.664 ;
        RECT 3.585 2.420 3.595 2.654 ;
        RECT 3.595 2.410 3.605 2.644 ;
        RECT 3.605 2.400 3.611 2.640 ;
        RECT 3.490 2.515 3.500 2.685 ;
        RECT 3.500 2.505 3.510 2.685 ;
        RECT 3.510 2.495 3.520 2.685 ;
        RECT 3.520 2.485 3.530 2.685 ;
        RECT 3.530 2.475 3.540 2.685 ;
        RECT 3.540 2.465 3.550 2.685 ;
        RECT 3.550 2.455 3.560 2.685 ;
        RECT 3.560 2.445 3.566 2.685 ;
        RECT 9.515 1.400 9.685 2.215 ;
        RECT 9.385 2.045 9.685 2.215 ;
        RECT 9.725 1.025 9.895 1.570 ;
        RECT 8.785 1.400 9.895 1.570 ;
        RECT 9.725 1.025 10.115 1.195 ;
        RECT 6.855 0.990 7.135 1.160 ;
        RECT 6.885 2.125 7.740 2.295 ;
        RECT 7.350 0.850 7.800 1.020 ;
        RECT 7.845 0.850 7.875 1.065 ;
        RECT 7.920 0.895 8.175 1.065 ;
        RECT 8.040 0.895 8.175 1.415 ;
        RECT 8.025 2.465 8.315 2.675 ;
        RECT 8.025 2.465 8.685 2.645 ;
        RECT 8.855 2.465 9.440 2.645 ;
        RECT 9.510 2.395 9.565 2.645 ;
        RECT 9.885 1.860 10.055 2.565 ;
        RECT 9.645 2.395 10.055 2.565 ;
        RECT 10.140 1.675 10.310 2.030 ;
        RECT 9.885 1.860 10.310 2.030 ;
        RECT 10.140 1.675 11.185 1.845 ;
        RECT 9.565 2.395 9.575 2.635 ;
        RECT 9.575 2.395 9.585 2.625 ;
        RECT 9.585 2.395 9.595 2.615 ;
        RECT 9.595 2.395 9.605 2.605 ;
        RECT 9.605 2.395 9.615 2.595 ;
        RECT 9.615 2.395 9.625 2.585 ;
        RECT 9.625 2.395 9.635 2.575 ;
        RECT 9.635 2.395 9.645 2.565 ;
        RECT 9.440 2.465 9.450 2.645 ;
        RECT 9.450 2.455 9.460 2.645 ;
        RECT 9.460 2.445 9.470 2.645 ;
        RECT 9.470 2.435 9.480 2.645 ;
        RECT 9.480 2.425 9.490 2.645 ;
        RECT 9.490 2.415 9.500 2.645 ;
        RECT 9.500 2.405 9.510 2.645 ;
        RECT 8.685 1.800 8.695 2.644 ;
        RECT 8.695 1.810 8.705 2.644 ;
        RECT 8.705 1.820 8.715 2.644 ;
        RECT 8.715 1.830 8.725 2.644 ;
        RECT 8.725 1.840 8.735 2.644 ;
        RECT 8.735 1.850 8.745 2.644 ;
        RECT 8.745 1.860 8.755 2.644 ;
        RECT 8.755 1.870 8.765 2.644 ;
        RECT 8.765 1.880 8.775 2.644 ;
        RECT 8.775 1.890 8.785 2.644 ;
        RECT 8.785 1.900 8.795 2.644 ;
        RECT 8.795 1.910 8.805 2.644 ;
        RECT 8.805 1.920 8.815 2.644 ;
        RECT 8.815 1.930 8.825 2.644 ;
        RECT 8.825 1.940 8.835 2.644 ;
        RECT 8.835 1.950 8.845 2.644 ;
        RECT 8.845 1.960 8.855 2.644 ;
        RECT 8.605 1.720 8.615 1.960 ;
        RECT 8.615 1.730 8.625 1.970 ;
        RECT 8.625 1.740 8.635 1.980 ;
        RECT 8.635 1.750 8.645 1.990 ;
        RECT 8.645 1.760 8.655 2.000 ;
        RECT 8.655 1.770 8.665 2.010 ;
        RECT 8.665 1.780 8.675 2.020 ;
        RECT 8.675 1.790 8.685 2.030 ;
        RECT 8.455 1.400 8.465 1.810 ;
        RECT 8.465 1.400 8.475 1.820 ;
        RECT 8.475 1.400 8.485 1.830 ;
        RECT 8.485 1.400 8.495 1.840 ;
        RECT 8.495 1.400 8.505 1.850 ;
        RECT 8.505 1.400 8.515 1.860 ;
        RECT 8.515 1.400 8.525 1.870 ;
        RECT 8.525 1.400 8.535 1.880 ;
        RECT 8.535 1.400 8.545 1.890 ;
        RECT 8.545 1.400 8.555 1.900 ;
        RECT 8.555 1.400 8.565 1.910 ;
        RECT 8.565 1.400 8.575 1.920 ;
        RECT 8.575 1.400 8.585 1.930 ;
        RECT 8.585 1.400 8.595 1.940 ;
        RECT 8.595 1.400 8.605 1.950 ;
        RECT 8.435 1.390 8.445 1.790 ;
        RECT 8.445 1.400 8.455 1.800 ;
        RECT 8.330 1.285 8.340 1.569 ;
        RECT 8.340 1.295 8.350 1.569 ;
        RECT 8.350 1.305 8.360 1.569 ;
        RECT 8.360 1.315 8.370 1.569 ;
        RECT 8.370 1.325 8.380 1.569 ;
        RECT 8.380 1.335 8.390 1.569 ;
        RECT 8.390 1.345 8.400 1.569 ;
        RECT 8.400 1.355 8.410 1.569 ;
        RECT 8.410 1.365 8.420 1.569 ;
        RECT 8.420 1.375 8.430 1.569 ;
        RECT 8.430 1.380 8.436 1.570 ;
        RECT 8.275 1.230 8.285 1.514 ;
        RECT 8.285 1.240 8.295 1.524 ;
        RECT 8.295 1.250 8.305 1.534 ;
        RECT 8.305 1.260 8.315 1.544 ;
        RECT 8.315 1.270 8.325 1.554 ;
        RECT 8.325 1.275 8.331 1.565 ;
        RECT 8.175 0.895 8.185 1.415 ;
        RECT 8.185 0.895 8.195 1.425 ;
        RECT 8.195 0.895 8.205 1.435 ;
        RECT 8.205 0.895 8.215 1.445 ;
        RECT 8.215 0.895 8.225 1.455 ;
        RECT 8.225 0.895 8.235 1.465 ;
        RECT 8.235 0.895 8.245 1.475 ;
        RECT 8.245 0.895 8.255 1.485 ;
        RECT 8.255 0.895 8.265 1.495 ;
        RECT 8.265 0.895 8.275 1.505 ;
        RECT 7.855 2.170 7.865 2.674 ;
        RECT 7.865 2.180 7.875 2.674 ;
        RECT 7.875 2.190 7.885 2.674 ;
        RECT 7.885 2.200 7.895 2.674 ;
        RECT 7.895 2.210 7.905 2.674 ;
        RECT 7.905 2.220 7.915 2.674 ;
        RECT 7.915 2.230 7.925 2.674 ;
        RECT 7.925 2.240 7.935 2.674 ;
        RECT 7.935 2.250 7.945 2.674 ;
        RECT 7.945 2.260 7.955 2.674 ;
        RECT 7.955 2.270 7.965 2.674 ;
        RECT 7.965 2.280 7.975 2.674 ;
        RECT 7.975 2.290 7.985 2.674 ;
        RECT 7.985 2.300 7.995 2.674 ;
        RECT 7.995 2.310 8.005 2.674 ;
        RECT 8.005 2.320 8.015 2.674 ;
        RECT 8.015 2.330 8.025 2.674 ;
        RECT 7.875 0.860 7.885 1.064 ;
        RECT 7.885 0.870 7.895 1.064 ;
        RECT 7.895 0.880 7.905 1.064 ;
        RECT 7.905 0.890 7.915 1.064 ;
        RECT 7.915 0.895 7.921 1.065 ;
        RECT 7.820 2.135 7.830 2.375 ;
        RECT 7.830 2.145 7.840 2.385 ;
        RECT 7.840 2.155 7.850 2.395 ;
        RECT 7.850 2.160 7.856 2.404 ;
        RECT 7.800 0.850 7.810 1.020 ;
        RECT 7.810 0.850 7.820 1.030 ;
        RECT 7.820 0.850 7.830 1.040 ;
        RECT 7.830 0.850 7.840 1.050 ;
        RECT 7.840 0.850 7.846 1.060 ;
        RECT 7.740 2.125 7.750 2.295 ;
        RECT 7.750 2.125 7.760 2.305 ;
        RECT 7.760 2.125 7.770 2.315 ;
        RECT 7.770 2.125 7.780 2.325 ;
        RECT 7.780 2.125 7.790 2.335 ;
        RECT 7.790 2.125 7.800 2.345 ;
        RECT 7.800 2.125 7.810 2.355 ;
        RECT 7.810 2.125 7.820 2.365 ;
        RECT 7.275 0.850 7.285 1.084 ;
        RECT 7.285 0.850 7.295 1.074 ;
        RECT 7.295 0.850 7.305 1.064 ;
        RECT 7.305 0.850 7.315 1.054 ;
        RECT 7.315 0.850 7.325 1.044 ;
        RECT 7.325 0.850 7.335 1.034 ;
        RECT 7.335 0.850 7.345 1.024 ;
        RECT 7.345 0.850 7.351 1.020 ;
        RECT 7.210 0.915 7.220 1.149 ;
        RECT 7.220 0.905 7.230 1.139 ;
        RECT 7.230 0.895 7.240 1.129 ;
        RECT 7.240 0.885 7.250 1.119 ;
        RECT 7.250 0.875 7.260 1.109 ;
        RECT 7.260 0.865 7.270 1.099 ;
        RECT 7.270 0.855 7.276 1.095 ;
        RECT 7.135 0.990 7.145 1.160 ;
        RECT 7.145 0.980 7.155 1.160 ;
        RECT 7.155 0.970 7.165 1.160 ;
        RECT 7.165 0.960 7.175 1.160 ;
        RECT 7.175 0.950 7.185 1.160 ;
        RECT 7.185 0.940 7.195 1.160 ;
        RECT 7.195 0.930 7.205 1.160 ;
        RECT 7.205 0.920 7.211 1.160 ;
  END 
END FFDSHQHD2XHT

MACRO FFDSHQHD1XHT
  CLASS  CORE ;
  FOREIGN FFDSHQHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.840 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.420 0.720 9.740 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.455 2.560 2.050 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.995 ;
        RECT 2.175 -0.300 2.475 1.230 ;
        RECT 4.055 -0.300 4.355 0.995 ;
        RECT 5.300 -0.300 5.600 0.530 ;
        RECT 7.235 -0.300 7.535 0.795 ;
        RECT 8.900 -0.300 9.200 1.055 ;
        RECT 0.000 -0.300 9.840 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.870 1.210 1.130 1.795 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.610 0.710 4.840 1.200 ;
        RECT 4.670 0.710 4.840 1.780 ;
        RECT 4.670 1.610 5.065 1.780 ;
        RECT 5.915 0.545 6.085 0.880 ;
        RECT 4.610 0.710 6.085 0.880 ;
        RECT 5.915 0.545 7.035 0.715 ;
        RECT 4.610 0.710 7.035 0.715 ;
        RECT 6.865 0.545 7.035 1.145 ;
        RECT 7.715 0.755 7.885 1.145 ;
        RECT 6.865 0.975 7.885 1.145 ;
        RECT 7.715 0.755 8.425 0.925 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 1.980 0.340 3.990 ;
        RECT 2.205 3.215 2.505 3.990 ;
        RECT 4.035 3.095 4.335 3.990 ;
        RECT 5.135 3.095 5.435 3.990 ;
        RECT 7.235 2.745 7.535 3.990 ;
        RECT 8.335 2.745 8.635 3.990 ;
        RECT 8.900 2.295 9.200 3.990 ;
        RECT 0.000 3.390 9.840 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.000 1.975 1.170 2.215 ;
        RECT 0.870 2.045 1.170 2.215 ;
        RECT 1.145 0.825 1.480 0.995 ;
        RECT 1.000 1.975 1.480 2.145 ;
        RECT 1.310 0.825 1.480 2.145 ;
        RECT 1.310 1.610 1.540 1.910 ;
        RECT 3.115 2.165 3.285 2.335 ;
        RECT 3.130 0.995 3.300 1.495 ;
        RECT 3.130 1.325 3.415 1.495 ;
        RECT 3.315 1.325 3.415 2.335 ;
        RECT 3.485 1.325 4.150 1.495 ;
        RECT 4.320 1.405 4.330 1.865 ;
        RECT 4.330 1.415 4.340 1.865 ;
        RECT 4.340 1.425 4.350 1.865 ;
        RECT 4.350 1.435 4.360 1.865 ;
        RECT 4.360 1.445 4.370 1.865 ;
        RECT 4.370 1.455 4.380 1.865 ;
        RECT 4.380 1.465 4.390 1.865 ;
        RECT 4.390 1.475 4.400 1.865 ;
        RECT 4.400 1.485 4.410 1.865 ;
        RECT 4.410 1.495 4.420 1.865 ;
        RECT 4.420 1.505 4.430 1.865 ;
        RECT 4.430 1.515 4.440 1.865 ;
        RECT 4.440 1.525 4.450 1.865 ;
        RECT 4.450 1.535 4.460 1.865 ;
        RECT 4.460 1.545 4.470 1.865 ;
        RECT 4.470 1.555 4.480 1.865 ;
        RECT 4.480 1.565 4.490 1.865 ;
        RECT 4.250 1.335 4.260 1.595 ;
        RECT 4.260 1.345 4.270 1.605 ;
        RECT 4.270 1.355 4.280 1.615 ;
        RECT 4.280 1.365 4.290 1.625 ;
        RECT 4.290 1.375 4.300 1.635 ;
        RECT 4.300 1.385 4.310 1.645 ;
        RECT 4.310 1.395 4.320 1.655 ;
        RECT 4.150 1.325 4.160 1.495 ;
        RECT 4.160 1.325 4.170 1.505 ;
        RECT 4.170 1.325 4.180 1.515 ;
        RECT 4.180 1.325 4.190 1.525 ;
        RECT 4.190 1.325 4.200 1.535 ;
        RECT 4.200 1.325 4.210 1.545 ;
        RECT 4.210 1.325 4.220 1.555 ;
        RECT 4.220 1.325 4.230 1.565 ;
        RECT 4.230 1.325 4.240 1.575 ;
        RECT 4.240 1.325 4.250 1.585 ;
        RECT 3.415 1.325 3.425 2.325 ;
        RECT 3.425 1.325 3.435 2.315 ;
        RECT 3.435 1.325 3.445 2.305 ;
        RECT 3.445 1.325 3.455 2.295 ;
        RECT 3.455 1.325 3.465 2.285 ;
        RECT 3.465 1.325 3.475 2.275 ;
        RECT 3.475 1.325 3.485 2.265 ;
        RECT 3.285 2.165 3.295 2.335 ;
        RECT 3.295 2.155 3.305 2.335 ;
        RECT 3.305 2.145 3.315 2.335 ;
        RECT 3.775 1.675 4.075 2.215 ;
        RECT 5.020 1.060 5.190 1.360 ;
        RECT 5.020 1.190 5.760 1.360 ;
        RECT 5.590 1.190 5.760 2.215 ;
        RECT 3.770 2.045 5.760 2.215 ;
        RECT 0.170 1.060 0.340 1.790 ;
        RECT 0.170 1.620 0.690 1.790 ;
        RECT 0.520 1.620 0.690 2.565 ;
        RECT 0.520 2.395 1.230 2.565 ;
        RECT 1.060 2.395 1.230 3.035 ;
        RECT 1.060 2.865 3.640 3.035 ;
        RECT 3.835 2.745 5.785 2.915 ;
        RECT 5.615 2.745 5.785 3.195 ;
        RECT 5.615 3.025 6.335 3.195 ;
        RECT 3.760 2.745 3.770 2.979 ;
        RECT 3.770 2.745 3.780 2.969 ;
        RECT 3.780 2.745 3.790 2.959 ;
        RECT 3.790 2.745 3.800 2.949 ;
        RECT 3.800 2.745 3.810 2.939 ;
        RECT 3.810 2.745 3.820 2.929 ;
        RECT 3.820 2.745 3.830 2.919 ;
        RECT 3.830 2.745 3.836 2.915 ;
        RECT 3.715 2.790 3.725 3.024 ;
        RECT 3.725 2.780 3.735 3.014 ;
        RECT 3.735 2.770 3.745 3.004 ;
        RECT 3.745 2.760 3.755 2.994 ;
        RECT 3.755 2.750 3.761 2.990 ;
        RECT 3.640 2.865 3.650 3.035 ;
        RECT 3.650 2.855 3.660 3.035 ;
        RECT 3.660 2.845 3.670 3.035 ;
        RECT 3.670 2.835 3.680 3.035 ;
        RECT 3.680 2.825 3.690 3.035 ;
        RECT 3.690 2.815 3.700 3.035 ;
        RECT 3.700 2.805 3.710 3.035 ;
        RECT 3.710 2.795 3.716 3.035 ;
        RECT 1.720 0.995 1.890 2.685 ;
        RECT 1.440 2.350 1.890 2.685 ;
        RECT 2.765 0.525 2.935 2.685 ;
        RECT 2.765 1.795 3.135 1.965 ;
        RECT 1.440 2.515 3.490 2.685 ;
        RECT 2.765 0.525 3.595 0.695 ;
        RECT 5.965 1.265 6.135 2.685 ;
        RECT 3.685 2.395 6.135 2.565 ;
        RECT 5.965 1.265 6.335 1.435 ;
        RECT 5.965 2.515 6.780 2.685 ;
        RECT 6.610 2.515 6.780 2.890 ;
        RECT 3.610 2.395 3.620 2.629 ;
        RECT 3.620 2.395 3.630 2.619 ;
        RECT 3.630 2.395 3.640 2.609 ;
        RECT 3.640 2.395 3.650 2.599 ;
        RECT 3.650 2.395 3.660 2.589 ;
        RECT 3.660 2.395 3.670 2.579 ;
        RECT 3.670 2.395 3.680 2.569 ;
        RECT 3.680 2.395 3.686 2.565 ;
        RECT 3.565 2.440 3.575 2.674 ;
        RECT 3.575 2.430 3.585 2.664 ;
        RECT 3.585 2.420 3.595 2.654 ;
        RECT 3.595 2.410 3.605 2.644 ;
        RECT 3.605 2.400 3.611 2.640 ;
        RECT 3.490 2.515 3.500 2.685 ;
        RECT 3.500 2.505 3.510 2.685 ;
        RECT 3.510 2.495 3.520 2.685 ;
        RECT 3.520 2.485 3.530 2.685 ;
        RECT 3.530 2.475 3.540 2.685 ;
        RECT 3.540 2.465 3.550 2.685 ;
        RECT 3.550 2.455 3.560 2.685 ;
        RECT 3.560 2.445 3.566 2.685 ;
        RECT 7.915 1.455 8.085 2.215 ;
        RECT 7.490 2.045 8.085 2.215 ;
        RECT 8.305 1.125 8.475 1.625 ;
        RECT 7.915 1.455 8.475 1.625 ;
        RECT 8.305 1.125 8.605 1.295 ;
        RECT 7.320 1.885 7.330 2.215 ;
        RECT 7.330 1.895 7.340 2.215 ;
        RECT 7.340 1.905 7.350 2.215 ;
        RECT 7.350 1.915 7.360 2.215 ;
        RECT 7.360 1.925 7.370 2.215 ;
        RECT 7.370 1.935 7.380 2.215 ;
        RECT 7.380 1.945 7.390 2.215 ;
        RECT 7.390 1.955 7.400 2.215 ;
        RECT 7.400 1.965 7.410 2.215 ;
        RECT 7.410 1.975 7.420 2.215 ;
        RECT 7.420 1.985 7.430 2.215 ;
        RECT 7.430 1.995 7.440 2.215 ;
        RECT 7.440 2.005 7.450 2.215 ;
        RECT 7.450 2.015 7.460 2.215 ;
        RECT 7.460 2.025 7.470 2.215 ;
        RECT 7.470 2.035 7.480 2.215 ;
        RECT 7.480 2.045 7.490 2.215 ;
        RECT 7.275 1.840 7.285 2.170 ;
        RECT 7.285 1.850 7.295 2.180 ;
        RECT 7.295 1.860 7.305 2.190 ;
        RECT 7.305 1.870 7.315 2.200 ;
        RECT 7.315 1.875 7.321 2.209 ;
        RECT 6.975 1.675 6.985 1.869 ;
        RECT 6.985 1.675 6.995 1.879 ;
        RECT 6.995 1.675 7.005 1.889 ;
        RECT 7.005 1.675 7.015 1.899 ;
        RECT 7.015 1.675 7.025 1.909 ;
        RECT 7.025 1.675 7.035 1.919 ;
        RECT 7.035 1.675 7.045 1.929 ;
        RECT 7.045 1.675 7.055 1.939 ;
        RECT 7.055 1.675 7.065 1.949 ;
        RECT 7.065 1.675 7.075 1.959 ;
        RECT 7.075 1.675 7.085 1.969 ;
        RECT 7.085 1.675 7.095 1.979 ;
        RECT 7.095 1.675 7.105 1.989 ;
        RECT 7.105 1.675 7.115 1.999 ;
        RECT 7.115 1.675 7.125 2.009 ;
        RECT 7.125 1.675 7.135 2.019 ;
        RECT 7.135 1.675 7.145 2.029 ;
        RECT 7.145 1.675 7.155 2.039 ;
        RECT 7.155 1.675 7.165 2.049 ;
        RECT 7.165 1.675 7.175 2.059 ;
        RECT 7.175 1.675 7.185 2.069 ;
        RECT 7.185 1.675 7.195 2.079 ;
        RECT 7.195 1.675 7.205 2.089 ;
        RECT 7.205 1.675 7.215 2.099 ;
        RECT 7.215 1.675 7.225 2.109 ;
        RECT 7.225 1.675 7.235 2.119 ;
        RECT 7.235 1.675 7.245 2.129 ;
        RECT 7.245 1.675 7.255 2.139 ;
        RECT 7.255 1.675 7.265 2.149 ;
        RECT 7.265 1.675 7.275 2.159 ;
        RECT 6.295 0.895 6.685 1.065 ;
        RECT 6.515 0.895 6.685 2.335 ;
        RECT 6.315 2.165 6.865 2.335 ;
        RECT 6.515 1.325 7.690 1.495 ;
        RECT 7.520 1.325 7.690 1.730 ;
        RECT 8.315 1.860 8.485 2.565 ;
        RECT 7.185 2.395 8.485 2.565 ;
        RECT 9.050 1.530 9.220 2.030 ;
        RECT 8.315 1.860 9.220 2.030 ;
        RECT 7.095 2.315 7.105 2.565 ;
        RECT 7.105 2.325 7.115 2.565 ;
        RECT 7.115 2.335 7.125 2.565 ;
        RECT 7.125 2.345 7.135 2.565 ;
        RECT 7.135 2.355 7.145 2.565 ;
        RECT 7.145 2.365 7.155 2.565 ;
        RECT 7.155 2.375 7.165 2.565 ;
        RECT 7.165 2.385 7.175 2.565 ;
        RECT 7.175 2.395 7.185 2.565 ;
        RECT 6.955 2.175 6.965 2.425 ;
        RECT 6.965 2.185 6.975 2.435 ;
        RECT 6.975 2.195 6.985 2.445 ;
        RECT 6.985 2.205 6.995 2.455 ;
        RECT 6.995 2.215 7.005 2.465 ;
        RECT 7.005 2.225 7.015 2.475 ;
        RECT 7.015 2.235 7.025 2.485 ;
        RECT 7.025 2.245 7.035 2.495 ;
        RECT 7.035 2.255 7.045 2.505 ;
        RECT 7.045 2.265 7.055 2.515 ;
        RECT 7.055 2.275 7.065 2.525 ;
        RECT 7.065 2.285 7.075 2.535 ;
        RECT 7.075 2.295 7.085 2.545 ;
        RECT 7.085 2.305 7.095 2.555 ;
        RECT 6.865 2.165 6.875 2.335 ;
        RECT 6.875 2.165 6.885 2.345 ;
        RECT 6.885 2.165 6.895 2.355 ;
        RECT 6.895 2.165 6.905 2.365 ;
        RECT 6.905 2.165 6.915 2.375 ;
        RECT 6.915 2.165 6.925 2.385 ;
        RECT 6.925 2.165 6.935 2.395 ;
        RECT 6.935 2.165 6.945 2.405 ;
        RECT 6.945 2.165 6.955 2.415 ;
  END 
END FFDSHQHD1XHT

MACRO FFEDQHD1XHT
  CLASS  CORE ;
  FOREIGN FFEDQHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.320 0.720 10.560 1.360 ;
        RECT 10.350 0.720 10.560 2.960 ;
        RECT 10.320 1.980 10.560 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 1.325 1.220 2.005 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.540 0.620 2.015 ;
        RECT 0.385 2.665 2.215 2.835 ;
        RECT 1.915 2.665 2.215 3.180 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.775 -0.300 1.075 0.710 ;
        RECT 2.535 -0.300 2.835 0.520 ;
        RECT 3.475 -0.300 3.775 0.520 ;
        RECT 5.930 -0.300 6.230 0.525 ;
        RECT 6.910 -0.300 7.210 0.565 ;
        RECT 8.800 -0.300 9.100 0.470 ;
        RECT 9.770 -0.300 9.940 0.710 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.900 1.525 3.485 1.950 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.735 3.035 1.035 3.990 ;
        RECT 2.685 2.840 3.665 3.990 ;
        RECT 6.115 3.160 7.095 3.990 ;
        RECT 8.810 2.830 9.110 3.990 ;
        RECT 9.735 2.975 10.035 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.205 0.975 1.600 1.145 ;
        RECT 1.430 0.975 1.600 2.430 ;
        RECT 0.205 2.260 1.600 2.430 ;
        RECT 1.430 1.705 1.700 2.005 ;
        RECT 3.045 1.125 3.845 1.295 ;
        RECT 3.665 1.125 3.845 2.300 ;
        RECT 3.045 2.130 3.845 2.300 ;
        RECT 3.665 1.525 3.940 1.825 ;
        RECT 4.025 1.065 4.325 1.235 ;
        RECT 4.120 1.065 4.300 2.280 ;
        RECT 4.090 1.980 4.300 2.280 ;
        RECT 4.120 1.065 4.325 1.850 ;
        RECT 4.120 1.550 4.420 1.850 ;
        RECT 1.780 0.945 2.225 1.245 ;
        RECT 2.055 0.945 2.225 2.485 ;
        RECT 1.780 2.185 2.225 2.485 ;
        RECT 2.620 2.305 2.790 2.660 ;
        RECT 1.780 2.305 2.790 2.485 ;
        RECT 4.615 1.060 4.785 2.660 ;
        RECT 2.620 2.480 4.785 2.660 ;
        RECT 4.535 1.060 4.835 1.230 ;
        RECT 5.165 1.060 5.335 2.280 ;
        RECT 5.100 1.060 5.400 1.230 ;
        RECT 6.300 1.675 6.600 1.930 ;
        RECT 5.165 1.760 6.600 1.930 ;
        RECT 5.820 1.325 6.120 1.540 ;
        RECT 6.510 1.125 6.810 1.495 ;
        RECT 5.820 1.325 7.320 1.495 ;
        RECT 7.150 1.325 7.320 2.280 ;
        RECT 6.480 2.110 7.320 2.280 ;
        RECT 5.535 2.810 5.705 3.145 ;
        RECT 3.845 2.975 5.705 3.145 ;
        RECT 5.535 2.810 7.900 2.980 ;
        RECT 4.965 2.460 5.135 2.770 ;
        RECT 7.500 1.310 7.670 2.630 ;
        RECT 7.500 1.310 7.900 1.480 ;
        RECT 4.965 2.460 8.355 2.630 ;
        RECT 8.185 2.460 8.355 2.970 ;
        RECT 2.510 0.700 2.680 1.825 ;
        RECT 2.510 0.700 5.735 0.880 ;
        RECT 5.620 0.765 7.620 0.890 ;
        RECT 5.630 0.765 7.620 0.900 ;
        RECT 5.640 0.765 7.620 0.910 ;
        RECT 5.650 0.765 7.620 0.920 ;
        RECT 5.660 0.765 7.620 0.930 ;
        RECT 5.670 0.765 7.620 0.940 ;
        RECT 5.675 0.700 5.735 0.945 ;
        RECT 2.510 0.710 5.745 0.880 ;
        RECT 2.510 0.720 5.755 0.880 ;
        RECT 2.510 0.730 5.765 0.880 ;
        RECT 2.510 0.740 5.775 0.880 ;
        RECT 2.510 0.750 5.785 0.880 ;
        RECT 5.675 0.765 7.620 0.944 ;
        RECT 2.510 0.760 5.795 0.880 ;
        RECT 7.450 0.575 7.620 0.945 ;
        RECT 5.795 0.765 7.620 0.945 ;
        RECT 7.450 0.575 8.620 0.760 ;
        RECT 8.450 0.575 8.620 1.480 ;
        RECT 8.450 1.310 9.665 1.480 ;
        RECT 9.335 0.875 9.505 1.480 ;
        RECT 9.495 1.310 9.665 2.215 ;
        RECT 9.240 2.045 9.665 2.215 ;
        RECT 7.850 0.940 8.250 1.110 ;
        RECT 8.080 0.940 8.250 2.215 ;
        RECT 7.850 2.045 8.250 2.215 ;
        RECT 8.890 1.675 9.060 2.650 ;
        RECT 8.080 1.675 9.315 1.845 ;
        RECT 9.970 1.520 10.140 2.650 ;
        RECT 8.890 2.480 10.140 2.650 ;
        RECT 9.970 1.520 10.160 1.820 ;
  END 
END FFEDQHD1XHT

MACRO FFEDHQHD3XHT
  CLASS  CORE ;
  FOREIGN FFEDHQHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.680 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 18.170 0.720 18.340 1.360 ;
        RECT 18.170 1.980 18.340 2.960 ;
        RECT 18.170 1.190 19.380 1.360 ;
        RECT 18.170 1.980 19.380 2.150 ;
        RECT 19.210 0.720 19.380 2.960 ;
        RECT 19.210 1.675 19.580 2.015 ;
        RECT 18.170 1.980 19.580 2.015 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.765 0.510 1.395 0.775 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.510 2.015 ;
        RECT 1.060 1.325 1.230 1.625 ;
        RECT 1.060 1.325 2.595 1.495 ;
        RECT 0.520 2.745 2.170 2.915 ;
        RECT 2.000 2.745 2.170 3.110 ;
        RECT 2.000 2.940 4.645 3.110 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.170 -0.300 0.340 1.360 ;
        RECT 1.685 -0.300 1.985 0.435 ;
        RECT 5.255 -0.300 6.235 0.435 ;
        RECT 7.175 -0.300 7.475 0.435 ;
        RECT 8.145 -0.300 8.445 0.435 ;
        RECT 11.545 -0.300 11.845 0.435 ;
        RECT 12.525 -0.300 12.825 0.435 ;
        RECT 13.585 -0.300 13.885 0.435 ;
        RECT 16.735 -0.300 17.035 0.595 ;
        RECT 17.585 -0.300 17.885 0.715 ;
        RECT 18.625 -0.300 18.925 0.715 ;
        RECT 0.000 -0.300 19.680 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 7.005 1.315 7.435 1.660 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.170 2.210 0.340 3.990 ;
        RECT 1.520 3.095 1.820 3.990 ;
        RECT 5.255 2.990 5.895 3.990 ;
        RECT 8.725 3.255 9.025 3.990 ;
        RECT 11.665 3.255 11.965 3.990 ;
        RECT 12.525 3.255 12.825 3.990 ;
        RECT 13.595 2.975 13.895 3.990 ;
        RECT 16.735 2.990 17.035 3.990 ;
        RECT 17.585 2.975 17.885 3.990 ;
        RECT 18.625 2.635 18.925 3.990 ;
        RECT 0.000 3.390 19.680 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 1.060 0.860 2.390 ;
        RECT 0.690 1.805 2.490 1.975 ;
        RECT 2.320 1.740 2.490 2.040 ;
        RECT 2.245 0.540 2.415 1.125 ;
        RECT 1.135 0.955 2.415 1.125 ;
        RECT 2.245 0.540 3.390 0.710 ;
        RECT 3.220 0.540 3.390 1.190 ;
        RECT 1.135 2.265 2.520 2.435 ;
        RECT 2.350 2.265 2.520 2.760 ;
        RECT 3.155 2.495 3.455 2.760 ;
        RECT 2.350 2.590 3.455 2.760 ;
        RECT 3.730 2.430 3.900 2.760 ;
        RECT 4.770 2.330 4.940 2.760 ;
        RECT 3.730 2.590 4.940 2.760 ;
        RECT 4.770 2.330 5.920 2.500 ;
        RECT 5.750 2.330 5.920 2.630 ;
        RECT 3.730 0.540 3.900 1.190 ;
        RECT 3.730 0.540 4.940 0.710 ;
        RECT 4.770 0.540 4.940 1.190 ;
        RECT 5.750 0.890 5.920 1.190 ;
        RECT 4.770 1.020 5.920 1.190 ;
        RECT 7.660 0.985 7.830 2.140 ;
        RECT 7.595 0.985 7.895 1.155 ;
        RECT 7.595 1.970 7.895 2.140 ;
        RECT 7.660 1.355 8.645 1.525 ;
        RECT 2.635 0.955 3.030 1.125 ;
        RECT 2.700 2.110 2.870 2.410 ;
        RECT 2.860 0.955 3.030 2.280 ;
        RECT 2.700 2.110 3.030 2.280 ;
        RECT 2.860 1.675 4.420 1.845 ;
        RECT 4.250 0.890 4.420 2.410 ;
        RECT 4.250 1.940 6.365 2.110 ;
        RECT 6.195 1.940 6.365 3.190 ;
        RECT 6.195 3.020 8.430 3.190 ;
        RECT 8.620 2.905 9.115 3.075 ;
        RECT 9.325 3.040 9.675 3.210 ;
        RECT 9.250 2.975 9.260 3.209 ;
        RECT 9.260 2.985 9.270 3.209 ;
        RECT 9.270 2.995 9.280 3.209 ;
        RECT 9.280 3.005 9.290 3.209 ;
        RECT 9.290 3.015 9.300 3.209 ;
        RECT 9.300 3.025 9.310 3.209 ;
        RECT 9.310 3.035 9.320 3.209 ;
        RECT 9.320 3.040 9.326 3.210 ;
        RECT 9.190 2.915 9.200 3.149 ;
        RECT 9.200 2.925 9.210 3.159 ;
        RECT 9.210 2.935 9.220 3.169 ;
        RECT 9.220 2.945 9.230 3.179 ;
        RECT 9.230 2.955 9.240 3.189 ;
        RECT 9.240 2.965 9.250 3.199 ;
        RECT 9.115 2.905 9.125 3.075 ;
        RECT 9.125 2.905 9.135 3.085 ;
        RECT 9.135 2.905 9.145 3.095 ;
        RECT 9.145 2.905 9.155 3.105 ;
        RECT 9.155 2.905 9.165 3.115 ;
        RECT 9.165 2.905 9.175 3.125 ;
        RECT 9.175 2.905 9.185 3.135 ;
        RECT 9.185 2.905 9.191 3.145 ;
        RECT 8.545 2.905 8.555 3.139 ;
        RECT 8.555 2.905 8.565 3.129 ;
        RECT 8.565 2.905 8.575 3.119 ;
        RECT 8.575 2.905 8.585 3.109 ;
        RECT 8.585 2.905 8.595 3.099 ;
        RECT 8.595 2.905 8.605 3.089 ;
        RECT 8.605 2.905 8.615 3.079 ;
        RECT 8.615 2.905 8.621 3.075 ;
        RECT 8.505 2.945 8.515 3.179 ;
        RECT 8.515 2.935 8.525 3.169 ;
        RECT 8.525 2.925 8.535 3.159 ;
        RECT 8.535 2.915 8.545 3.149 ;
        RECT 8.430 3.020 8.440 3.190 ;
        RECT 8.440 3.010 8.450 3.190 ;
        RECT 8.450 3.000 8.460 3.190 ;
        RECT 8.460 2.990 8.470 3.190 ;
        RECT 8.470 2.980 8.480 3.190 ;
        RECT 8.480 2.970 8.490 3.190 ;
        RECT 8.490 2.960 8.500 3.190 ;
        RECT 8.500 2.950 8.506 3.190 ;
        RECT 10.260 1.185 10.430 2.275 ;
        RECT 9.765 1.965 10.430 2.135 ;
        RECT 10.195 1.185 10.495 1.355 ;
        RECT 10.225 2.105 10.525 2.275 ;
        RECT 9.645 0.985 9.895 1.155 ;
        RECT 10.120 0.835 10.575 1.005 ;
        RECT 10.820 0.985 10.980 2.340 ;
        RECT 10.820 0.985 11.045 1.155 ;
        RECT 11.980 1.520 12.150 1.920 ;
        RECT 10.820 1.750 12.150 1.920 ;
        RECT 10.810 0.985 10.820 2.339 ;
        RECT 10.725 0.900 10.735 1.154 ;
        RECT 10.735 0.910 10.745 1.154 ;
        RECT 10.745 0.920 10.755 1.154 ;
        RECT 10.755 0.930 10.765 1.154 ;
        RECT 10.765 0.940 10.775 1.154 ;
        RECT 10.775 0.950 10.785 1.154 ;
        RECT 10.785 0.960 10.795 1.154 ;
        RECT 10.795 0.970 10.805 1.154 ;
        RECT 10.805 0.975 10.811 1.155 ;
        RECT 10.670 0.845 10.680 1.099 ;
        RECT 10.680 0.855 10.690 1.109 ;
        RECT 10.690 0.865 10.700 1.119 ;
        RECT 10.700 0.875 10.710 1.129 ;
        RECT 10.710 0.885 10.720 1.139 ;
        RECT 10.720 0.890 10.726 1.150 ;
        RECT 10.575 0.835 10.585 1.005 ;
        RECT 10.585 0.835 10.595 1.015 ;
        RECT 10.595 0.835 10.605 1.025 ;
        RECT 10.605 0.835 10.615 1.035 ;
        RECT 10.615 0.835 10.625 1.045 ;
        RECT 10.625 0.835 10.635 1.055 ;
        RECT 10.635 0.835 10.645 1.065 ;
        RECT 10.645 0.835 10.655 1.075 ;
        RECT 10.655 0.835 10.665 1.085 ;
        RECT 10.665 0.835 10.671 1.095 ;
        RECT 10.045 0.835 10.055 1.069 ;
        RECT 10.055 0.835 10.065 1.059 ;
        RECT 10.065 0.835 10.075 1.049 ;
        RECT 10.075 0.835 10.085 1.039 ;
        RECT 10.085 0.835 10.095 1.029 ;
        RECT 10.095 0.835 10.105 1.019 ;
        RECT 10.105 0.835 10.115 1.009 ;
        RECT 10.115 0.835 10.121 1.005 ;
        RECT 9.970 0.910 9.980 1.144 ;
        RECT 9.980 0.900 9.990 1.134 ;
        RECT 9.990 0.890 10.000 1.124 ;
        RECT 10.000 0.880 10.010 1.114 ;
        RECT 10.010 0.870 10.020 1.104 ;
        RECT 10.020 0.860 10.030 1.094 ;
        RECT 10.030 0.850 10.040 1.084 ;
        RECT 10.040 0.840 10.046 1.080 ;
        RECT 9.895 0.985 9.905 1.155 ;
        RECT 9.905 0.975 9.915 1.155 ;
        RECT 9.915 0.965 9.925 1.155 ;
        RECT 9.925 0.955 9.935 1.155 ;
        RECT 9.935 0.945 9.945 1.155 ;
        RECT 9.945 0.935 9.955 1.155 ;
        RECT 9.955 0.925 9.965 1.155 ;
        RECT 9.965 0.915 9.971 1.155 ;
        RECT 11.470 1.030 11.640 1.570 ;
        RECT 11.405 1.400 11.705 1.570 ;
        RECT 11.470 1.030 12.500 1.200 ;
        RECT 12.330 1.030 12.500 2.315 ;
        RECT 12.095 2.145 12.500 2.315 ;
        RECT 12.330 1.515 14.015 1.685 ;
        RECT 13.035 2.215 15.535 2.385 ;
        RECT 13.035 1.030 14.390 1.200 ;
        RECT 14.660 0.835 15.110 1.005 ;
        RECT 15.175 0.835 15.185 1.070 ;
        RECT 15.250 0.900 15.585 1.070 ;
        RECT 15.185 0.845 15.195 1.069 ;
        RECT 15.195 0.855 15.205 1.069 ;
        RECT 15.205 0.865 15.215 1.069 ;
        RECT 15.215 0.875 15.225 1.069 ;
        RECT 15.225 0.885 15.235 1.069 ;
        RECT 15.235 0.895 15.245 1.069 ;
        RECT 15.245 0.900 15.251 1.070 ;
        RECT 15.110 0.835 15.120 1.005 ;
        RECT 15.120 0.835 15.130 1.015 ;
        RECT 15.130 0.835 15.140 1.025 ;
        RECT 15.140 0.835 15.150 1.035 ;
        RECT 15.150 0.835 15.160 1.045 ;
        RECT 15.160 0.835 15.170 1.055 ;
        RECT 15.170 0.835 15.176 1.065 ;
        RECT 14.585 0.835 14.595 1.069 ;
        RECT 14.595 0.835 14.605 1.059 ;
        RECT 14.605 0.835 14.615 1.049 ;
        RECT 14.615 0.835 14.625 1.039 ;
        RECT 14.625 0.835 14.635 1.029 ;
        RECT 14.635 0.835 14.645 1.019 ;
        RECT 14.645 0.835 14.655 1.009 ;
        RECT 14.655 0.835 14.661 1.005 ;
        RECT 14.535 0.885 14.545 1.119 ;
        RECT 14.545 0.875 14.555 1.109 ;
        RECT 14.555 0.865 14.565 1.099 ;
        RECT 14.565 0.855 14.575 1.089 ;
        RECT 14.575 0.845 14.585 1.079 ;
        RECT 14.390 1.030 14.400 1.200 ;
        RECT 14.400 1.020 14.410 1.200 ;
        RECT 14.410 1.010 14.420 1.200 ;
        RECT 14.420 1.000 14.430 1.200 ;
        RECT 14.430 0.990 14.440 1.200 ;
        RECT 14.440 0.980 14.450 1.200 ;
        RECT 14.450 0.970 14.460 1.200 ;
        RECT 14.460 0.960 14.470 1.200 ;
        RECT 14.470 0.950 14.480 1.200 ;
        RECT 14.480 0.940 14.490 1.200 ;
        RECT 14.490 0.930 14.500 1.200 ;
        RECT 14.500 0.920 14.510 1.200 ;
        RECT 14.510 0.910 14.520 1.200 ;
        RECT 14.520 0.900 14.530 1.200 ;
        RECT 14.530 0.890 14.536 1.200 ;
        RECT 6.625 0.965 6.795 2.840 ;
        RECT 6.625 0.965 6.925 1.135 ;
        RECT 6.625 2.670 8.255 2.840 ;
        RECT 8.445 2.555 9.270 2.725 ;
        RECT 9.480 2.690 9.760 2.860 ;
        RECT 13.205 2.625 13.375 3.075 ;
        RECT 10.055 2.905 13.375 3.075 ;
        RECT 13.205 2.625 14.295 2.795 ;
        RECT 14.125 2.625 14.295 3.085 ;
        RECT 14.125 2.915 15.905 3.085 ;
        RECT 9.975 2.835 9.985 3.075 ;
        RECT 9.985 2.845 9.995 3.075 ;
        RECT 9.995 2.855 10.005 3.075 ;
        RECT 10.005 2.865 10.015 3.075 ;
        RECT 10.015 2.875 10.025 3.075 ;
        RECT 10.025 2.885 10.035 3.075 ;
        RECT 10.035 2.895 10.045 3.075 ;
        RECT 10.045 2.905 10.055 3.075 ;
        RECT 9.840 2.700 9.850 2.940 ;
        RECT 9.850 2.710 9.860 2.950 ;
        RECT 9.860 2.720 9.870 2.960 ;
        RECT 9.870 2.730 9.880 2.970 ;
        RECT 9.880 2.740 9.890 2.980 ;
        RECT 9.890 2.750 9.900 2.990 ;
        RECT 9.900 2.760 9.910 3.000 ;
        RECT 9.910 2.770 9.920 3.010 ;
        RECT 9.920 2.780 9.930 3.020 ;
        RECT 9.930 2.790 9.940 3.030 ;
        RECT 9.940 2.800 9.950 3.040 ;
        RECT 9.950 2.810 9.960 3.050 ;
        RECT 9.960 2.820 9.970 3.060 ;
        RECT 9.970 2.825 9.976 3.069 ;
        RECT 9.760 2.690 9.770 2.860 ;
        RECT 9.770 2.690 9.780 2.870 ;
        RECT 9.780 2.690 9.790 2.880 ;
        RECT 9.790 2.690 9.800 2.890 ;
        RECT 9.800 2.690 9.810 2.900 ;
        RECT 9.810 2.690 9.820 2.910 ;
        RECT 9.820 2.690 9.830 2.920 ;
        RECT 9.830 2.690 9.840 2.930 ;
        RECT 9.405 2.625 9.415 2.859 ;
        RECT 9.415 2.635 9.425 2.859 ;
        RECT 9.425 2.645 9.435 2.859 ;
        RECT 9.435 2.655 9.445 2.859 ;
        RECT 9.445 2.665 9.455 2.859 ;
        RECT 9.455 2.675 9.465 2.859 ;
        RECT 9.465 2.685 9.475 2.859 ;
        RECT 9.475 2.690 9.481 2.860 ;
        RECT 9.345 2.565 9.355 2.799 ;
        RECT 9.355 2.575 9.365 2.809 ;
        RECT 9.365 2.585 9.375 2.819 ;
        RECT 9.375 2.595 9.385 2.829 ;
        RECT 9.385 2.605 9.395 2.839 ;
        RECT 9.395 2.615 9.405 2.849 ;
        RECT 9.270 2.555 9.280 2.725 ;
        RECT 9.280 2.555 9.290 2.735 ;
        RECT 9.290 2.555 9.300 2.745 ;
        RECT 9.300 2.555 9.310 2.755 ;
        RECT 9.310 2.555 9.320 2.765 ;
        RECT 9.320 2.555 9.330 2.775 ;
        RECT 9.330 2.555 9.340 2.785 ;
        RECT 9.340 2.555 9.346 2.795 ;
        RECT 8.370 2.555 8.380 2.789 ;
        RECT 8.380 2.555 8.390 2.779 ;
        RECT 8.390 2.555 8.400 2.769 ;
        RECT 8.400 2.555 8.410 2.759 ;
        RECT 8.410 2.555 8.420 2.749 ;
        RECT 8.420 2.555 8.430 2.739 ;
        RECT 8.430 2.555 8.440 2.729 ;
        RECT 8.440 2.555 8.446 2.725 ;
        RECT 8.330 2.595 8.340 2.829 ;
        RECT 8.340 2.585 8.350 2.819 ;
        RECT 8.350 2.575 8.360 2.809 ;
        RECT 8.360 2.565 8.370 2.799 ;
        RECT 8.255 2.670 8.265 2.840 ;
        RECT 8.265 2.660 8.275 2.840 ;
        RECT 8.275 2.650 8.285 2.840 ;
        RECT 8.285 2.640 8.295 2.840 ;
        RECT 8.295 2.630 8.305 2.840 ;
        RECT 8.305 2.620 8.315 2.840 ;
        RECT 8.315 2.610 8.325 2.840 ;
        RECT 8.325 2.600 8.331 2.840 ;
        RECT 7.095 1.900 7.265 2.490 ;
        RECT 7.095 2.320 8.055 2.490 ;
        RECT 8.685 0.985 9.015 1.155 ;
        RECT 8.845 0.985 9.015 2.310 ;
        RECT 8.310 2.140 9.360 2.310 ;
        RECT 8.845 1.315 9.375 1.485 ;
        RECT 9.635 2.340 9.925 2.510 ;
        RECT 12.680 1.865 12.850 2.725 ;
        RECT 10.220 2.555 12.850 2.725 ;
        RECT 14.385 1.380 14.555 2.035 ;
        RECT 12.680 1.865 16.295 2.035 ;
        RECT 10.140 2.485 10.150 2.725 ;
        RECT 10.150 2.495 10.160 2.725 ;
        RECT 10.160 2.505 10.170 2.725 ;
        RECT 10.170 2.515 10.180 2.725 ;
        RECT 10.180 2.525 10.190 2.725 ;
        RECT 10.190 2.535 10.200 2.725 ;
        RECT 10.200 2.545 10.210 2.725 ;
        RECT 10.210 2.555 10.220 2.725 ;
        RECT 10.005 2.350 10.015 2.590 ;
        RECT 10.015 2.360 10.025 2.600 ;
        RECT 10.025 2.370 10.035 2.610 ;
        RECT 10.035 2.380 10.045 2.620 ;
        RECT 10.045 2.390 10.055 2.630 ;
        RECT 10.055 2.400 10.065 2.640 ;
        RECT 10.065 2.410 10.075 2.650 ;
        RECT 10.075 2.420 10.085 2.660 ;
        RECT 10.085 2.430 10.095 2.670 ;
        RECT 10.095 2.440 10.105 2.680 ;
        RECT 10.105 2.450 10.115 2.690 ;
        RECT 10.115 2.460 10.125 2.700 ;
        RECT 10.125 2.470 10.135 2.710 ;
        RECT 10.135 2.475 10.141 2.719 ;
        RECT 9.925 2.340 9.935 2.510 ;
        RECT 9.935 2.340 9.945 2.520 ;
        RECT 9.945 2.340 9.955 2.530 ;
        RECT 9.955 2.340 9.965 2.540 ;
        RECT 9.965 2.340 9.975 2.550 ;
        RECT 9.975 2.340 9.985 2.560 ;
        RECT 9.985 2.340 9.995 2.570 ;
        RECT 9.995 2.340 10.005 2.580 ;
        RECT 9.560 2.275 9.570 2.509 ;
        RECT 9.570 2.285 9.580 2.509 ;
        RECT 9.580 2.295 9.590 2.509 ;
        RECT 9.590 2.305 9.600 2.509 ;
        RECT 9.600 2.315 9.610 2.509 ;
        RECT 9.610 2.325 9.620 2.509 ;
        RECT 9.620 2.335 9.630 2.509 ;
        RECT 9.630 2.340 9.636 2.510 ;
        RECT 9.435 2.150 9.445 2.384 ;
        RECT 9.445 2.160 9.455 2.394 ;
        RECT 9.455 2.170 9.465 2.404 ;
        RECT 9.465 2.180 9.475 2.414 ;
        RECT 9.475 2.190 9.485 2.424 ;
        RECT 9.485 2.200 9.495 2.434 ;
        RECT 9.495 2.210 9.505 2.444 ;
        RECT 9.505 2.220 9.515 2.454 ;
        RECT 9.515 2.230 9.525 2.464 ;
        RECT 9.525 2.240 9.535 2.474 ;
        RECT 9.535 2.250 9.545 2.484 ;
        RECT 9.545 2.260 9.555 2.494 ;
        RECT 9.555 2.265 9.561 2.505 ;
        RECT 9.360 2.140 9.370 2.310 ;
        RECT 9.370 2.140 9.380 2.320 ;
        RECT 9.380 2.140 9.390 2.330 ;
        RECT 9.390 2.140 9.400 2.340 ;
        RECT 9.400 2.140 9.410 2.350 ;
        RECT 9.410 2.140 9.420 2.360 ;
        RECT 9.420 2.140 9.430 2.370 ;
        RECT 9.430 2.140 9.436 2.380 ;
        RECT 8.235 2.140 8.245 2.374 ;
        RECT 8.245 2.140 8.255 2.364 ;
        RECT 8.255 2.140 8.265 2.354 ;
        RECT 8.265 2.140 8.275 2.344 ;
        RECT 8.275 2.140 8.285 2.334 ;
        RECT 8.285 2.140 8.295 2.324 ;
        RECT 8.295 2.140 8.305 2.314 ;
        RECT 8.305 2.140 8.311 2.310 ;
        RECT 8.130 2.245 8.140 2.479 ;
        RECT 8.140 2.235 8.150 2.469 ;
        RECT 8.150 2.225 8.160 2.459 ;
        RECT 8.160 2.215 8.170 2.449 ;
        RECT 8.170 2.205 8.180 2.439 ;
        RECT 8.180 2.195 8.190 2.429 ;
        RECT 8.190 2.185 8.200 2.419 ;
        RECT 8.200 2.175 8.210 2.409 ;
        RECT 8.210 2.165 8.220 2.399 ;
        RECT 8.220 2.155 8.230 2.389 ;
        RECT 8.230 2.145 8.236 2.385 ;
        RECT 8.055 2.320 8.065 2.490 ;
        RECT 8.065 2.310 8.075 2.490 ;
        RECT 8.075 2.300 8.085 2.490 ;
        RECT 8.085 2.290 8.095 2.490 ;
        RECT 8.095 2.280 8.105 2.490 ;
        RECT 8.105 2.270 8.115 2.490 ;
        RECT 8.115 2.260 8.125 2.490 ;
        RECT 8.125 2.250 8.131 2.490 ;
        RECT 6.100 0.615 6.270 1.755 ;
        RECT 5.045 1.585 6.270 1.755 ;
        RECT 6.100 0.615 9.760 0.785 ;
        RECT 9.970 0.480 10.775 0.650 ;
        RECT 10.985 0.615 14.300 0.785 ;
        RECT 14.515 0.480 15.260 0.650 ;
        RECT 15.330 0.480 15.335 0.720 ;
        RECT 16.255 0.480 16.555 0.720 ;
        RECT 15.405 0.550 16.555 0.720 ;
        RECT 16.385 0.480 16.555 0.985 ;
        RECT 16.385 0.815 17.400 0.985 ;
        RECT 17.230 0.815 17.400 2.405 ;
        RECT 17.165 2.235 17.465 2.405 ;
        RECT 15.335 0.490 15.345 0.720 ;
        RECT 15.345 0.500 15.355 0.720 ;
        RECT 15.355 0.510 15.365 0.720 ;
        RECT 15.365 0.520 15.375 0.720 ;
        RECT 15.375 0.530 15.385 0.720 ;
        RECT 15.385 0.540 15.395 0.720 ;
        RECT 15.395 0.550 15.405 0.720 ;
        RECT 15.260 0.480 15.270 0.650 ;
        RECT 15.270 0.480 15.280 0.660 ;
        RECT 15.280 0.480 15.290 0.670 ;
        RECT 15.290 0.480 15.300 0.680 ;
        RECT 15.300 0.480 15.310 0.690 ;
        RECT 15.310 0.480 15.320 0.700 ;
        RECT 15.320 0.480 15.330 0.710 ;
        RECT 14.435 0.480 14.445 0.720 ;
        RECT 14.445 0.480 14.455 0.710 ;
        RECT 14.455 0.480 14.465 0.700 ;
        RECT 14.465 0.480 14.475 0.690 ;
        RECT 14.475 0.480 14.485 0.680 ;
        RECT 14.485 0.480 14.495 0.670 ;
        RECT 14.495 0.480 14.505 0.660 ;
        RECT 14.505 0.480 14.515 0.650 ;
        RECT 14.380 0.535 14.390 0.775 ;
        RECT 14.390 0.525 14.400 0.765 ;
        RECT 14.400 0.515 14.410 0.755 ;
        RECT 14.410 0.505 14.420 0.745 ;
        RECT 14.420 0.495 14.430 0.735 ;
        RECT 14.430 0.485 14.436 0.729 ;
        RECT 14.300 0.615 14.310 0.785 ;
        RECT 14.310 0.605 14.320 0.785 ;
        RECT 14.320 0.595 14.330 0.785 ;
        RECT 14.330 0.585 14.340 0.785 ;
        RECT 14.340 0.575 14.350 0.785 ;
        RECT 14.350 0.565 14.360 0.785 ;
        RECT 14.360 0.555 14.370 0.785 ;
        RECT 14.370 0.545 14.380 0.785 ;
        RECT 10.910 0.550 10.920 0.784 ;
        RECT 10.920 0.560 10.930 0.784 ;
        RECT 10.930 0.570 10.940 0.784 ;
        RECT 10.940 0.580 10.950 0.784 ;
        RECT 10.950 0.590 10.960 0.784 ;
        RECT 10.960 0.600 10.970 0.784 ;
        RECT 10.970 0.610 10.980 0.784 ;
        RECT 10.980 0.615 10.986 0.785 ;
        RECT 10.850 0.490 10.860 0.724 ;
        RECT 10.860 0.500 10.870 0.734 ;
        RECT 10.870 0.510 10.880 0.744 ;
        RECT 10.880 0.520 10.890 0.754 ;
        RECT 10.890 0.530 10.900 0.764 ;
        RECT 10.900 0.540 10.910 0.774 ;
        RECT 10.775 0.480 10.785 0.650 ;
        RECT 10.785 0.480 10.795 0.660 ;
        RECT 10.795 0.480 10.805 0.670 ;
        RECT 10.805 0.480 10.815 0.680 ;
        RECT 10.815 0.480 10.825 0.690 ;
        RECT 10.825 0.480 10.835 0.700 ;
        RECT 10.835 0.480 10.845 0.710 ;
        RECT 10.845 0.480 10.851 0.720 ;
        RECT 9.895 0.480 9.905 0.714 ;
        RECT 9.905 0.480 9.915 0.704 ;
        RECT 9.915 0.480 9.925 0.694 ;
        RECT 9.925 0.480 9.935 0.684 ;
        RECT 9.935 0.480 9.945 0.674 ;
        RECT 9.945 0.480 9.955 0.664 ;
        RECT 9.955 0.480 9.965 0.654 ;
        RECT 9.965 0.480 9.971 0.650 ;
        RECT 9.835 0.540 9.845 0.774 ;
        RECT 9.845 0.530 9.855 0.764 ;
        RECT 9.855 0.520 9.865 0.754 ;
        RECT 9.865 0.510 9.875 0.744 ;
        RECT 9.875 0.500 9.885 0.734 ;
        RECT 9.885 0.490 9.895 0.724 ;
        RECT 9.760 0.615 9.770 0.785 ;
        RECT 9.770 0.605 9.780 0.785 ;
        RECT 9.780 0.595 9.790 0.785 ;
        RECT 9.790 0.585 9.800 0.785 ;
        RECT 9.800 0.575 9.810 0.785 ;
        RECT 9.810 0.565 9.820 0.785 ;
        RECT 9.820 0.555 9.830 0.785 ;
        RECT 9.830 0.545 9.836 0.785 ;
        RECT 14.865 1.185 15.035 1.485 ;
        RECT 14.735 1.185 15.035 1.355 ;
        RECT 15.815 1.175 15.985 1.485 ;
        RECT 14.865 1.315 15.985 1.485 ;
        RECT 15.880 2.215 16.050 2.735 ;
        RECT 14.685 2.565 16.050 2.735 ;
        RECT 15.815 1.175 16.835 1.345 ;
        RECT 15.880 2.215 16.835 2.385 ;
        RECT 16.665 1.175 16.835 2.795 ;
        RECT 17.645 1.575 17.815 2.795 ;
        RECT 16.665 2.625 17.815 2.795 ;
        RECT 17.645 1.575 18.905 1.745 ;
  END 
END FFEDHQHD3XHT

MACRO FFEDHQHD2XHT
  CLASS  CORE ;
  FOREIGN FFEDHQHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.040 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 17.040 0.720 17.210 1.405 ;
        RECT 17.040 1.980 17.210 2.960 ;
        RECT 17.040 1.235 17.940 1.405 ;
        RECT 17.730 1.235 17.940 2.150 ;
        RECT 17.040 1.980 17.940 2.150 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 0.510 1.505 0.855 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.510 2.015 ;
        RECT 0.520 2.745 2.170 2.915 ;
        RECT 2.000 2.745 2.170 3.090 ;
        RECT 2.000 2.920 4.645 3.090 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.170 -0.300 0.340 1.360 ;
        RECT 1.685 -0.300 1.985 0.745 ;
        RECT 5.255 -0.300 6.235 0.435 ;
        RECT 7.180 -0.300 8.160 0.435 ;
        RECT 10.565 -0.300 12.225 0.435 ;
        RECT 15.515 -0.300 15.815 0.595 ;
        RECT 16.455 -0.300 16.755 1.055 ;
        RECT 17.495 -0.300 17.795 1.055 ;
        RECT 0.000 -0.300 18.040 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 7.070 1.265 7.370 1.685 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.170 2.210 0.340 3.990 ;
        RECT 1.520 3.095 1.820 3.990 ;
        RECT 5.255 2.990 6.170 3.990 ;
        RECT 10.565 3.255 12.665 3.990 ;
        RECT 15.515 2.990 15.815 3.990 ;
        RECT 16.455 2.975 16.755 3.990 ;
        RECT 17.495 2.635 17.795 3.990 ;
        RECT 0.000 3.390 18.040 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 1.060 0.860 2.390 ;
        RECT 0.690 1.785 2.520 1.955 ;
        RECT 2.350 1.720 2.520 2.020 ;
        RECT 1.135 2.265 2.520 2.435 ;
        RECT 2.350 2.265 2.520 2.740 ;
        RECT 3.220 2.390 3.390 2.740 ;
        RECT 2.350 2.570 3.390 2.740 ;
        RECT 2.245 0.710 2.415 1.295 ;
        RECT 1.135 1.125 2.415 1.295 ;
        RECT 2.245 0.710 3.390 0.880 ;
        RECT 3.220 0.710 3.390 1.360 ;
        RECT 3.730 2.390 3.900 2.740 ;
        RECT 4.770 2.330 4.940 2.740 ;
        RECT 3.730 2.570 4.940 2.740 ;
        RECT 4.770 2.330 5.920 2.500 ;
        RECT 5.750 2.330 5.920 2.630 ;
        RECT 3.730 0.530 3.900 1.180 ;
        RECT 3.730 0.530 4.940 0.700 ;
        RECT 4.770 0.530 4.940 1.180 ;
        RECT 5.750 0.880 5.920 1.180 ;
        RECT 4.770 1.010 5.920 1.180 ;
        RECT 7.630 0.965 7.800 2.140 ;
        RECT 7.565 0.965 7.865 1.135 ;
        RECT 7.565 1.970 7.865 2.140 ;
        RECT 7.630 1.335 8.525 1.505 ;
        RECT 2.700 1.060 2.870 2.390 ;
        RECT 2.700 1.675 4.420 1.845 ;
        RECT 4.250 0.880 4.420 2.390 ;
        RECT 4.250 1.945 6.350 2.115 ;
        RECT 6.810 3.040 7.615 3.210 ;
        RECT 7.635 3.020 7.690 3.210 ;
        RECT 7.710 3.020 8.595 3.190 ;
        RECT 8.615 3.020 8.670 3.210 ;
        RECT 8.690 3.040 9.385 3.210 ;
        RECT 8.670 3.030 8.680 3.210 ;
        RECT 8.680 3.040 8.690 3.210 ;
        RECT 8.595 3.020 8.605 3.190 ;
        RECT 8.605 3.020 8.615 3.200 ;
        RECT 7.690 3.020 7.700 3.200 ;
        RECT 7.700 3.020 7.710 3.190 ;
        RECT 7.615 3.040 7.625 3.210 ;
        RECT 7.625 3.030 7.635 3.210 ;
        RECT 6.695 2.935 6.705 3.209 ;
        RECT 6.705 2.945 6.715 3.209 ;
        RECT 6.715 2.955 6.725 3.209 ;
        RECT 6.725 2.965 6.735 3.209 ;
        RECT 6.735 2.975 6.745 3.209 ;
        RECT 6.745 2.985 6.755 3.209 ;
        RECT 6.755 2.995 6.765 3.209 ;
        RECT 6.765 3.005 6.775 3.209 ;
        RECT 6.775 3.015 6.785 3.209 ;
        RECT 6.785 3.025 6.795 3.209 ;
        RECT 6.795 3.035 6.805 3.209 ;
        RECT 6.805 3.040 6.811 3.210 ;
        RECT 6.520 2.760 6.530 3.034 ;
        RECT 6.530 2.770 6.540 3.044 ;
        RECT 6.540 2.780 6.550 3.054 ;
        RECT 6.550 2.790 6.560 3.064 ;
        RECT 6.560 2.800 6.570 3.074 ;
        RECT 6.570 2.810 6.580 3.084 ;
        RECT 6.580 2.820 6.590 3.094 ;
        RECT 6.590 2.830 6.600 3.104 ;
        RECT 6.600 2.840 6.610 3.114 ;
        RECT 6.610 2.850 6.620 3.124 ;
        RECT 6.620 2.860 6.630 3.134 ;
        RECT 6.630 2.870 6.640 3.144 ;
        RECT 6.640 2.880 6.650 3.154 ;
        RECT 6.650 2.890 6.660 3.164 ;
        RECT 6.660 2.900 6.670 3.174 ;
        RECT 6.670 2.910 6.680 3.184 ;
        RECT 6.680 2.920 6.690 3.194 ;
        RECT 6.690 2.925 6.696 3.205 ;
        RECT 6.350 1.945 6.360 2.865 ;
        RECT 6.360 1.945 6.370 2.875 ;
        RECT 6.370 1.945 6.380 2.885 ;
        RECT 6.380 1.945 6.390 2.895 ;
        RECT 6.390 1.945 6.400 2.905 ;
        RECT 6.400 1.945 6.410 2.915 ;
        RECT 6.410 1.945 6.420 2.925 ;
        RECT 6.420 1.945 6.430 2.935 ;
        RECT 6.430 1.945 6.440 2.945 ;
        RECT 6.440 1.945 6.450 2.955 ;
        RECT 6.450 1.945 6.460 2.965 ;
        RECT 6.460 1.945 6.470 2.975 ;
        RECT 6.470 1.945 6.480 2.985 ;
        RECT 6.480 1.945 6.490 2.995 ;
        RECT 6.490 1.945 6.500 3.005 ;
        RECT 6.500 1.945 6.510 3.015 ;
        RECT 6.510 1.945 6.520 3.025 ;
        RECT 9.190 0.920 9.360 2.155 ;
        RECT 9.085 1.985 9.385 2.155 ;
        RECT 9.710 0.920 9.880 2.155 ;
        RECT 9.710 1.770 9.915 2.155 ;
        RECT 9.615 1.985 9.915 2.155 ;
        RECT 10.880 1.520 11.050 1.940 ;
        RECT 9.710 1.770 11.050 1.940 ;
        RECT 10.370 0.985 10.540 1.590 ;
        RECT 10.370 0.985 11.400 1.155 ;
        RECT 11.230 0.985 11.400 2.315 ;
        RECT 10.995 2.145 11.400 2.315 ;
        RECT 11.230 1.535 12.575 1.705 ;
        RECT 11.935 2.535 14.255 2.705 ;
        RECT 12.915 0.875 13.215 1.155 ;
        RECT 11.935 0.985 13.215 1.155 ;
        RECT 13.860 0.875 14.030 1.065 ;
        RECT 12.915 0.875 14.030 1.045 ;
        RECT 13.860 0.895 14.335 1.065 ;
        RECT 6.625 0.965 6.710 1.135 ;
        RECT 6.880 0.965 6.925 1.135 ;
        RECT 6.880 1.970 7.295 2.140 ;
        RECT 6.990 2.690 7.450 2.860 ;
        RECT 7.470 2.670 7.540 2.860 ;
        RECT 7.560 2.670 8.750 2.840 ;
        RECT 8.770 2.670 8.840 2.860 ;
        RECT 9.955 2.690 10.125 3.025 ;
        RECT 8.860 2.690 10.125 2.860 ;
        RECT 11.585 2.855 11.755 3.055 ;
        RECT 9.955 2.855 11.755 3.025 ;
        RECT 11.585 2.885 14.555 3.055 ;
        RECT 14.385 2.885 14.555 3.075 ;
        RECT 14.385 2.905 14.685 3.075 ;
        RECT 8.840 2.680 8.850 2.860 ;
        RECT 8.850 2.690 8.860 2.860 ;
        RECT 8.750 2.670 8.760 2.840 ;
        RECT 8.760 2.670 8.770 2.850 ;
        RECT 7.540 2.670 7.550 2.850 ;
        RECT 7.550 2.670 7.560 2.840 ;
        RECT 7.450 2.690 7.460 2.860 ;
        RECT 7.460 2.680 7.470 2.860 ;
        RECT 6.915 2.625 6.925 2.859 ;
        RECT 6.925 2.635 6.935 2.859 ;
        RECT 6.935 2.645 6.945 2.859 ;
        RECT 6.945 2.655 6.955 2.859 ;
        RECT 6.955 2.665 6.965 2.859 ;
        RECT 6.965 2.675 6.975 2.859 ;
        RECT 6.975 2.685 6.985 2.859 ;
        RECT 6.985 2.690 6.991 2.860 ;
        RECT 6.880 2.590 6.890 2.824 ;
        RECT 6.890 2.600 6.900 2.834 ;
        RECT 6.900 2.610 6.910 2.844 ;
        RECT 6.910 2.615 6.916 2.855 ;
        RECT 6.710 0.965 6.720 2.655 ;
        RECT 6.720 0.965 6.730 2.665 ;
        RECT 6.730 0.965 6.740 2.675 ;
        RECT 6.740 0.965 6.750 2.685 ;
        RECT 6.750 0.965 6.760 2.695 ;
        RECT 6.760 0.965 6.770 2.705 ;
        RECT 6.770 0.965 6.780 2.715 ;
        RECT 6.780 0.965 6.790 2.725 ;
        RECT 6.790 0.965 6.800 2.735 ;
        RECT 6.800 0.965 6.810 2.745 ;
        RECT 6.810 0.965 6.820 2.755 ;
        RECT 6.820 0.965 6.830 2.765 ;
        RECT 6.830 0.965 6.840 2.775 ;
        RECT 6.840 0.965 6.850 2.785 ;
        RECT 6.850 0.965 6.860 2.795 ;
        RECT 6.860 0.965 6.870 2.805 ;
        RECT 6.870 0.965 6.880 2.815 ;
        RECT 7.070 2.320 7.370 2.510 ;
        RECT 8.610 1.665 8.780 2.490 ;
        RECT 8.545 0.965 8.955 1.135 ;
        RECT 8.930 2.340 10.695 2.500 ;
        RECT 8.785 0.965 8.955 1.835 ;
        RECT 8.610 1.665 8.955 1.835 ;
        RECT 8.785 1.270 8.990 1.570 ;
        RECT 7.070 2.320 8.995 2.490 ;
        RECT 7.070 2.330 9.005 2.490 ;
        RECT 10.525 2.340 10.695 2.675 ;
        RECT 8.940 2.340 10.695 2.510 ;
        RECT 11.585 1.885 11.755 2.675 ;
        RECT 10.525 2.505 11.755 2.675 ;
        RECT 13.120 1.460 13.290 2.055 ;
        RECT 11.585 1.885 13.290 2.055 ;
        RECT 13.120 1.815 15.075 1.985 ;
        RECT 6.110 0.615 6.280 1.755 ;
        RECT 5.045 1.585 6.280 1.755 ;
        RECT 8.655 0.505 8.825 0.785 ;
        RECT 6.110 0.615 8.825 0.785 ;
        RECT 8.655 0.505 10.290 0.675 ;
        RECT 10.120 0.505 10.290 0.805 ;
        RECT 12.485 0.500 12.655 0.805 ;
        RECT 10.120 0.635 12.655 0.805 ;
        RECT 12.485 0.500 14.690 0.670 ;
        RECT 14.520 0.500 14.690 0.945 ;
        RECT 14.520 0.775 16.180 0.945 ;
        RECT 16.010 0.775 16.180 2.355 ;
        RECT 15.945 2.185 16.245 2.355 ;
        RECT 13.615 1.245 13.785 1.520 ;
        RECT 13.485 1.245 13.785 1.415 ;
        RECT 14.595 1.125 14.765 1.520 ;
        RECT 13.615 1.350 14.765 1.520 ;
        RECT 14.595 1.125 15.615 1.295 ;
        RECT 13.435 2.185 15.615 2.355 ;
        RECT 15.445 1.125 15.615 2.760 ;
        RECT 16.450 1.585 16.620 2.760 ;
        RECT 15.445 2.590 16.620 2.760 ;
        RECT 16.450 1.585 17.435 1.755 ;
  END 
END FFEDHQHD2XHT

MACRO FFEDHQHD1XHT
  CLASS  CORE ;
  FOREIGN FFEDHQHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.890 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.415 0.720 11.585 2.960 ;
        RECT 11.415 1.675 11.790 2.075 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.865 1.260 1.130 2.000 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.585 2.020 ;
        RECT 0.285 2.645 1.365 2.815 ;
        RECT 1.195 2.645 1.365 3.210 ;
        RECT 1.195 3.040 2.075 3.210 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.730 ;
        RECT 2.415 -0.300 2.715 0.435 ;
        RECT 4.210 -0.300 4.510 0.435 ;
        RECT 6.960 -0.300 7.260 0.435 ;
        RECT 8.020 -0.300 8.320 0.435 ;
        RECT 9.890 -0.300 10.190 0.565 ;
        RECT 10.830 -0.300 11.130 1.055 ;
        RECT 0.000 -0.300 11.890 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 3.505 1.330 4.140 1.570 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.995 0.955 3.990 ;
        RECT 2.515 3.040 2.815 3.990 ;
        RECT 5.275 3.255 5.575 3.990 ;
        RECT 7.080 3.205 7.380 3.990 ;
        RECT 8.020 3.205 8.320 3.990 ;
        RECT 9.890 2.995 10.190 3.990 ;
        RECT 10.800 2.995 11.100 3.990 ;
        RECT 0.000 3.390 11.890 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.910 0.340 1.360 ;
        RECT 0.170 0.910 1.480 1.080 ;
        RECT 1.310 0.910 1.480 2.445 ;
        RECT 0.105 2.275 1.480 2.445 ;
        RECT 1.310 1.785 1.645 1.955 ;
        RECT 2.720 1.125 2.890 2.445 ;
        RECT 2.720 1.125 3.265 1.295 ;
        RECT 2.720 2.275 3.600 2.445 ;
        RECT 3.430 2.210 3.600 2.510 ;
        RECT 3.640 0.965 4.490 1.135 ;
        RECT 4.320 0.965 4.490 2.055 ;
        RECT 4.130 1.885 4.490 2.055 ;
        RECT 4.320 1.335 5.090 1.505 ;
        RECT 3.155 1.785 3.950 1.955 ;
        RECT 3.780 1.785 3.950 2.405 ;
        RECT 4.670 1.685 4.840 2.405 ;
        RECT 3.780 2.235 4.840 2.405 ;
        RECT 4.760 0.965 5.455 1.135 ;
        RECT 5.195 1.685 5.365 2.120 ;
        RECT 5.275 0.965 5.455 1.865 ;
        RECT 4.670 1.685 5.455 1.865 ;
        RECT 5.275 1.270 5.510 1.570 ;
        RECT 1.660 1.060 1.995 1.360 ;
        RECT 1.660 2.165 1.995 2.465 ;
        RECT 1.825 1.060 1.995 2.860 ;
        RECT 1.825 2.690 3.715 2.860 ;
        RECT 3.735 2.670 3.820 2.860 ;
        RECT 3.840 2.670 4.840 2.840 ;
        RECT 5.545 2.155 5.715 2.725 ;
        RECT 5.035 2.555 5.715 2.725 ;
        RECT 5.705 0.965 5.875 2.325 ;
        RECT 5.640 0.965 5.940 1.135 ;
        RECT 5.545 2.155 5.940 2.325 ;
        RECT 4.955 2.555 4.965 2.795 ;
        RECT 4.965 2.555 4.975 2.785 ;
        RECT 4.975 2.555 4.985 2.775 ;
        RECT 4.985 2.555 4.995 2.765 ;
        RECT 4.995 2.555 5.005 2.755 ;
        RECT 5.005 2.555 5.015 2.745 ;
        RECT 5.015 2.555 5.025 2.735 ;
        RECT 5.025 2.555 5.035 2.725 ;
        RECT 4.920 2.590 4.930 2.830 ;
        RECT 4.930 2.580 4.940 2.820 ;
        RECT 4.940 2.570 4.950 2.810 ;
        RECT 4.950 2.560 4.956 2.804 ;
        RECT 4.840 2.670 4.850 2.840 ;
        RECT 4.850 2.660 4.860 2.840 ;
        RECT 4.860 2.650 4.870 2.840 ;
        RECT 4.870 2.640 4.880 2.840 ;
        RECT 4.880 2.630 4.890 2.840 ;
        RECT 4.890 2.620 4.900 2.840 ;
        RECT 4.900 2.610 4.910 2.840 ;
        RECT 4.910 2.600 4.920 2.840 ;
        RECT 3.820 2.670 3.830 2.850 ;
        RECT 3.830 2.670 3.840 2.840 ;
        RECT 3.715 2.690 3.725 2.860 ;
        RECT 3.725 2.680 3.735 2.860 ;
        RECT 6.225 0.965 6.395 2.325 ;
        RECT 6.160 0.965 6.460 1.135 ;
        RECT 6.160 2.155 6.460 2.325 ;
        RECT 6.225 1.785 7.630 1.955 ;
        RECT 7.575 0.965 7.745 1.605 ;
        RECT 7.510 0.965 7.810 1.135 ;
        RECT 7.810 1.435 7.980 2.325 ;
        RECT 7.510 2.155 7.980 2.325 ;
        RECT 6.840 1.435 8.530 1.605 ;
        RECT 3.365 3.040 3.925 3.210 ;
        RECT 3.945 3.020 4.060 3.210 ;
        RECT 4.080 3.020 5.000 3.190 ;
        RECT 5.195 2.905 5.730 3.075 ;
        RECT 6.500 2.855 6.800 3.195 ;
        RECT 5.930 3.025 6.800 3.195 ;
        RECT 6.500 2.855 9.010 3.025 ;
        RECT 8.710 2.855 9.010 3.195 ;
        RECT 5.850 2.955 5.860 3.195 ;
        RECT 5.860 2.965 5.870 3.195 ;
        RECT 5.870 2.975 5.880 3.195 ;
        RECT 5.880 2.985 5.890 3.195 ;
        RECT 5.890 2.995 5.900 3.195 ;
        RECT 5.900 3.005 5.910 3.195 ;
        RECT 5.910 3.015 5.920 3.195 ;
        RECT 5.920 3.025 5.930 3.195 ;
        RECT 5.810 2.915 5.820 3.155 ;
        RECT 5.820 2.925 5.830 3.165 ;
        RECT 5.830 2.935 5.840 3.175 ;
        RECT 5.840 2.945 5.850 3.185 ;
        RECT 5.730 2.905 5.740 3.075 ;
        RECT 5.740 2.905 5.750 3.085 ;
        RECT 5.750 2.905 5.760 3.095 ;
        RECT 5.760 2.905 5.770 3.105 ;
        RECT 5.770 2.905 5.780 3.115 ;
        RECT 5.780 2.905 5.790 3.125 ;
        RECT 5.790 2.905 5.800 3.135 ;
        RECT 5.800 2.905 5.810 3.145 ;
        RECT 5.115 2.905 5.125 3.145 ;
        RECT 5.125 2.905 5.135 3.135 ;
        RECT 5.135 2.905 5.145 3.125 ;
        RECT 5.145 2.905 5.155 3.115 ;
        RECT 5.155 2.905 5.165 3.105 ;
        RECT 5.165 2.905 5.175 3.095 ;
        RECT 5.175 2.905 5.185 3.085 ;
        RECT 5.185 2.905 5.195 3.075 ;
        RECT 5.080 2.940 5.090 3.180 ;
        RECT 5.090 2.930 5.100 3.170 ;
        RECT 5.100 2.920 5.110 3.160 ;
        RECT 5.110 2.910 5.116 3.154 ;
        RECT 5.000 3.020 5.010 3.190 ;
        RECT 5.010 3.010 5.020 3.190 ;
        RECT 5.020 3.000 5.030 3.190 ;
        RECT 5.030 2.990 5.040 3.190 ;
        RECT 5.040 2.980 5.050 3.190 ;
        RECT 5.050 2.970 5.060 3.190 ;
        RECT 5.060 2.960 5.070 3.190 ;
        RECT 5.070 2.950 5.080 3.190 ;
        RECT 4.060 3.020 4.070 3.200 ;
        RECT 4.070 3.020 4.080 3.190 ;
        RECT 3.925 3.040 3.935 3.210 ;
        RECT 3.935 3.030 3.945 3.210 ;
        RECT 5.980 2.505 6.300 2.815 ;
        RECT 8.590 1.785 8.760 2.675 ;
        RECT 8.710 1.315 8.880 1.955 ;
        RECT 8.590 1.785 8.880 1.955 ;
        RECT 8.710 1.315 9.010 1.485 ;
        RECT 5.980 2.505 9.425 2.675 ;
        RECT 9.255 2.505 9.425 3.195 ;
        RECT 9.190 3.025 9.490 3.195 ;
        RECT 2.370 0.615 2.540 1.820 ;
        RECT 8.545 0.500 8.715 0.785 ;
        RECT 2.370 0.615 8.715 0.785 ;
        RECT 8.545 0.500 9.710 0.670 ;
        RECT 9.540 0.500 9.710 1.755 ;
        RECT 9.540 1.585 10.555 1.755 ;
        RECT 10.385 0.880 10.555 2.465 ;
        RECT 10.320 2.295 10.620 2.465 ;
        RECT 8.940 0.945 9.360 1.115 ;
        RECT 9.190 0.945 9.360 2.305 ;
        RECT 8.940 2.135 10.115 2.305 ;
        RECT 9.935 2.135 10.115 2.815 ;
        RECT 11.000 1.520 11.170 2.815 ;
        RECT 9.935 2.645 11.170 2.815 ;
  END 
END FFEDHQHD1XHT

MACRO FFEDHDMXHT
  CLASS  CORE ;
  FOREIGN FFEDHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.480 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.130 0.970 11.380 1.270 ;
        RECT 11.210 0.970 11.380 2.445 ;
        RECT 11.130 1.980 11.380 2.445 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.940 0.820 10.260 1.205 ;
        RECT 10.090 0.820 10.260 1.470 ;
        RECT 10.090 2.000 10.260 2.300 ;
        RECT 10.090 1.290 10.545 1.470 ;
        RECT 10.345 1.290 10.545 2.235 ;
        RECT 10.090 2.000 10.545 2.235 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 1.325 1.195 2.005 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.545 0.625 2.010 ;
        RECT 0.330 2.695 2.160 2.865 ;
        RECT 1.860 2.695 2.160 3.180 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 -0.300 1.020 0.795 ;
        RECT 2.510 -0.300 2.810 0.520 ;
        RECT 3.480 -0.300 3.780 0.520 ;
        RECT 6.010 -0.300 6.310 0.525 ;
        RECT 7.035 -0.300 7.335 0.565 ;
        RECT 8.935 -0.300 9.235 1.110 ;
        RECT 10.545 -0.300 10.845 1.055 ;
        RECT 0.000 -0.300 11.480 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.970 1.525 3.490 2.015 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 3.045 1.020 3.990 ;
        RECT 2.680 2.905 3.660 3.990 ;
        RECT 6.130 3.160 6.430 3.990 ;
        RECT 7.045 3.160 7.345 3.990 ;
        RECT 8.945 2.830 9.245 3.990 ;
        RECT 10.515 2.925 10.815 3.990 ;
        RECT 0.000 3.390 11.480 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.150 0.975 1.545 1.145 ;
        RECT 1.375 0.975 1.545 2.430 ;
        RECT 0.150 2.260 1.545 2.430 ;
        RECT 1.375 1.705 1.645 2.005 ;
        RECT 3.020 1.125 3.905 1.295 ;
        RECT 3.735 1.125 3.905 2.365 ;
        RECT 2.990 2.195 3.905 2.365 ;
        RECT 3.735 1.525 3.970 1.825 ;
        RECT 4.085 1.125 4.385 1.295 ;
        RECT 4.150 1.125 4.320 2.280 ;
        RECT 4.150 1.125 4.385 1.850 ;
        RECT 4.150 1.550 4.485 1.850 ;
        RECT 1.745 1.045 2.055 1.345 ;
        RECT 1.885 1.045 2.055 2.515 ;
        RECT 1.725 2.215 2.055 2.515 ;
        RECT 1.725 2.345 2.695 2.515 ;
        RECT 2.525 2.345 2.695 2.725 ;
        RECT 4.665 1.060 4.845 2.725 ;
        RECT 2.525 2.545 4.845 2.725 ;
        RECT 4.595 1.060 4.895 1.230 ;
        RECT 5.245 1.060 5.415 2.280 ;
        RECT 5.180 1.060 5.480 1.230 ;
        RECT 6.380 1.675 6.680 1.930 ;
        RECT 5.245 1.760 6.680 1.930 ;
        RECT 5.900 1.325 6.200 1.540 ;
        RECT 6.590 1.125 6.890 1.495 ;
        RECT 5.900 1.325 7.455 1.495 ;
        RECT 7.285 1.325 7.455 2.280 ;
        RECT 6.560 2.110 7.455 2.280 ;
        RECT 5.615 2.810 5.785 3.145 ;
        RECT 3.875 2.975 5.785 3.145 ;
        RECT 5.615 2.810 8.035 2.980 ;
        RECT 5.035 2.460 5.205 2.770 ;
        RECT 7.635 1.310 7.805 2.630 ;
        RECT 7.635 1.310 8.035 1.480 ;
        RECT 5.035 2.460 8.415 2.630 ;
        RECT 8.235 2.460 8.415 2.935 ;
        RECT 8.235 2.765 8.555 2.935 ;
        RECT 2.455 0.700 2.625 1.825 ;
        RECT 5.710 0.700 5.880 0.945 ;
        RECT 2.455 0.700 5.880 0.880 ;
        RECT 7.580 0.575 7.750 0.945 ;
        RECT 5.710 0.765 7.750 0.945 ;
        RECT 7.580 0.575 8.755 0.760 ;
        RECT 8.585 0.575 8.755 1.480 ;
        RECT 9.580 0.875 9.655 1.480 ;
        RECT 8.585 1.310 9.655 1.480 ;
        RECT 9.740 0.875 9.750 2.215 ;
        RECT 9.485 2.045 9.750 2.215 ;
        RECT 9.910 1.650 10.135 1.820 ;
        RECT 9.750 1.320 9.760 2.214 ;
        RECT 9.760 1.330 9.770 2.214 ;
        RECT 9.770 1.340 9.780 2.214 ;
        RECT 9.780 1.350 9.790 2.214 ;
        RECT 9.790 1.360 9.800 2.214 ;
        RECT 9.800 1.370 9.810 2.214 ;
        RECT 9.810 1.380 9.820 2.214 ;
        RECT 9.820 1.390 9.830 2.214 ;
        RECT 9.830 1.400 9.840 2.214 ;
        RECT 9.840 1.410 9.850 2.214 ;
        RECT 9.850 1.420 9.860 2.214 ;
        RECT 9.860 1.430 9.870 2.214 ;
        RECT 9.870 1.440 9.880 2.214 ;
        RECT 9.880 1.450 9.890 2.214 ;
        RECT 9.890 1.460 9.900 2.214 ;
        RECT 9.900 1.470 9.910 2.214 ;
        RECT 9.655 0.875 9.665 1.479 ;
        RECT 9.665 0.875 9.675 1.489 ;
        RECT 9.675 0.875 9.685 1.499 ;
        RECT 9.685 0.875 9.695 1.509 ;
        RECT 9.695 0.875 9.705 1.519 ;
        RECT 9.705 0.875 9.715 1.529 ;
        RECT 9.715 0.875 9.725 1.539 ;
        RECT 9.725 0.875 9.735 1.549 ;
        RECT 9.735 0.875 9.741 1.559 ;
        RECT 7.985 0.940 8.385 1.110 ;
        RECT 8.215 0.940 8.385 2.215 ;
        RECT 7.985 2.045 8.385 2.215 ;
        RECT 9.135 1.675 9.305 2.650 ;
        RECT 8.215 1.675 9.560 1.845 ;
        RECT 10.780 1.520 10.950 2.650 ;
        RECT 9.135 2.480 10.950 2.650 ;
        RECT 10.780 1.520 10.970 1.820 ;
  END 
END FFEDHDMXHT

MACRO FFEDHDLXHT
  CLASS  CORE ;
  FOREIGN FFEDHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.480 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.065 0.885 11.380 1.055 ;
        RECT 11.170 0.885 11.380 2.280 ;
        RECT 11.130 1.980 11.380 2.280 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.940 0.820 10.325 1.195 ;
        RECT 10.090 2.000 10.260 2.300 ;
        RECT 10.145 0.820 10.325 1.470 ;
        RECT 10.145 1.290 10.600 1.470 ;
        RECT 10.430 1.290 10.600 2.170 ;
        RECT 10.090 2.000 10.600 2.170 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 1.325 1.195 2.005 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.575 0.565 2.015 ;
        RECT 0.330 2.665 2.160 2.835 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 -0.300 1.020 0.795 ;
        RECT 2.715 -0.300 3.695 0.520 ;
        RECT 6.205 -0.300 7.185 0.575 ;
        RECT 8.915 -0.300 9.215 0.725 ;
        RECT 10.545 -0.300 10.845 1.055 ;
        RECT 0.000 -0.300 11.480 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.870 1.525 3.555 1.950 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.720 3.015 1.020 3.990 ;
        RECT 2.700 2.840 3.680 3.990 ;
        RECT 6.230 3.160 7.210 3.990 ;
        RECT 8.915 2.830 9.215 3.990 ;
        RECT 10.515 2.830 10.815 3.990 ;
        RECT 0.000 3.390 11.480 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.150 0.975 1.545 1.145 ;
        RECT 1.375 0.975 1.545 2.430 ;
        RECT 0.150 2.260 1.545 2.430 ;
        RECT 1.375 1.705 1.645 2.005 ;
        RECT 3.020 1.125 3.905 1.295 ;
        RECT 3.735 1.125 3.905 2.300 ;
        RECT 2.990 2.130 3.905 2.300 ;
        RECT 3.735 1.525 3.970 1.825 ;
        RECT 4.085 1.125 4.385 1.295 ;
        RECT 4.150 1.125 4.320 2.280 ;
        RECT 4.150 1.125 4.385 1.850 ;
        RECT 4.150 1.550 4.450 1.850 ;
        RECT 1.745 1.045 2.055 1.345 ;
        RECT 1.885 1.045 2.055 2.485 ;
        RECT 1.725 2.185 2.055 2.485 ;
        RECT 2.575 2.315 2.745 2.660 ;
        RECT 1.725 2.315 2.745 2.485 ;
        RECT 4.665 1.060 4.845 2.660 ;
        RECT 2.575 2.480 4.845 2.660 ;
        RECT 4.595 1.060 4.895 1.230 ;
        RECT 5.245 1.060 5.415 2.280 ;
        RECT 5.180 1.060 5.480 1.230 ;
        RECT 6.380 1.675 6.680 1.930 ;
        RECT 5.245 1.760 6.680 1.930 ;
        RECT 5.900 1.325 6.200 1.540 ;
        RECT 6.590 1.125 6.890 1.495 ;
        RECT 5.900 1.325 7.435 1.495 ;
        RECT 7.265 1.325 7.435 2.280 ;
        RECT 6.560 2.110 7.435 2.280 ;
        RECT 3.875 2.840 4.175 3.145 ;
        RECT 5.550 2.810 5.730 3.145 ;
        RECT 3.875 2.975 5.730 3.145 ;
        RECT 5.550 2.810 7.905 2.980 ;
        RECT 5.035 2.460 5.205 2.770 ;
        RECT 7.615 1.310 7.785 2.630 ;
        RECT 7.615 1.310 8.015 1.480 ;
        RECT 5.035 2.460 8.420 2.630 ;
        RECT 8.250 2.460 8.420 2.885 ;
        RECT 2.455 0.700 2.625 1.825 ;
        RECT 5.680 0.700 5.850 0.945 ;
        RECT 2.455 0.700 5.850 0.880 ;
        RECT 7.490 0.555 7.660 0.945 ;
        RECT 5.680 0.765 7.660 0.945 ;
        RECT 7.490 0.555 8.735 0.740 ;
        RECT 8.565 0.555 8.735 1.480 ;
        RECT 9.560 0.855 9.660 1.480 ;
        RECT 8.565 1.310 9.660 1.480 ;
        RECT 9.720 0.855 9.730 2.215 ;
        RECT 9.720 1.310 9.750 2.215 ;
        RECT 9.465 2.045 9.750 2.215 ;
        RECT 9.890 1.650 10.250 1.820 ;
        RECT 9.750 1.320 9.760 2.214 ;
        RECT 9.760 1.330 9.770 2.214 ;
        RECT 9.770 1.340 9.780 2.214 ;
        RECT 9.780 1.350 9.790 2.214 ;
        RECT 9.790 1.360 9.800 2.214 ;
        RECT 9.800 1.370 9.810 2.214 ;
        RECT 9.810 1.380 9.820 2.214 ;
        RECT 9.820 1.390 9.830 2.214 ;
        RECT 9.830 1.400 9.840 2.214 ;
        RECT 9.840 1.410 9.850 2.214 ;
        RECT 9.850 1.420 9.860 2.214 ;
        RECT 9.860 1.430 9.870 2.214 ;
        RECT 9.870 1.440 9.880 2.214 ;
        RECT 9.880 1.450 9.890 2.214 ;
        RECT 9.660 0.855 9.670 1.479 ;
        RECT 9.670 0.855 9.680 1.489 ;
        RECT 9.680 0.855 9.690 1.499 ;
        RECT 9.690 0.855 9.700 1.509 ;
        RECT 9.700 0.855 9.710 1.519 ;
        RECT 9.710 0.855 9.720 1.529 ;
        RECT 7.965 0.920 8.365 1.090 ;
        RECT 8.195 0.920 8.365 2.215 ;
        RECT 7.965 2.045 8.365 2.215 ;
        RECT 8.970 1.675 9.140 2.650 ;
        RECT 8.195 1.675 9.540 1.845 ;
        RECT 10.780 1.520 10.950 2.650 ;
        RECT 8.970 2.480 10.950 2.650 ;
        RECT 10.780 1.520 10.970 1.820 ;
  END 
END FFEDHDLXHT

MACRO FFEDHD2XHT
  CLASS  CORE ;
  FOREIGN FFEDHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.710 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.200 2.045 11.500 2.555 ;
        RECT 11.200 1.125 11.795 1.295 ;
        RECT 11.615 1.125 11.795 2.425 ;
        RECT 11.200 2.045 11.795 2.425 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.100 1.125 10.560 1.295 ;
        RECT 10.350 0.775 10.560 2.215 ;
        RECT 10.100 2.045 10.560 2.215 ;
        RECT 10.350 0.775 12.535 0.945 ;
        RECT 12.365 0.720 12.535 2.960 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.875 1.265 1.130 2.015 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.675 0.605 2.015 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.675 -0.300 0.975 0.735 ;
        RECT 2.435 -0.300 2.735 0.525 ;
        RECT 3.495 -0.300 3.795 0.525 ;
        RECT 5.860 -0.300 6.160 0.525 ;
        RECT 6.830 -0.300 7.130 0.565 ;
        RECT 9.040 -0.300 9.340 0.470 ;
        RECT 10.650 -0.300 10.950 0.595 ;
        RECT 11.750 -0.300 12.050 0.595 ;
        RECT 0.000 -0.300 12.710 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.870 1.525 3.425 1.950 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.685 2.640 0.985 3.990 ;
        RECT 2.585 2.905 3.565 3.990 ;
        RECT 6.060 3.160 7.040 3.990 ;
        RECT 8.955 2.765 9.255 3.990 ;
        RECT 10.650 3.095 10.950 3.990 ;
        RECT 11.750 3.095 12.050 3.990 ;
        RECT 0.000 3.390 12.710 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 0.915 0.405 1.145 ;
        RECT 0.105 0.915 1.500 1.085 ;
        RECT 1.330 0.915 1.500 2.430 ;
        RECT 0.105 2.260 1.500 2.430 ;
        RECT 1.330 1.705 1.600 2.005 ;
        RECT 2.945 1.125 3.775 1.295 ;
        RECT 3.605 1.125 3.775 2.300 ;
        RECT 2.945 2.130 3.775 2.300 ;
        RECT 3.605 1.525 3.840 1.825 ;
        RECT 3.955 1.125 4.255 1.295 ;
        RECT 4.020 1.125 4.190 2.280 ;
        RECT 4.020 1.125 4.255 1.850 ;
        RECT 4.020 1.550 4.320 1.850 ;
        RECT 1.680 0.945 2.010 1.245 ;
        RECT 1.840 0.945 2.010 2.875 ;
        RECT 1.680 2.235 2.010 2.875 ;
        RECT 4.535 1.980 4.705 2.725 ;
        RECT 1.680 2.545 4.705 2.725 ;
        RECT 4.545 1.060 4.715 2.380 ;
        RECT 4.535 1.980 4.715 2.380 ;
        RECT 4.465 1.060 4.765 1.230 ;
        RECT 5.095 1.060 5.265 2.280 ;
        RECT 5.030 1.060 5.330 1.230 ;
        RECT 6.230 1.675 6.530 1.930 ;
        RECT 5.095 1.760 6.530 1.930 ;
        RECT 5.750 1.325 6.050 1.540 ;
        RECT 6.440 1.125 6.740 1.495 ;
        RECT 5.750 1.325 7.245 1.495 ;
        RECT 7.075 1.325 7.245 2.280 ;
        RECT 6.410 2.110 7.245 2.280 ;
        RECT 4.885 2.460 5.055 2.770 ;
        RECT 4.885 2.460 8.305 2.630 ;
        RECT 8.135 2.460 8.305 2.795 ;
        RECT 3.745 2.975 4.045 3.185 ;
        RECT 5.465 2.810 5.635 3.145 ;
        RECT 3.745 2.975 5.635 3.145 ;
        RECT 5.465 2.810 7.850 2.980 ;
        RECT 7.680 2.810 7.850 3.210 ;
        RECT 8.220 1.350 8.665 1.520 ;
        RECT 8.485 1.350 8.665 3.210 ;
        RECT 7.680 3.040 8.665 3.210 ;
        RECT 2.410 0.710 2.580 1.825 ;
        RECT 2.410 0.710 5.695 0.880 ;
        RECT 5.570 0.765 7.560 0.890 ;
        RECT 5.580 0.765 7.560 0.900 ;
        RECT 5.590 0.765 7.560 0.910 ;
        RECT 5.600 0.765 7.560 0.920 ;
        RECT 5.610 0.765 7.560 0.930 ;
        RECT 5.620 0.765 7.560 0.940 ;
        RECT 5.625 0.710 5.695 0.945 ;
        RECT 2.410 0.720 5.705 0.880 ;
        RECT 2.410 0.730 5.715 0.880 ;
        RECT 2.410 0.740 5.725 0.880 ;
        RECT 2.410 0.750 5.735 0.880 ;
        RECT 5.625 0.765 7.560 0.944 ;
        RECT 2.410 0.760 5.745 0.880 ;
        RECT 7.390 0.650 7.560 0.945 ;
        RECT 5.745 0.765 7.560 0.945 ;
        RECT 8.540 0.480 8.840 0.820 ;
        RECT 7.390 0.650 9.635 0.820 ;
        RECT 9.465 0.650 9.635 1.295 ;
        RECT 9.465 1.125 9.920 1.295 ;
        RECT 9.750 1.125 9.920 2.215 ;
        RECT 9.560 2.045 9.920 2.215 ;
        RECT 9.750 1.650 10.170 1.820 ;
        RECT 7.760 1.000 7.940 2.240 ;
        RECT 7.760 2.070 8.080 2.240 ;
        RECT 7.760 1.000 9.090 1.170 ;
        RECT 8.920 1.000 9.090 1.815 ;
        RECT 9.210 1.645 9.380 2.565 ;
        RECT 8.920 1.645 9.570 1.815 ;
        RECT 10.800 1.605 10.970 2.565 ;
        RECT 9.210 2.395 10.970 2.565 ;
        RECT 10.800 1.605 11.435 1.775 ;
        RECT 10.115 2.745 10.285 3.210 ;
        RECT 9.820 3.040 10.285 3.210 ;
        RECT 12.015 1.585 12.185 2.915 ;
        RECT 10.115 2.745 12.185 2.915 ;
  END 
END FFEDHD2XHT

MACRO FFEDHD1XHT
  CLASS  CORE ;
  FOREIGN FFEDHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.480 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.130 0.720 11.300 2.960 ;
        RECT 11.130 2.040 11.380 2.445 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.870 0.510 10.325 0.720 ;
        RECT 10.090 2.000 10.260 2.300 ;
        RECT 10.090 0.510 10.325 1.470 ;
        RECT 10.090 1.290 10.545 1.470 ;
        RECT 10.345 1.290 10.545 2.235 ;
        RECT 10.090 2.000 10.545 2.235 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 1.325 1.220 2.005 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.625 0.620 2.015 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.775 -0.300 1.075 0.795 ;
        RECT 2.750 -0.300 3.730 0.525 ;
        RECT 6.250 -0.300 7.230 0.575 ;
        RECT 8.935 -0.300 9.235 1.110 ;
        RECT 10.610 -0.300 10.780 1.120 ;
        RECT 0.000 -0.300 11.480 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 2.970 1.525 3.555 2.015 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.785 2.640 1.085 3.990 ;
        RECT 2.715 2.905 3.695 3.990 ;
        RECT 6.265 3.160 7.245 3.990 ;
        RECT 8.945 2.830 9.245 3.990 ;
        RECT 10.545 2.975 10.845 3.990 ;
        RECT 0.000 3.390 11.480 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.205 0.975 1.600 1.145 ;
        RECT 1.430 0.975 1.600 2.430 ;
        RECT 0.205 2.260 1.600 2.430 ;
        RECT 1.430 1.770 1.765 1.940 ;
        RECT 3.045 1.125 3.905 1.295 ;
        RECT 3.735 1.125 3.905 2.365 ;
        RECT 3.045 2.195 3.905 2.365 ;
        RECT 3.735 1.525 3.970 1.825 ;
        RECT 4.085 1.125 4.385 1.295 ;
        RECT 4.150 1.125 4.320 2.280 ;
        RECT 4.150 1.125 4.385 1.850 ;
        RECT 4.150 1.550 4.450 1.850 ;
        RECT 1.780 2.120 1.950 2.760 ;
        RECT 1.780 0.945 2.255 1.245 ;
        RECT 2.085 0.945 2.255 2.725 ;
        RECT 1.780 2.120 2.255 2.725 ;
        RECT 4.675 1.060 4.845 2.725 ;
        RECT 1.780 2.545 4.845 2.725 ;
        RECT 4.595 1.060 4.895 1.230 ;
        RECT 5.245 1.060 5.415 2.280 ;
        RECT 5.180 1.060 5.480 1.230 ;
        RECT 6.380 1.675 6.680 1.930 ;
        RECT 5.245 1.760 6.680 1.930 ;
        RECT 5.900 1.325 6.200 1.540 ;
        RECT 6.590 1.125 6.890 1.495 ;
        RECT 5.900 1.325 7.455 1.495 ;
        RECT 7.285 1.325 7.455 2.280 ;
        RECT 6.560 2.110 7.455 2.280 ;
        RECT 5.550 2.810 5.850 3.120 ;
        RECT 3.875 2.950 5.850 3.120 ;
        RECT 5.550 2.810 8.035 2.980 ;
        RECT 5.035 2.460 5.205 2.770 ;
        RECT 7.635 1.310 7.805 2.630 ;
        RECT 7.635 1.310 8.035 1.480 ;
        RECT 5.035 2.460 8.490 2.630 ;
        RECT 8.320 2.460 8.490 2.945 ;
        RECT 2.510 0.705 2.680 1.825 ;
        RECT 2.510 0.705 4.295 0.885 ;
        RECT 4.300 0.705 4.320 0.880 ;
        RECT 4.325 0.700 5.860 0.880 ;
        RECT 5.690 0.700 5.860 0.945 ;
        RECT 2.510 0.705 5.860 0.879 ;
        RECT 7.580 0.575 7.750 0.945 ;
        RECT 5.690 0.765 7.750 0.945 ;
        RECT 7.580 0.575 8.735 0.760 ;
        RECT 8.565 0.575 8.735 1.480 ;
        RECT 8.565 1.310 9.910 1.480 ;
        RECT 9.580 0.875 9.750 1.480 ;
        RECT 9.740 1.310 9.910 2.215 ;
        RECT 9.485 2.045 9.910 2.215 ;
        RECT 9.740 1.650 10.135 1.820 ;
        RECT 7.985 0.940 8.385 1.110 ;
        RECT 8.215 0.940 8.385 2.215 ;
        RECT 7.985 2.045 8.385 2.215 ;
        RECT 9.135 1.675 9.305 2.650 ;
        RECT 8.215 1.675 9.560 1.845 ;
        RECT 10.780 1.520 10.950 2.650 ;
        RECT 9.135 2.480 10.950 2.650 ;
  END 
END FFEDHD1XHT

MACRO FFEDCRHDMXHT
  CLASS  CORE ;
  FOREIGN FFEDCRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.530 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.055 0.955 13.225 2.620 ;
        RECT 13.055 1.645 13.255 2.620 ;
        RECT 13.055 1.645 13.430 2.040 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.985 0.805 12.200 1.480 ;
        RECT 11.985 1.300 12.470 1.480 ;
        RECT 12.270 1.300 12.470 2.215 ;
        RECT 11.950 2.045 12.470 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.595 2.970 2.355 3.210 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.215 2.560 0.830 2.770 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.620 1.560 2.800 2.430 ;
        RECT 2.510 2.085 2.800 2.430 ;
        RECT 2.620 1.560 3.020 1.860 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.750 ;
        RECT 2.510 -0.300 2.680 0.810 ;
        RECT 3.535 -0.300 4.555 0.555 ;
        RECT 5.550 -0.300 6.530 0.555 ;
        RECT 8.205 -0.300 8.505 0.575 ;
        RECT 9.185 -0.300 9.355 0.890 ;
        RECT 10.990 -0.300 11.290 0.800 ;
        RECT 12.470 -0.300 12.770 1.040 ;
        RECT 0.000 -0.300 13.530 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 4.895 1.545 5.325 1.965 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 2.960 0.835 3.990 ;
        RECT 2.535 2.970 2.835 3.990 ;
        RECT 3.325 2.970 3.625 3.990 ;
        RECT 5.335 2.915 5.635 3.990 ;
        RECT 6.300 2.905 6.600 3.990 ;
        RECT 8.050 2.900 8.350 3.990 ;
        RECT 9.120 2.900 9.420 3.990 ;
        RECT 10.990 2.870 11.290 3.990 ;
        RECT 12.470 2.860 12.770 3.990 ;
        RECT 0.000 3.390 13.530 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.010 0.340 2.300 ;
        RECT 0.170 1.585 1.340 1.755 ;
        RECT 1.170 0.605 1.340 2.650 ;
        RECT 1.170 0.605 1.525 0.775 ;
        RECT 1.170 2.480 1.895 2.650 ;
        RECT 1.595 2.480 1.895 2.745 ;
        RECT 2.900 1.125 3.680 1.295 ;
        RECT 3.510 1.125 3.680 2.350 ;
        RECT 2.980 2.050 3.680 2.350 ;
        RECT 3.510 1.585 3.835 1.755 ;
        RECT 1.520 1.010 1.700 2.300 ;
        RECT 1.520 1.010 1.730 1.310 ;
        RECT 1.520 2.120 2.330 2.300 ;
        RECT 2.160 2.120 2.330 2.780 ;
        RECT 2.160 2.610 4.030 2.780 ;
        RECT 3.850 2.610 4.030 3.080 ;
        RECT 3.850 2.910 4.365 3.080 ;
        RECT 4.850 1.125 5.685 1.295 ;
        RECT 5.505 1.125 5.685 2.335 ;
        RECT 4.780 2.165 5.685 2.335 ;
        RECT 5.505 1.695 5.790 1.995 ;
        RECT 3.860 1.125 4.480 1.295 ;
        RECT 4.310 1.125 4.480 2.725 ;
        RECT 6.550 1.660 6.720 2.725 ;
        RECT 4.310 2.555 6.720 2.725 ;
        RECT 7.285 1.200 7.455 2.445 ;
        RECT 7.250 1.200 7.550 1.370 ;
        RECT 7.285 1.930 8.315 2.100 ;
        RECT 8.525 1.685 8.655 1.985 ;
        RECT 8.420 1.685 8.430 2.079 ;
        RECT 8.430 1.685 8.440 2.069 ;
        RECT 8.440 1.685 8.450 2.059 ;
        RECT 8.450 1.685 8.460 2.049 ;
        RECT 8.460 1.685 8.470 2.039 ;
        RECT 8.470 1.685 8.480 2.029 ;
        RECT 8.480 1.685 8.490 2.019 ;
        RECT 8.490 1.685 8.500 2.009 ;
        RECT 8.500 1.685 8.510 1.999 ;
        RECT 8.510 1.685 8.520 1.989 ;
        RECT 8.520 1.685 8.526 1.985 ;
        RECT 8.410 1.835 8.420 2.089 ;
        RECT 8.315 1.930 8.325 2.100 ;
        RECT 8.325 1.920 8.335 2.100 ;
        RECT 8.335 1.910 8.345 2.100 ;
        RECT 8.345 1.900 8.355 2.100 ;
        RECT 8.355 1.890 8.365 2.100 ;
        RECT 8.365 1.880 8.375 2.100 ;
        RECT 8.375 1.870 8.385 2.100 ;
        RECT 8.385 1.860 8.395 2.100 ;
        RECT 8.395 1.850 8.405 2.100 ;
        RECT 8.405 1.840 8.411 2.100 ;
        RECT 2.990 0.490 3.290 0.945 ;
        RECT 2.990 0.775 6.635 0.945 ;
        RECT 7.015 0.480 7.760 0.650 ;
        RECT 8.705 0.490 9.005 0.935 ;
        RECT 8.130 0.765 9.005 0.935 ;
        RECT 8.045 0.690 8.055 0.934 ;
        RECT 8.055 0.700 8.065 0.934 ;
        RECT 8.065 0.710 8.075 0.934 ;
        RECT 8.075 0.720 8.085 0.934 ;
        RECT 8.085 0.730 8.095 0.934 ;
        RECT 8.095 0.740 8.105 0.934 ;
        RECT 8.105 0.750 8.115 0.934 ;
        RECT 8.115 0.760 8.125 0.934 ;
        RECT 8.125 0.765 8.131 0.935 ;
        RECT 7.845 0.490 7.855 0.734 ;
        RECT 7.855 0.500 7.865 0.744 ;
        RECT 7.865 0.510 7.875 0.754 ;
        RECT 7.875 0.520 7.885 0.764 ;
        RECT 7.885 0.530 7.895 0.774 ;
        RECT 7.895 0.540 7.905 0.784 ;
        RECT 7.905 0.550 7.915 0.794 ;
        RECT 7.915 0.560 7.925 0.804 ;
        RECT 7.925 0.570 7.935 0.814 ;
        RECT 7.935 0.580 7.945 0.824 ;
        RECT 7.945 0.590 7.955 0.834 ;
        RECT 7.955 0.600 7.965 0.844 ;
        RECT 7.965 0.610 7.975 0.854 ;
        RECT 7.975 0.620 7.985 0.864 ;
        RECT 7.985 0.630 7.995 0.874 ;
        RECT 7.995 0.640 8.005 0.884 ;
        RECT 8.005 0.650 8.015 0.894 ;
        RECT 8.015 0.660 8.025 0.904 ;
        RECT 8.025 0.670 8.035 0.914 ;
        RECT 8.035 0.680 8.045 0.924 ;
        RECT 7.760 0.480 7.770 0.650 ;
        RECT 7.770 0.480 7.780 0.660 ;
        RECT 7.780 0.480 7.790 0.670 ;
        RECT 7.790 0.480 7.800 0.680 ;
        RECT 7.800 0.480 7.810 0.690 ;
        RECT 7.810 0.480 7.820 0.700 ;
        RECT 7.820 0.480 7.830 0.710 ;
        RECT 7.830 0.480 7.840 0.720 ;
        RECT 7.840 0.480 7.846 0.730 ;
        RECT 6.930 0.480 6.940 0.724 ;
        RECT 6.940 0.480 6.950 0.714 ;
        RECT 6.950 0.480 6.960 0.704 ;
        RECT 6.960 0.480 6.970 0.694 ;
        RECT 6.970 0.480 6.980 0.684 ;
        RECT 6.980 0.480 6.990 0.674 ;
        RECT 6.990 0.480 7.000 0.664 ;
        RECT 7.000 0.480 7.010 0.654 ;
        RECT 7.010 0.480 7.016 0.650 ;
        RECT 6.720 0.690 6.730 0.934 ;
        RECT 6.730 0.680 6.740 0.924 ;
        RECT 6.740 0.670 6.750 0.914 ;
        RECT 6.750 0.660 6.760 0.904 ;
        RECT 6.760 0.650 6.770 0.894 ;
        RECT 6.770 0.640 6.780 0.884 ;
        RECT 6.780 0.630 6.790 0.874 ;
        RECT 6.790 0.620 6.800 0.864 ;
        RECT 6.800 0.610 6.810 0.854 ;
        RECT 6.810 0.600 6.820 0.844 ;
        RECT 6.820 0.590 6.830 0.834 ;
        RECT 6.830 0.580 6.840 0.824 ;
        RECT 6.840 0.570 6.850 0.814 ;
        RECT 6.850 0.560 6.860 0.804 ;
        RECT 6.860 0.550 6.870 0.794 ;
        RECT 6.870 0.540 6.880 0.784 ;
        RECT 6.880 0.530 6.890 0.774 ;
        RECT 6.890 0.520 6.900 0.764 ;
        RECT 6.900 0.510 6.910 0.754 ;
        RECT 6.910 0.500 6.920 0.744 ;
        RECT 6.920 0.490 6.930 0.734 ;
        RECT 6.635 0.775 6.645 0.945 ;
        RECT 6.645 0.765 6.655 0.945 ;
        RECT 6.655 0.755 6.665 0.945 ;
        RECT 6.665 0.745 6.675 0.945 ;
        RECT 6.675 0.735 6.685 0.945 ;
        RECT 6.685 0.725 6.695 0.945 ;
        RECT 6.695 0.715 6.705 0.945 ;
        RECT 6.705 0.705 6.715 0.945 ;
        RECT 6.715 0.695 6.721 0.945 ;
        RECT 8.060 1.125 8.240 1.750 ;
        RECT 7.940 1.580 8.240 1.750 ;
        RECT 8.060 1.125 9.155 1.295 ;
        RECT 8.985 1.125 9.155 2.340 ;
        RECT 8.600 2.170 9.155 2.340 ;
        RECT 8.985 1.570 9.550 1.740 ;
        RECT 5.970 1.125 6.140 2.365 ;
        RECT 5.910 1.125 6.900 1.295 ;
        RECT 7.075 2.625 7.245 2.955 ;
        RECT 7.185 0.830 7.680 1.000 ;
        RECT 7.635 2.530 7.805 2.795 ;
        RECT 7.070 2.625 7.805 2.795 ;
        RECT 9.755 0.580 9.925 2.700 ;
        RECT 7.635 2.530 9.925 2.700 ;
        RECT 9.755 0.580 10.065 0.880 ;
        RECT 9.760 2.575 10.485 2.745 ;
        RECT 10.315 2.575 10.485 2.885 ;
        RECT 7.100 0.830 7.110 1.074 ;
        RECT 7.110 0.830 7.120 1.064 ;
        RECT 7.120 0.830 7.130 1.054 ;
        RECT 7.130 0.830 7.140 1.044 ;
        RECT 7.140 0.830 7.150 1.034 ;
        RECT 7.150 0.830 7.160 1.024 ;
        RECT 7.160 0.830 7.170 1.014 ;
        RECT 7.170 0.830 7.180 1.004 ;
        RECT 7.180 0.830 7.186 1.000 ;
        RECT 7.070 0.860 7.080 1.104 ;
        RECT 7.080 0.850 7.090 1.094 ;
        RECT 7.090 0.840 7.100 1.084 ;
        RECT 6.900 1.030 6.910 2.794 ;
        RECT 6.910 1.020 6.920 2.794 ;
        RECT 6.920 1.010 6.930 2.794 ;
        RECT 6.930 1.000 6.940 2.794 ;
        RECT 6.940 0.990 6.950 2.794 ;
        RECT 6.950 0.980 6.960 2.794 ;
        RECT 6.960 0.970 6.970 2.794 ;
        RECT 6.970 0.960 6.980 2.794 ;
        RECT 6.980 0.950 6.990 2.794 ;
        RECT 6.990 0.940 7.000 2.794 ;
        RECT 7.000 0.930 7.010 2.794 ;
        RECT 7.010 0.920 7.020 2.794 ;
        RECT 7.020 0.910 7.030 2.794 ;
        RECT 7.030 0.900 7.040 2.794 ;
        RECT 7.040 0.890 7.050 2.794 ;
        RECT 7.050 0.880 7.060 2.794 ;
        RECT 7.060 0.870 7.070 2.794 ;
        RECT 11.420 1.125 11.760 1.295 ;
        RECT 11.590 0.500 11.760 2.330 ;
        RECT 11.420 2.160 11.760 2.330 ;
        RECT 11.590 0.500 11.795 0.800 ;
        RECT 11.590 1.665 12.090 1.835 ;
        RECT 10.105 1.060 10.275 1.845 ;
        RECT 10.130 1.675 10.310 2.395 ;
        RECT 10.860 1.675 11.030 2.680 ;
        RECT 10.105 1.675 11.410 1.845 ;
        RECT 12.705 1.535 12.875 2.680 ;
        RECT 10.860 2.510 12.875 2.680 ;
  END 
END FFEDCRHDMXHT

MACRO FFEDCRHDLXHT
  CLASS  CORE ;
  FOREIGN FFEDCRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.530 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.145 1.060 13.430 2.280 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 12.050 0.850 12.260 1.445 ;
        RECT 12.050 1.265 12.615 1.445 ;
        RECT 12.435 1.265 12.615 2.215 ;
        RECT 12.020 2.045 12.615 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.115 1.265 2.440 1.795 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.225 2.560 0.870 2.770 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.620 1.625 2.800 2.430 ;
        RECT 2.510 2.085 2.800 2.430 ;
        RECT 2.620 1.625 2.980 1.795 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.685 ;
        RECT 2.350 -0.300 2.650 0.815 ;
        RECT 3.525 -0.300 4.545 0.555 ;
        RECT 5.530 -0.300 6.510 0.555 ;
        RECT 8.235 -0.300 8.535 0.575 ;
        RECT 9.205 -0.300 9.375 0.930 ;
        RECT 11.050 -0.300 11.350 0.825 ;
        RECT 12.570 -0.300 12.870 0.745 ;
        RECT 0.000 -0.300 13.530 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 4.895 1.545 5.325 1.965 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.960 0.955 3.990 ;
        RECT 2.425 2.970 2.725 3.990 ;
        RECT 3.325 2.970 3.625 3.990 ;
        RECT 5.325 2.915 5.625 3.990 ;
        RECT 6.300 2.905 6.600 3.990 ;
        RECT 8.080 2.900 8.380 3.990 ;
        RECT 9.140 2.900 9.440 3.990 ;
        RECT 11.080 2.870 11.380 3.990 ;
        RECT 12.560 2.860 12.860 3.990 ;
        RECT 0.000 3.390 13.530 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.010 0.340 2.300 ;
        RECT 0.170 1.585 1.340 1.755 ;
        RECT 1.170 0.660 1.340 2.650 ;
        RECT 1.170 0.660 1.525 0.830 ;
        RECT 1.170 2.480 1.940 2.650 ;
        RECT 1.770 2.480 1.940 2.810 ;
        RECT 2.980 2.000 3.150 2.300 ;
        RECT 2.900 1.125 3.455 1.295 ;
        RECT 3.285 1.125 3.455 2.170 ;
        RECT 2.980 2.000 3.455 2.170 ;
        RECT 3.285 1.575 3.835 1.745 ;
        RECT 1.565 1.010 1.735 2.300 ;
        RECT 1.565 2.120 2.330 2.300 ;
        RECT 2.160 2.120 2.330 2.780 ;
        RECT 2.160 2.610 4.030 2.780 ;
        RECT 3.850 2.610 4.030 3.075 ;
        RECT 3.850 2.905 4.365 3.075 ;
        RECT 4.860 1.125 5.685 1.295 ;
        RECT 5.505 1.125 5.685 2.335 ;
        RECT 4.780 2.165 5.685 2.335 ;
        RECT 5.505 1.600 5.790 1.900 ;
        RECT 3.860 1.125 4.480 1.295 ;
        RECT 4.310 1.125 4.480 2.725 ;
        RECT 6.550 1.660 6.720 2.725 ;
        RECT 4.310 2.555 6.720 2.725 ;
        RECT 7.285 1.200 7.455 2.495 ;
        RECT 7.250 1.200 7.550 1.370 ;
        RECT 7.285 1.930 8.340 2.100 ;
        RECT 8.545 1.685 8.660 1.985 ;
        RECT 8.450 1.685 8.460 2.069 ;
        RECT 8.460 1.685 8.470 2.059 ;
        RECT 8.470 1.685 8.480 2.049 ;
        RECT 8.480 1.685 8.490 2.039 ;
        RECT 8.490 1.685 8.500 2.029 ;
        RECT 8.500 1.685 8.510 2.019 ;
        RECT 8.510 1.685 8.520 2.009 ;
        RECT 8.520 1.685 8.530 1.999 ;
        RECT 8.530 1.685 8.540 1.989 ;
        RECT 8.540 1.685 8.546 1.985 ;
        RECT 8.430 1.840 8.440 2.090 ;
        RECT 8.440 1.830 8.450 2.080 ;
        RECT 8.340 1.930 8.350 2.100 ;
        RECT 8.350 1.920 8.360 2.100 ;
        RECT 8.360 1.910 8.370 2.100 ;
        RECT 8.370 1.900 8.380 2.100 ;
        RECT 8.380 1.890 8.390 2.100 ;
        RECT 8.390 1.880 8.400 2.100 ;
        RECT 8.400 1.870 8.410 2.100 ;
        RECT 8.410 1.860 8.420 2.100 ;
        RECT 8.420 1.850 8.430 2.100 ;
        RECT 2.990 0.490 3.290 0.945 ;
        RECT 2.990 0.775 6.610 0.945 ;
        RECT 6.990 0.480 7.760 0.650 ;
        RECT 8.720 0.510 9.020 0.935 ;
        RECT 8.130 0.765 9.020 0.935 ;
        RECT 8.045 0.690 8.055 0.934 ;
        RECT 8.055 0.700 8.065 0.934 ;
        RECT 8.065 0.710 8.075 0.934 ;
        RECT 8.075 0.720 8.085 0.934 ;
        RECT 8.085 0.730 8.095 0.934 ;
        RECT 8.095 0.740 8.105 0.934 ;
        RECT 8.105 0.750 8.115 0.934 ;
        RECT 8.115 0.760 8.125 0.934 ;
        RECT 8.125 0.765 8.131 0.935 ;
        RECT 7.845 0.490 7.855 0.734 ;
        RECT 7.855 0.500 7.865 0.744 ;
        RECT 7.865 0.510 7.875 0.754 ;
        RECT 7.875 0.520 7.885 0.764 ;
        RECT 7.885 0.530 7.895 0.774 ;
        RECT 7.895 0.540 7.905 0.784 ;
        RECT 7.905 0.550 7.915 0.794 ;
        RECT 7.915 0.560 7.925 0.804 ;
        RECT 7.925 0.570 7.935 0.814 ;
        RECT 7.935 0.580 7.945 0.824 ;
        RECT 7.945 0.590 7.955 0.834 ;
        RECT 7.955 0.600 7.965 0.844 ;
        RECT 7.965 0.610 7.975 0.854 ;
        RECT 7.975 0.620 7.985 0.864 ;
        RECT 7.985 0.630 7.995 0.874 ;
        RECT 7.995 0.640 8.005 0.884 ;
        RECT 8.005 0.650 8.015 0.894 ;
        RECT 8.015 0.660 8.025 0.904 ;
        RECT 8.025 0.670 8.035 0.914 ;
        RECT 8.035 0.680 8.045 0.924 ;
        RECT 7.760 0.480 7.770 0.650 ;
        RECT 7.770 0.480 7.780 0.660 ;
        RECT 7.780 0.480 7.790 0.670 ;
        RECT 7.790 0.480 7.800 0.680 ;
        RECT 7.800 0.480 7.810 0.690 ;
        RECT 7.810 0.480 7.820 0.700 ;
        RECT 7.820 0.480 7.830 0.710 ;
        RECT 7.830 0.480 7.840 0.720 ;
        RECT 7.840 0.480 7.846 0.730 ;
        RECT 6.905 0.480 6.915 0.724 ;
        RECT 6.915 0.480 6.925 0.714 ;
        RECT 6.925 0.480 6.935 0.704 ;
        RECT 6.935 0.480 6.945 0.694 ;
        RECT 6.945 0.480 6.955 0.684 ;
        RECT 6.955 0.480 6.965 0.674 ;
        RECT 6.965 0.480 6.975 0.664 ;
        RECT 6.975 0.480 6.985 0.654 ;
        RECT 6.985 0.480 6.991 0.650 ;
        RECT 6.695 0.690 6.705 0.934 ;
        RECT 6.705 0.680 6.715 0.924 ;
        RECT 6.715 0.670 6.725 0.914 ;
        RECT 6.725 0.660 6.735 0.904 ;
        RECT 6.735 0.650 6.745 0.894 ;
        RECT 6.745 0.640 6.755 0.884 ;
        RECT 6.755 0.630 6.765 0.874 ;
        RECT 6.765 0.620 6.775 0.864 ;
        RECT 6.775 0.610 6.785 0.854 ;
        RECT 6.785 0.600 6.795 0.844 ;
        RECT 6.795 0.590 6.805 0.834 ;
        RECT 6.805 0.580 6.815 0.824 ;
        RECT 6.815 0.570 6.825 0.814 ;
        RECT 6.825 0.560 6.835 0.804 ;
        RECT 6.835 0.550 6.845 0.794 ;
        RECT 6.845 0.540 6.855 0.784 ;
        RECT 6.855 0.530 6.865 0.774 ;
        RECT 6.865 0.520 6.875 0.764 ;
        RECT 6.875 0.510 6.885 0.754 ;
        RECT 6.885 0.500 6.895 0.744 ;
        RECT 6.895 0.490 6.905 0.734 ;
        RECT 6.610 0.775 6.620 0.945 ;
        RECT 6.620 0.765 6.630 0.945 ;
        RECT 6.630 0.755 6.640 0.945 ;
        RECT 6.640 0.745 6.650 0.945 ;
        RECT 6.650 0.735 6.660 0.945 ;
        RECT 6.660 0.725 6.670 0.945 ;
        RECT 6.670 0.715 6.680 0.945 ;
        RECT 6.680 0.705 6.690 0.945 ;
        RECT 6.690 0.695 6.696 0.945 ;
        RECT 8.080 1.125 8.250 1.700 ;
        RECT 7.945 1.530 8.250 1.700 ;
        RECT 8.080 1.125 9.010 1.295 ;
        RECT 8.840 1.125 9.010 2.340 ;
        RECT 8.630 2.170 9.010 2.340 ;
        RECT 8.840 1.570 9.600 1.740 ;
        RECT 5.970 1.125 6.140 2.365 ;
        RECT 5.910 1.125 6.900 1.295 ;
        RECT 7.185 0.830 7.680 1.000 ;
        RECT 7.690 2.530 7.860 2.905 ;
        RECT 7.070 2.735 7.860 2.905 ;
        RECT 9.785 0.710 9.955 2.780 ;
        RECT 7.690 2.530 9.955 2.700 ;
        RECT 9.785 0.710 10.160 0.880 ;
        RECT 9.785 2.610 10.640 2.780 ;
        RECT 7.100 0.830 7.110 1.074 ;
        RECT 7.110 0.830 7.120 1.064 ;
        RECT 7.120 0.830 7.130 1.054 ;
        RECT 7.130 0.830 7.140 1.044 ;
        RECT 7.140 0.830 7.150 1.034 ;
        RECT 7.150 0.830 7.160 1.024 ;
        RECT 7.160 0.830 7.170 1.014 ;
        RECT 7.170 0.830 7.180 1.004 ;
        RECT 7.180 0.830 7.186 1.000 ;
        RECT 7.070 0.860 7.080 1.104 ;
        RECT 7.080 0.850 7.090 1.094 ;
        RECT 7.090 0.840 7.100 1.084 ;
        RECT 6.900 1.030 6.910 2.904 ;
        RECT 6.910 1.020 6.920 2.904 ;
        RECT 6.920 1.010 6.930 2.904 ;
        RECT 6.930 1.000 6.940 2.904 ;
        RECT 6.940 0.990 6.950 2.904 ;
        RECT 6.950 0.980 6.960 2.904 ;
        RECT 6.960 0.970 6.970 2.904 ;
        RECT 6.970 0.960 6.980 2.904 ;
        RECT 6.980 0.950 6.990 2.904 ;
        RECT 6.990 0.940 7.000 2.904 ;
        RECT 7.000 0.930 7.010 2.904 ;
        RECT 7.010 0.920 7.020 2.904 ;
        RECT 7.020 0.910 7.030 2.904 ;
        RECT 7.030 0.900 7.040 2.904 ;
        RECT 7.040 0.890 7.050 2.904 ;
        RECT 7.050 0.880 7.060 2.904 ;
        RECT 7.060 0.870 7.070 2.904 ;
        RECT 11.510 1.125 11.810 1.295 ;
        RECT 11.640 0.500 11.810 2.330 ;
        RECT 11.510 2.160 11.810 2.330 ;
        RECT 11.640 0.500 11.950 0.670 ;
        RECT 11.640 1.665 12.255 1.835 ;
        RECT 10.135 1.060 10.345 1.360 ;
        RECT 10.165 1.060 10.345 2.420 ;
        RECT 10.165 1.675 11.425 1.845 ;
        RECT 11.160 1.675 11.330 2.680 ;
        RECT 11.255 1.610 11.425 1.910 ;
        RECT 11.160 1.675 11.425 1.910 ;
        RECT 12.795 1.610 12.965 2.680 ;
        RECT 11.160 2.510 12.965 2.680 ;
  END 
END FFEDCRHDLXHT

MACRO FFEDCRHD1XHT
  CLASS  CORE ;
  FOREIGN FFEDCRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.530 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.055 0.720 13.225 2.960 ;
        RECT 13.055 1.645 13.430 2.040 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.985 1.300 12.470 1.480 ;
        RECT 11.985 0.720 12.270 1.480 ;
        RECT 12.270 1.300 12.470 2.215 ;
        RECT 11.950 2.045 12.470 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.115 1.265 2.440 1.795 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.225 2.560 0.830 2.770 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.620 1.625 2.800 2.430 ;
        RECT 2.510 2.085 2.800 2.430 ;
        RECT 2.620 1.625 2.980 1.795 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.685 ;
        RECT 2.425 -0.300 2.725 0.745 ;
        RECT 3.470 -0.300 3.770 0.595 ;
        RECT 4.385 -0.300 4.685 0.595 ;
        RECT 5.445 -0.300 5.745 0.595 ;
        RECT 6.220 -0.300 6.520 0.595 ;
        RECT 8.205 -0.300 8.505 0.575 ;
        RECT 9.185 -0.300 9.355 1.220 ;
        RECT 10.990 -0.300 11.290 0.735 ;
        RECT 12.535 -0.300 12.705 1.120 ;
        RECT 0.000 -0.300 13.530 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 4.895 1.545 5.325 1.965 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 2.960 0.835 3.990 ;
        RECT 2.425 2.970 2.725 3.990 ;
        RECT 3.325 2.970 3.625 3.990 ;
        RECT 5.335 2.915 5.635 3.990 ;
        RECT 6.300 2.905 6.600 3.990 ;
        RECT 8.050 2.900 8.350 3.990 ;
        RECT 9.120 2.900 9.420 3.990 ;
        RECT 10.990 2.870 11.290 3.990 ;
        RECT 12.470 2.975 12.770 3.990 ;
        RECT 0.000 3.390 13.530 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.010 0.340 2.300 ;
        RECT 0.170 1.585 1.340 1.755 ;
        RECT 1.170 0.605 1.340 3.040 ;
        RECT 1.170 0.605 1.525 0.775 ;
        RECT 1.170 2.870 1.940 3.040 ;
        RECT 1.770 2.870 1.940 3.170 ;
        RECT 2.980 2.000 3.150 2.300 ;
        RECT 2.900 1.125 3.475 1.295 ;
        RECT 3.305 1.125 3.475 2.170 ;
        RECT 2.980 2.000 3.475 2.170 ;
        RECT 3.305 1.575 3.835 1.745 ;
        RECT 1.520 1.010 1.690 2.640 ;
        RECT 2.160 2.460 2.330 2.780 ;
        RECT 1.520 2.460 2.330 2.640 ;
        RECT 2.160 2.610 4.020 2.780 ;
        RECT 3.850 2.610 4.020 3.075 ;
        RECT 3.850 2.905 4.365 3.075 ;
        RECT 4.895 1.125 5.675 1.295 ;
        RECT 5.505 1.125 5.675 2.335 ;
        RECT 4.780 2.165 5.675 2.335 ;
        RECT 5.505 1.530 5.790 1.830 ;
        RECT 4.310 1.980 4.545 2.280 ;
        RECT 3.860 1.125 4.490 1.295 ;
        RECT 4.310 1.125 4.490 2.280 ;
        RECT 4.375 1.980 4.545 2.725 ;
        RECT 6.550 1.660 6.720 2.725 ;
        RECT 4.375 2.555 6.720 2.725 ;
        RECT 7.285 1.200 7.455 2.445 ;
        RECT 7.250 1.200 7.550 1.370 ;
        RECT 7.285 1.930 8.310 2.100 ;
        RECT 8.515 1.685 8.655 1.985 ;
        RECT 8.485 1.685 8.495 2.005 ;
        RECT 8.495 1.685 8.505 1.995 ;
        RECT 8.505 1.685 8.515 1.985 ;
        RECT 8.400 1.840 8.410 2.090 ;
        RECT 8.410 1.830 8.420 2.080 ;
        RECT 8.420 1.820 8.430 2.070 ;
        RECT 8.430 1.810 8.440 2.060 ;
        RECT 8.440 1.800 8.450 2.050 ;
        RECT 8.450 1.790 8.460 2.040 ;
        RECT 8.460 1.780 8.470 2.030 ;
        RECT 8.470 1.770 8.480 2.020 ;
        RECT 8.480 1.760 8.486 2.014 ;
        RECT 8.310 1.930 8.320 2.100 ;
        RECT 8.320 1.920 8.330 2.100 ;
        RECT 8.330 1.910 8.340 2.100 ;
        RECT 8.340 1.900 8.350 2.100 ;
        RECT 8.350 1.890 8.360 2.100 ;
        RECT 8.360 1.880 8.370 2.100 ;
        RECT 8.370 1.870 8.380 2.100 ;
        RECT 8.380 1.860 8.390 2.100 ;
        RECT 8.390 1.850 8.400 2.100 ;
        RECT 2.990 0.490 3.290 0.945 ;
        RECT 2.990 0.775 6.635 0.945 ;
        RECT 7.015 0.480 7.760 0.650 ;
        RECT 8.705 0.490 9.005 0.935 ;
        RECT 8.130 0.765 9.005 0.935 ;
        RECT 8.045 0.690 8.055 0.934 ;
        RECT 8.055 0.700 8.065 0.934 ;
        RECT 8.065 0.710 8.075 0.934 ;
        RECT 8.075 0.720 8.085 0.934 ;
        RECT 8.085 0.730 8.095 0.934 ;
        RECT 8.095 0.740 8.105 0.934 ;
        RECT 8.105 0.750 8.115 0.934 ;
        RECT 8.115 0.760 8.125 0.934 ;
        RECT 8.125 0.765 8.131 0.935 ;
        RECT 7.845 0.490 7.855 0.734 ;
        RECT 7.855 0.500 7.865 0.744 ;
        RECT 7.865 0.510 7.875 0.754 ;
        RECT 7.875 0.520 7.885 0.764 ;
        RECT 7.885 0.530 7.895 0.774 ;
        RECT 7.895 0.540 7.905 0.784 ;
        RECT 7.905 0.550 7.915 0.794 ;
        RECT 7.915 0.560 7.925 0.804 ;
        RECT 7.925 0.570 7.935 0.814 ;
        RECT 7.935 0.580 7.945 0.824 ;
        RECT 7.945 0.590 7.955 0.834 ;
        RECT 7.955 0.600 7.965 0.844 ;
        RECT 7.965 0.610 7.975 0.854 ;
        RECT 7.975 0.620 7.985 0.864 ;
        RECT 7.985 0.630 7.995 0.874 ;
        RECT 7.995 0.640 8.005 0.884 ;
        RECT 8.005 0.650 8.015 0.894 ;
        RECT 8.015 0.660 8.025 0.904 ;
        RECT 8.025 0.670 8.035 0.914 ;
        RECT 8.035 0.680 8.045 0.924 ;
        RECT 7.760 0.480 7.770 0.650 ;
        RECT 7.770 0.480 7.780 0.660 ;
        RECT 7.780 0.480 7.790 0.670 ;
        RECT 7.790 0.480 7.800 0.680 ;
        RECT 7.800 0.480 7.810 0.690 ;
        RECT 7.810 0.480 7.820 0.700 ;
        RECT 7.820 0.480 7.830 0.710 ;
        RECT 7.830 0.480 7.840 0.720 ;
        RECT 7.840 0.480 7.846 0.730 ;
        RECT 6.930 0.480 6.940 0.724 ;
        RECT 6.940 0.480 6.950 0.714 ;
        RECT 6.950 0.480 6.960 0.704 ;
        RECT 6.960 0.480 6.970 0.694 ;
        RECT 6.970 0.480 6.980 0.684 ;
        RECT 6.980 0.480 6.990 0.674 ;
        RECT 6.990 0.480 7.000 0.664 ;
        RECT 7.000 0.480 7.010 0.654 ;
        RECT 7.010 0.480 7.016 0.650 ;
        RECT 6.720 0.690 6.730 0.934 ;
        RECT 6.730 0.680 6.740 0.924 ;
        RECT 6.740 0.670 6.750 0.914 ;
        RECT 6.750 0.660 6.760 0.904 ;
        RECT 6.760 0.650 6.770 0.894 ;
        RECT 6.770 0.640 6.780 0.884 ;
        RECT 6.780 0.630 6.790 0.874 ;
        RECT 6.790 0.620 6.800 0.864 ;
        RECT 6.800 0.610 6.810 0.854 ;
        RECT 6.810 0.600 6.820 0.844 ;
        RECT 6.820 0.590 6.830 0.834 ;
        RECT 6.830 0.580 6.840 0.824 ;
        RECT 6.840 0.570 6.850 0.814 ;
        RECT 6.850 0.560 6.860 0.804 ;
        RECT 6.860 0.550 6.870 0.794 ;
        RECT 6.870 0.540 6.880 0.784 ;
        RECT 6.880 0.530 6.890 0.774 ;
        RECT 6.890 0.520 6.900 0.764 ;
        RECT 6.900 0.510 6.910 0.754 ;
        RECT 6.910 0.500 6.920 0.744 ;
        RECT 6.920 0.490 6.930 0.734 ;
        RECT 6.635 0.775 6.645 0.945 ;
        RECT 6.645 0.765 6.655 0.945 ;
        RECT 6.655 0.755 6.665 0.945 ;
        RECT 6.665 0.745 6.675 0.945 ;
        RECT 6.675 0.735 6.685 0.945 ;
        RECT 6.685 0.725 6.695 0.945 ;
        RECT 6.695 0.715 6.705 0.945 ;
        RECT 6.705 0.705 6.715 0.945 ;
        RECT 6.715 0.695 6.721 0.945 ;
        RECT 8.060 1.125 8.230 1.750 ;
        RECT 7.930 1.580 8.230 1.750 ;
        RECT 8.060 1.125 9.005 1.295 ;
        RECT 8.835 1.125 9.005 2.340 ;
        RECT 8.600 2.170 9.005 2.340 ;
        RECT 8.835 1.570 9.550 1.740 ;
        RECT 5.970 1.125 6.140 2.365 ;
        RECT 5.910 1.125 6.900 1.295 ;
        RECT 7.105 2.645 7.275 3.115 ;
        RECT 7.185 0.830 7.680 1.000 ;
        RECT 7.635 2.530 7.805 2.815 ;
        RECT 7.070 2.645 7.805 2.815 ;
        RECT 7.635 2.530 9.930 2.700 ;
        RECT 9.760 0.615 9.930 2.955 ;
        RECT 9.760 0.615 10.130 0.785 ;
        RECT 9.760 2.785 10.550 2.955 ;
        RECT 10.250 2.785 10.550 3.020 ;
        RECT 7.100 0.830 7.110 1.074 ;
        RECT 7.110 0.830 7.120 1.064 ;
        RECT 7.120 0.830 7.130 1.054 ;
        RECT 7.130 0.830 7.140 1.044 ;
        RECT 7.140 0.830 7.150 1.034 ;
        RECT 7.150 0.830 7.160 1.024 ;
        RECT 7.160 0.830 7.170 1.014 ;
        RECT 7.170 0.830 7.180 1.004 ;
        RECT 7.180 0.830 7.186 1.000 ;
        RECT 7.070 0.860 7.080 1.104 ;
        RECT 7.080 0.850 7.090 1.094 ;
        RECT 7.090 0.840 7.100 1.084 ;
        RECT 6.900 1.030 6.910 2.814 ;
        RECT 6.910 1.020 6.920 2.814 ;
        RECT 6.920 1.010 6.930 2.814 ;
        RECT 6.930 1.000 6.940 2.814 ;
        RECT 6.940 0.990 6.950 2.814 ;
        RECT 6.950 0.980 6.960 2.814 ;
        RECT 6.960 0.970 6.970 2.814 ;
        RECT 6.970 0.960 6.980 2.814 ;
        RECT 6.980 0.950 6.990 2.814 ;
        RECT 6.990 0.940 7.000 2.814 ;
        RECT 7.000 0.930 7.010 2.814 ;
        RECT 7.010 0.920 7.020 2.814 ;
        RECT 7.020 0.910 7.030 2.814 ;
        RECT 7.030 0.900 7.040 2.814 ;
        RECT 7.040 0.890 7.050 2.814 ;
        RECT 7.050 0.880 7.060 2.814 ;
        RECT 7.060 0.870 7.070 2.814 ;
        RECT 11.420 1.125 11.760 1.295 ;
        RECT 11.590 0.500 11.760 2.330 ;
        RECT 11.420 2.160 11.760 2.330 ;
        RECT 11.590 0.500 11.795 0.800 ;
        RECT 11.590 1.665 12.090 1.835 ;
        RECT 10.130 1.060 10.310 2.395 ;
        RECT 10.860 1.675 11.030 2.680 ;
        RECT 10.130 1.675 11.410 1.845 ;
        RECT 12.705 1.520 12.875 2.680 ;
        RECT 10.860 2.510 12.875 2.680 ;
  END 
END FFEDCRHD1XHT

MACRO FFDSRHQHDMXHT
  CLASS  CORE ;
  FOREIGN FFDSRHQHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.480 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.760 1.980 11.300 2.430 ;
        RECT 10.970 1.060 11.300 1.360 ;
        RECT 11.090 1.060 11.300 2.620 ;
        RECT 11.065 1.980 11.300 2.620 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.600 2.560 2.050 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 9.940 1.260 10.215 1.735 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.995 ;
        RECT 2.175 -0.300 2.475 1.230 ;
        RECT 4.035 -0.300 4.335 1.065 ;
        RECT 6.160 -0.300 6.460 0.715 ;
        RECT 8.050 -0.300 8.350 0.795 ;
        RECT 10.420 -0.300 10.720 1.285 ;
        RECT 0.000 -0.300 11.480 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.870 1.260 1.130 1.730 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 8.230 1.330 8.825 1.540 ;
        RECT 8.425 1.330 8.825 1.815 ;
        RECT 6.545 2.625 6.611 2.805 ;
        RECT 6.555 2.625 6.611 2.815 ;
        RECT 6.565 2.625 6.611 2.825 ;
        RECT 6.575 2.625 6.611 2.835 ;
        RECT 6.640 3.020 7.800 3.189 ;
        RECT 5.810 2.625 5.980 2.925 ;
        RECT 6.585 2.625 6.611 2.845 ;
        RECT 6.585 2.835 6.820 2.845 ;
        RECT 6.595 2.625 6.611 2.855 ;
        RECT 6.595 2.835 6.820 2.855 ;
        RECT 6.605 2.625 6.611 2.865 ;
        RECT 6.605 2.835 6.820 2.865 ;
        RECT 6.610 2.625 6.611 2.869 ;
        RECT 5.810 2.625 6.611 2.795 ;
        RECT 6.610 2.635 6.620 2.869 ;
        RECT 6.610 2.835 6.820 2.869 ;
        RECT 5.810 2.635 6.620 2.795 ;
        RECT 6.620 2.645 6.630 2.879 ;
        RECT 6.620 2.835 6.820 2.879 ;
        RECT 5.810 2.645 6.630 2.795 ;
        RECT 6.630 2.655 6.640 2.889 ;
        RECT 6.630 2.835 6.820 2.889 ;
        RECT 5.810 2.655 6.640 2.795 ;
        RECT 6.640 2.665 6.650 3.189 ;
        RECT 5.810 2.665 6.650 2.795 ;
        RECT 6.640 2.675 6.660 3.189 ;
        RECT 5.810 2.675 6.660 2.795 ;
        RECT 6.640 2.685 6.670 3.189 ;
        RECT 5.810 2.685 6.670 2.795 ;
        RECT 6.640 2.695 6.680 3.189 ;
        RECT 5.810 2.695 6.680 2.795 ;
        RECT 6.640 2.705 6.690 3.189 ;
        RECT 5.810 2.705 6.690 2.795 ;
        RECT 6.640 2.715 6.700 3.189 ;
        RECT 5.810 2.715 6.700 2.795 ;
        RECT 6.640 2.725 6.710 3.189 ;
        RECT 5.810 2.725 6.710 2.795 ;
        RECT 6.640 2.735 6.720 3.189 ;
        RECT 5.810 2.735 6.720 2.795 ;
        RECT 6.640 2.745 6.730 3.189 ;
        RECT 5.810 2.745 6.730 2.795 ;
        RECT 6.640 2.755 6.740 3.189 ;
        RECT 5.810 2.755 6.740 2.795 ;
        RECT 6.640 2.765 6.750 3.189 ;
        RECT 5.810 2.765 6.750 2.795 ;
        RECT 6.640 2.775 6.760 3.189 ;
        RECT 5.810 2.775 6.760 2.795 ;
        RECT 6.640 2.785 6.770 3.189 ;
        RECT 5.810 2.785 6.770 2.795 ;
        RECT 6.640 2.795 6.780 3.189 ;
        RECT 6.545 2.795 6.780 2.805 ;
        RECT 6.640 2.805 6.790 3.189 ;
        RECT 6.555 2.805 6.790 2.815 ;
        RECT 6.640 2.815 6.800 3.189 ;
        RECT 6.565 2.815 6.800 2.825 ;
        RECT 6.640 2.825 6.810 3.189 ;
        RECT 6.575 2.825 6.810 2.835 ;
        RECT 6.640 2.835 6.820 3.189 ;
        RECT 7.790 2.950 7.800 3.190 ;
        RECT 7.790 2.950 8.930 3.055 ;
        RECT 6.820 3.020 7.800 3.190 ;
        RECT 7.800 2.940 7.810 3.180 ;
        RECT 7.780 2.960 8.930 3.055 ;
        RECT 6.640 3.020 7.810 3.180 ;
        RECT 7.810 2.930 7.820 3.170 ;
        RECT 7.770 2.970 8.930 3.055 ;
        RECT 6.640 3.020 7.820 3.170 ;
        RECT 7.820 2.920 7.830 3.160 ;
        RECT 7.760 2.980 8.930 3.055 ;
        RECT 6.640 3.020 7.830 3.160 ;
        RECT 7.830 2.910 7.840 3.150 ;
        RECT 7.750 2.990 8.930 3.055 ;
        RECT 6.640 3.020 7.840 3.150 ;
        RECT 7.840 2.900 7.850 3.140 ;
        RECT 7.740 3.000 8.930 3.055 ;
        RECT 6.640 3.020 7.850 3.140 ;
        RECT 7.850 2.890 7.856 3.134 ;
        RECT 7.730 3.010 8.930 3.055 ;
        RECT 7.855 2.885 7.856 3.134 ;
        RECT 6.640 3.020 7.856 3.134 ;
        RECT 7.855 2.885 7.865 3.125 ;
        RECT 6.640 3.020 7.865 3.125 ;
        RECT 7.855 2.885 7.875 3.115 ;
        RECT 6.640 3.020 7.875 3.115 ;
        RECT 7.855 2.885 7.885 3.105 ;
        RECT 6.640 3.020 7.885 3.105 ;
        RECT 7.855 2.885 7.895 3.095 ;
        RECT 6.640 3.020 7.895 3.095 ;
        RECT 7.855 2.885 7.905 3.085 ;
        RECT 6.640 3.020 7.905 3.085 ;
        RECT 7.855 2.885 7.915 3.075 ;
        RECT 6.640 3.020 7.915 3.075 ;
        RECT 7.855 2.885 7.925 3.065 ;
        RECT 6.640 3.020 7.925 3.065 ;
        RECT 7.855 2.885 8.930 3.055 ;
        RECT 8.630 2.885 8.930 3.185 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 1.980 0.340 3.990 ;
        RECT 2.205 3.215 2.505 3.990 ;
        RECT 3.915 3.155 4.215 3.990 ;
        RECT 6.160 2.975 6.460 3.990 ;
        RECT 8.050 3.255 8.350 3.990 ;
        RECT 9.480 2.745 9.780 3.990 ;
        RECT 10.420 2.800 10.720 3.990 ;
        RECT 0.000 3.390 11.480 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.000 1.910 1.170 2.215 ;
        RECT 0.870 2.045 1.170 2.215 ;
        RECT 1.145 0.825 1.480 0.995 ;
        RECT 1.000 1.910 1.480 2.080 ;
        RECT 1.310 0.825 1.480 2.080 ;
        RECT 1.310 1.610 1.540 1.910 ;
        RECT 3.115 2.165 3.285 2.335 ;
        RECT 3.130 0.995 3.300 1.495 ;
        RECT 3.130 1.325 3.415 1.495 ;
        RECT 3.315 1.325 3.415 2.335 ;
        RECT 3.485 1.325 4.150 1.495 ;
        RECT 4.425 1.675 5.035 1.845 ;
        RECT 4.255 1.360 4.265 1.844 ;
        RECT 4.265 1.370 4.275 1.844 ;
        RECT 4.275 1.380 4.285 1.844 ;
        RECT 4.285 1.390 4.295 1.844 ;
        RECT 4.295 1.400 4.305 1.844 ;
        RECT 4.305 1.410 4.315 1.844 ;
        RECT 4.315 1.420 4.325 1.844 ;
        RECT 4.325 1.430 4.335 1.844 ;
        RECT 4.335 1.440 4.345 1.844 ;
        RECT 4.345 1.450 4.355 1.844 ;
        RECT 4.355 1.460 4.365 1.844 ;
        RECT 4.365 1.470 4.375 1.844 ;
        RECT 4.375 1.480 4.385 1.844 ;
        RECT 4.385 1.490 4.395 1.844 ;
        RECT 4.395 1.500 4.405 1.844 ;
        RECT 4.405 1.510 4.415 1.844 ;
        RECT 4.415 1.520 4.425 1.844 ;
        RECT 4.230 1.335 4.240 1.575 ;
        RECT 4.240 1.345 4.250 1.585 ;
        RECT 4.250 1.350 4.256 1.594 ;
        RECT 4.150 1.325 4.160 1.495 ;
        RECT 4.160 1.325 4.170 1.505 ;
        RECT 4.170 1.325 4.180 1.515 ;
        RECT 4.180 1.325 4.190 1.525 ;
        RECT 4.190 1.325 4.200 1.535 ;
        RECT 4.200 1.325 4.210 1.545 ;
        RECT 4.210 1.325 4.220 1.555 ;
        RECT 4.220 1.325 4.230 1.565 ;
        RECT 3.415 1.325 3.425 2.325 ;
        RECT 3.425 1.325 3.435 2.315 ;
        RECT 3.435 1.325 3.445 2.305 ;
        RECT 3.445 1.325 3.455 2.295 ;
        RECT 3.455 1.325 3.465 2.285 ;
        RECT 3.465 1.325 3.475 2.275 ;
        RECT 3.475 1.325 3.485 2.265 ;
        RECT 3.285 2.165 3.295 2.335 ;
        RECT 3.295 2.155 3.305 2.335 ;
        RECT 3.305 2.145 3.315 2.335 ;
        RECT 0.170 1.060 0.340 1.790 ;
        RECT 0.170 1.620 0.690 1.790 ;
        RECT 0.520 1.620 0.690 2.565 ;
        RECT 0.520 2.395 1.230 2.565 ;
        RECT 1.060 2.395 1.230 3.035 ;
        RECT 1.060 2.865 3.705 3.035 ;
        RECT 3.765 2.805 3.780 3.035 ;
        RECT 3.840 2.805 4.425 2.975 ;
        RECT 4.750 3.040 5.565 3.210 ;
        RECT 4.660 2.960 4.670 3.210 ;
        RECT 4.670 2.970 4.680 3.210 ;
        RECT 4.680 2.980 4.690 3.210 ;
        RECT 4.690 2.990 4.700 3.210 ;
        RECT 4.700 3.000 4.710 3.210 ;
        RECT 4.710 3.010 4.720 3.210 ;
        RECT 4.720 3.020 4.730 3.210 ;
        RECT 4.730 3.030 4.740 3.210 ;
        RECT 4.740 3.040 4.750 3.210 ;
        RECT 4.515 2.815 4.525 3.065 ;
        RECT 4.525 2.825 4.535 3.075 ;
        RECT 4.535 2.835 4.545 3.085 ;
        RECT 4.545 2.845 4.555 3.095 ;
        RECT 4.555 2.855 4.565 3.105 ;
        RECT 4.565 2.865 4.575 3.115 ;
        RECT 4.575 2.875 4.585 3.125 ;
        RECT 4.585 2.885 4.595 3.135 ;
        RECT 4.595 2.895 4.605 3.145 ;
        RECT 4.605 2.905 4.615 3.155 ;
        RECT 4.615 2.915 4.625 3.165 ;
        RECT 4.625 2.925 4.635 3.175 ;
        RECT 4.635 2.935 4.645 3.185 ;
        RECT 4.645 2.945 4.655 3.195 ;
        RECT 4.655 2.950 4.661 3.204 ;
        RECT 4.425 2.805 4.435 2.975 ;
        RECT 4.435 2.805 4.445 2.985 ;
        RECT 4.445 2.805 4.455 2.995 ;
        RECT 4.455 2.805 4.465 3.005 ;
        RECT 4.465 2.805 4.475 3.015 ;
        RECT 4.475 2.805 4.485 3.025 ;
        RECT 4.485 2.805 4.495 3.035 ;
        RECT 4.495 2.805 4.505 3.045 ;
        RECT 4.505 2.805 4.515 3.055 ;
        RECT 3.780 2.805 3.790 3.025 ;
        RECT 3.790 2.805 3.800 3.015 ;
        RECT 3.800 2.805 3.810 3.005 ;
        RECT 3.810 2.805 3.820 2.995 ;
        RECT 3.820 2.805 3.830 2.985 ;
        RECT 3.830 2.805 3.840 2.975 ;
        RECT 3.705 2.865 3.715 3.035 ;
        RECT 3.715 2.855 3.725 3.035 ;
        RECT 3.725 2.845 3.735 3.035 ;
        RECT 3.735 2.835 3.745 3.035 ;
        RECT 3.745 2.825 3.755 3.035 ;
        RECT 3.755 2.815 3.765 3.035 ;
        RECT 3.775 1.685 4.075 2.225 ;
        RECT 3.775 2.055 5.090 2.225 ;
        RECT 4.915 2.055 5.090 2.275 ;
        RECT 5.060 1.125 5.230 1.295 ;
        RECT 5.395 1.125 5.400 2.095 ;
        RECT 6.430 1.525 6.600 2.095 ;
        RECT 5.395 1.925 6.600 2.095 ;
        RECT 5.230 1.125 5.240 2.249 ;
        RECT 5.240 1.125 5.250 2.239 ;
        RECT 5.250 1.125 5.260 2.229 ;
        RECT 5.260 1.125 5.270 2.219 ;
        RECT 5.270 1.125 5.280 2.209 ;
        RECT 5.280 1.125 5.290 2.199 ;
        RECT 5.290 1.125 5.300 2.189 ;
        RECT 5.300 1.125 5.310 2.179 ;
        RECT 5.310 1.125 5.320 2.169 ;
        RECT 5.320 1.125 5.330 2.159 ;
        RECT 5.330 1.125 5.340 2.149 ;
        RECT 5.340 1.125 5.350 2.139 ;
        RECT 5.350 1.125 5.360 2.129 ;
        RECT 5.360 1.125 5.370 2.119 ;
        RECT 5.370 1.125 5.380 2.109 ;
        RECT 5.380 1.125 5.390 2.099 ;
        RECT 5.390 1.125 5.396 2.095 ;
        RECT 5.215 1.930 5.225 2.264 ;
        RECT 5.225 1.920 5.231 2.260 ;
        RECT 5.090 2.055 5.100 2.275 ;
        RECT 5.100 2.045 5.110 2.275 ;
        RECT 5.110 2.035 5.120 2.275 ;
        RECT 5.120 2.025 5.130 2.275 ;
        RECT 5.130 2.015 5.140 2.275 ;
        RECT 5.140 2.005 5.150 2.275 ;
        RECT 5.150 1.995 5.160 2.275 ;
        RECT 5.160 1.985 5.170 2.275 ;
        RECT 5.170 1.975 5.180 2.275 ;
        RECT 5.180 1.965 5.190 2.275 ;
        RECT 5.190 1.955 5.200 2.275 ;
        RECT 5.200 1.945 5.210 2.275 ;
        RECT 5.210 1.935 5.216 2.275 ;
        RECT 1.720 0.995 1.890 2.685 ;
        RECT 1.440 2.350 1.890 2.685 ;
        RECT 2.765 0.525 2.935 2.685 ;
        RECT 2.765 1.795 3.135 1.965 ;
        RECT 1.440 2.515 3.490 2.685 ;
        RECT 3.550 2.455 3.570 2.685 ;
        RECT 2.765 0.525 3.595 0.695 ;
        RECT 3.630 2.455 4.650 2.625 ;
        RECT 4.660 2.455 4.810 2.635 ;
        RECT 4.820 2.465 5.305 2.635 ;
        RECT 5.630 2.275 6.735 2.445 ;
        RECT 6.950 1.265 7.150 1.435 ;
        RECT 7.185 2.535 7.355 2.825 ;
        RECT 7.075 2.535 7.355 2.705 ;
        RECT 7.185 2.655 7.660 2.825 ;
        RECT 6.995 2.465 7.005 2.705 ;
        RECT 7.005 2.475 7.015 2.705 ;
        RECT 7.015 2.485 7.025 2.705 ;
        RECT 7.025 2.495 7.035 2.705 ;
        RECT 7.035 2.505 7.045 2.705 ;
        RECT 7.045 2.515 7.055 2.705 ;
        RECT 7.055 2.525 7.065 2.705 ;
        RECT 7.065 2.535 7.075 2.705 ;
        RECT 6.950 2.420 6.960 2.660 ;
        RECT 6.960 2.430 6.970 2.670 ;
        RECT 6.970 2.440 6.980 2.680 ;
        RECT 6.980 2.450 6.990 2.690 ;
        RECT 6.990 2.455 6.996 2.699 ;
        RECT 6.780 1.265 6.790 2.489 ;
        RECT 6.790 1.265 6.800 2.499 ;
        RECT 6.800 1.265 6.810 2.509 ;
        RECT 6.810 1.265 6.820 2.519 ;
        RECT 6.820 1.265 6.830 2.529 ;
        RECT 6.830 1.265 6.840 2.539 ;
        RECT 6.840 1.265 6.850 2.549 ;
        RECT 6.850 1.265 6.860 2.559 ;
        RECT 6.860 1.265 6.870 2.569 ;
        RECT 6.870 1.265 6.880 2.579 ;
        RECT 6.880 1.265 6.890 2.589 ;
        RECT 6.890 1.265 6.900 2.599 ;
        RECT 6.900 1.265 6.910 2.609 ;
        RECT 6.910 1.265 6.920 2.619 ;
        RECT 6.920 1.265 6.930 2.629 ;
        RECT 6.930 1.265 6.940 2.639 ;
        RECT 6.940 1.265 6.950 2.649 ;
        RECT 6.735 2.275 6.745 2.445 ;
        RECT 6.745 2.275 6.755 2.455 ;
        RECT 6.755 2.275 6.765 2.465 ;
        RECT 6.765 2.275 6.775 2.475 ;
        RECT 6.775 2.275 6.781 2.485 ;
        RECT 5.495 2.275 5.505 2.569 ;
        RECT 5.505 2.275 5.515 2.559 ;
        RECT 5.515 2.275 5.525 2.549 ;
        RECT 5.525 2.275 5.535 2.539 ;
        RECT 5.535 2.275 5.545 2.529 ;
        RECT 5.545 2.275 5.555 2.519 ;
        RECT 5.555 2.275 5.565 2.509 ;
        RECT 5.565 2.275 5.575 2.499 ;
        RECT 5.575 2.275 5.585 2.489 ;
        RECT 5.585 2.275 5.595 2.479 ;
        RECT 5.595 2.275 5.605 2.469 ;
        RECT 5.605 2.275 5.615 2.459 ;
        RECT 5.615 2.275 5.625 2.449 ;
        RECT 5.625 2.275 5.631 2.445 ;
        RECT 5.440 2.330 5.450 2.624 ;
        RECT 5.450 2.320 5.460 2.614 ;
        RECT 5.460 2.310 5.470 2.604 ;
        RECT 5.470 2.300 5.480 2.594 ;
        RECT 5.480 2.290 5.490 2.584 ;
        RECT 5.490 2.280 5.496 2.580 ;
        RECT 5.305 2.465 5.315 2.635 ;
        RECT 5.315 2.455 5.325 2.635 ;
        RECT 5.325 2.445 5.335 2.635 ;
        RECT 5.335 2.435 5.345 2.635 ;
        RECT 5.345 2.425 5.355 2.635 ;
        RECT 5.355 2.415 5.365 2.635 ;
        RECT 5.365 2.405 5.375 2.635 ;
        RECT 5.375 2.395 5.385 2.635 ;
        RECT 5.385 2.385 5.395 2.635 ;
        RECT 5.395 2.375 5.405 2.635 ;
        RECT 5.405 2.365 5.415 2.635 ;
        RECT 5.415 2.355 5.425 2.635 ;
        RECT 5.425 2.345 5.435 2.635 ;
        RECT 5.435 2.335 5.441 2.635 ;
        RECT 4.810 2.465 4.820 2.635 ;
        RECT 4.650 2.455 4.660 2.625 ;
        RECT 3.570 2.455 3.580 2.675 ;
        RECT 3.580 2.455 3.590 2.665 ;
        RECT 3.590 2.455 3.600 2.655 ;
        RECT 3.600 2.455 3.610 2.645 ;
        RECT 3.610 2.455 3.620 2.635 ;
        RECT 3.620 2.455 3.630 2.625 ;
        RECT 3.490 2.515 3.500 2.685 ;
        RECT 3.500 2.505 3.510 2.685 ;
        RECT 3.510 2.495 3.520 2.685 ;
        RECT 3.520 2.485 3.530 2.685 ;
        RECT 3.530 2.475 3.540 2.685 ;
        RECT 3.540 2.465 3.550 2.685 ;
        RECT 9.165 1.125 9.335 2.215 ;
        RECT 8.305 2.045 9.335 2.215 ;
        RECT 9.070 1.125 9.370 1.295 ;
        RECT 8.135 1.885 8.145 2.215 ;
        RECT 8.145 1.895 8.155 2.215 ;
        RECT 8.155 1.905 8.165 2.215 ;
        RECT 8.165 1.915 8.175 2.215 ;
        RECT 8.175 1.925 8.185 2.215 ;
        RECT 8.185 1.935 8.195 2.215 ;
        RECT 8.195 1.945 8.205 2.215 ;
        RECT 8.205 1.955 8.215 2.215 ;
        RECT 8.215 1.965 8.225 2.215 ;
        RECT 8.225 1.975 8.235 2.215 ;
        RECT 8.235 1.985 8.245 2.215 ;
        RECT 8.245 1.995 8.255 2.215 ;
        RECT 8.255 2.005 8.265 2.215 ;
        RECT 8.265 2.015 8.275 2.215 ;
        RECT 8.275 2.025 8.285 2.215 ;
        RECT 8.285 2.035 8.295 2.215 ;
        RECT 8.295 2.045 8.305 2.215 ;
        RECT 8.090 1.840 8.100 2.170 ;
        RECT 8.100 1.850 8.110 2.180 ;
        RECT 8.110 1.860 8.120 2.190 ;
        RECT 8.120 1.870 8.130 2.200 ;
        RECT 8.130 1.875 8.136 2.209 ;
        RECT 7.790 1.675 7.800 1.869 ;
        RECT 7.800 1.675 7.810 1.879 ;
        RECT 7.810 1.675 7.820 1.889 ;
        RECT 7.820 1.675 7.830 1.899 ;
        RECT 7.830 1.675 7.840 1.909 ;
        RECT 7.840 1.675 7.850 1.919 ;
        RECT 7.850 1.675 7.860 1.929 ;
        RECT 7.860 1.675 7.870 1.939 ;
        RECT 7.870 1.675 7.880 1.949 ;
        RECT 7.880 1.675 7.890 1.959 ;
        RECT 7.890 1.675 7.900 1.969 ;
        RECT 7.900 1.675 7.910 1.979 ;
        RECT 7.910 1.675 7.920 1.989 ;
        RECT 7.920 1.675 7.930 1.999 ;
        RECT 7.930 1.675 7.940 2.009 ;
        RECT 7.940 1.675 7.950 2.019 ;
        RECT 7.950 1.675 7.960 2.029 ;
        RECT 7.960 1.675 7.970 2.039 ;
        RECT 7.970 1.675 7.980 2.049 ;
        RECT 7.980 1.675 7.990 2.059 ;
        RECT 7.990 1.675 8.000 2.069 ;
        RECT 8.000 1.675 8.010 2.079 ;
        RECT 8.010 1.675 8.020 2.089 ;
        RECT 8.020 1.675 8.030 2.099 ;
        RECT 8.030 1.675 8.040 2.109 ;
        RECT 8.040 1.675 8.050 2.119 ;
        RECT 8.050 1.675 8.060 2.129 ;
        RECT 8.060 1.675 8.070 2.139 ;
        RECT 8.070 1.675 8.080 2.149 ;
        RECT 8.080 1.675 8.090 2.159 ;
        RECT 4.645 0.730 4.815 1.400 ;
        RECT 5.660 0.730 5.830 1.065 ;
        RECT 4.645 0.730 5.830 0.900 ;
        RECT 6.760 0.545 6.930 1.065 ;
        RECT 5.660 0.895 6.930 1.065 ;
        RECT 6.760 0.545 7.850 0.715 ;
        RECT 7.680 0.545 7.850 1.145 ;
        RECT 8.685 0.745 8.855 1.145 ;
        RECT 7.680 0.975 8.855 1.145 ;
        RECT 9.550 0.745 9.720 2.215 ;
        RECT 8.685 0.745 10.170 0.945 ;
        RECT 9.550 2.045 10.170 2.215 ;
        RECT 7.110 0.895 7.500 1.065 ;
        RECT 7.330 0.895 7.500 2.335 ;
        RECT 7.130 2.165 7.680 2.335 ;
        RECT 8.720 2.395 9.020 2.705 ;
        RECT 10.410 1.610 10.580 2.565 ;
        RECT 8.000 2.395 10.580 2.565 ;
        RECT 10.410 1.610 10.830 1.780 ;
        RECT 7.910 2.315 7.920 2.565 ;
        RECT 7.920 2.325 7.930 2.565 ;
        RECT 7.930 2.335 7.940 2.565 ;
        RECT 7.940 2.345 7.950 2.565 ;
        RECT 7.950 2.355 7.960 2.565 ;
        RECT 7.960 2.365 7.970 2.565 ;
        RECT 7.970 2.375 7.980 2.565 ;
        RECT 7.980 2.385 7.990 2.565 ;
        RECT 7.990 2.395 8.000 2.565 ;
        RECT 7.770 2.175 7.780 2.425 ;
        RECT 7.780 2.185 7.790 2.435 ;
        RECT 7.790 2.195 7.800 2.445 ;
        RECT 7.800 2.205 7.810 2.455 ;
        RECT 7.810 2.215 7.820 2.465 ;
        RECT 7.820 2.225 7.830 2.475 ;
        RECT 7.830 2.235 7.840 2.485 ;
        RECT 7.840 2.245 7.850 2.495 ;
        RECT 7.850 2.255 7.860 2.505 ;
        RECT 7.860 2.265 7.870 2.515 ;
        RECT 7.870 2.275 7.880 2.525 ;
        RECT 7.880 2.285 7.890 2.535 ;
        RECT 7.890 2.295 7.900 2.545 ;
        RECT 7.900 2.305 7.910 2.555 ;
        RECT 7.680 2.165 7.690 2.335 ;
        RECT 7.690 2.165 7.700 2.345 ;
        RECT 7.700 2.165 7.710 2.355 ;
        RECT 7.710 2.165 7.720 2.365 ;
        RECT 7.720 2.165 7.730 2.375 ;
        RECT 7.730 2.165 7.740 2.385 ;
        RECT 7.740 2.165 7.750 2.395 ;
        RECT 7.750 2.165 7.760 2.405 ;
        RECT 7.760 2.165 7.770 2.415 ;
  END 
END FFDSRHQHDMXHT

MACRO FFDSRHQHD3XHT
  CLASS  CORE ;
  FOREIGN FFDSRHQHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.400 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 14.755 0.785 15.055 1.405 ;
        RECT 14.755 1.980 15.055 2.960 ;
        RECT 14.755 1.235 16.095 1.405 ;
        RECT 15.415 1.235 16.095 2.435 ;
        RECT 14.755 1.980 16.095 2.435 ;
        RECT 15.795 0.720 16.095 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.670 1.600 3.180 2.020 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 13.630 1.260 14.100 1.790 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 0.965 ;
        RECT 1.145 -0.300 1.445 0.965 ;
        RECT 2.715 -0.300 3.015 1.230 ;
        RECT 4.575 -0.300 4.875 1.055 ;
        RECT 8.010 -0.300 8.310 0.435 ;
        RECT 9.155 -0.300 9.455 0.435 ;
        RECT 11.765 -0.300 12.065 0.715 ;
        RECT 14.235 -0.300 14.535 1.055 ;
        RECT 15.275 -0.300 15.575 1.055 ;
        RECT 0.000 -0.300 16.400 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 1.090 1.230 1.665 1.700 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 12.275 2.885 12.905 3.185 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.280 0.860 3.990 ;
        RECT 1.675 2.965 1.975 3.990 ;
        RECT 2.685 2.965 2.985 3.990 ;
        RECT 4.490 3.095 4.790 3.990 ;
        RECT 6.600 3.095 6.900 3.990 ;
        RECT 7.575 3.025 7.875 3.990 ;
        RECT 8.675 2.900 8.975 3.990 ;
        RECT 11.765 2.845 12.065 3.990 ;
        RECT 13.175 2.825 13.475 3.990 ;
        RECT 14.235 2.975 14.535 3.990 ;
        RECT 15.275 2.635 15.575 3.990 ;
        RECT 0.000 3.390 16.400 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 2.280 0.340 3.175 ;
        RECT 0.105 3.005 0.405 3.175 ;
        RECT 1.665 0.795 2.020 0.965 ;
        RECT 1.850 0.795 2.020 1.700 ;
        RECT 1.850 1.400 2.080 1.700 ;
        RECT 3.710 2.135 3.825 2.435 ;
        RECT 4.025 1.325 4.965 1.495 ;
        RECT 4.795 1.325 4.965 1.845 ;
        RECT 4.795 1.675 5.895 1.845 ;
        RECT 3.935 1.325 3.945 2.385 ;
        RECT 3.945 1.325 3.955 2.375 ;
        RECT 3.955 1.325 3.965 2.365 ;
        RECT 3.965 1.325 3.975 2.355 ;
        RECT 3.975 1.325 3.985 2.345 ;
        RECT 3.985 1.325 3.995 2.335 ;
        RECT 3.995 1.325 4.005 2.325 ;
        RECT 4.005 1.325 4.015 2.315 ;
        RECT 4.015 1.325 4.025 2.305 ;
        RECT 3.895 1.295 3.905 2.425 ;
        RECT 3.905 1.305 3.915 2.415 ;
        RECT 3.915 1.315 3.925 2.405 ;
        RECT 3.925 1.325 3.935 2.395 ;
        RECT 3.855 1.255 3.865 2.435 ;
        RECT 3.865 1.265 3.875 2.435 ;
        RECT 3.875 1.275 3.885 2.435 ;
        RECT 3.885 1.285 3.895 2.435 ;
        RECT 3.840 1.240 3.850 1.480 ;
        RECT 3.850 1.245 3.856 1.489 ;
        RECT 3.825 2.135 3.835 2.435 ;
        RECT 3.835 2.125 3.845 2.435 ;
        RECT 3.845 2.115 3.855 2.435 ;
        RECT 3.670 0.995 3.680 1.309 ;
        RECT 3.680 0.995 3.690 1.319 ;
        RECT 3.690 0.995 3.700 1.329 ;
        RECT 3.700 0.995 3.710 1.339 ;
        RECT 3.710 0.995 3.720 1.349 ;
        RECT 3.720 0.995 3.730 1.359 ;
        RECT 3.730 0.995 3.740 1.369 ;
        RECT 3.740 0.995 3.750 1.379 ;
        RECT 3.750 0.995 3.760 1.389 ;
        RECT 3.760 0.995 3.770 1.399 ;
        RECT 3.770 0.995 3.780 1.409 ;
        RECT 3.780 0.995 3.790 1.419 ;
        RECT 3.790 0.995 3.800 1.429 ;
        RECT 3.800 0.995 3.810 1.439 ;
        RECT 3.810 0.995 3.820 1.449 ;
        RECT 3.820 0.995 3.830 1.459 ;
        RECT 3.830 0.995 3.840 1.469 ;
        RECT 5.155 0.775 5.455 1.085 ;
        RECT 5.155 0.775 7.645 0.945 ;
        RECT 4.315 1.675 4.615 2.215 ;
        RECT 6.075 1.125 6.245 2.215 ;
        RECT 4.315 2.045 6.870 2.215 ;
        RECT 6.945 1.970 6.950 2.215 ;
        RECT 5.695 1.125 7.095 1.295 ;
        RECT 7.025 1.970 7.425 2.140 ;
        RECT 7.860 1.495 9.185 1.665 ;
        RECT 7.715 1.495 7.725 1.799 ;
        RECT 7.725 1.495 7.735 1.789 ;
        RECT 7.735 1.495 7.745 1.779 ;
        RECT 7.745 1.495 7.755 1.769 ;
        RECT 7.755 1.495 7.765 1.759 ;
        RECT 7.765 1.495 7.775 1.749 ;
        RECT 7.775 1.495 7.785 1.739 ;
        RECT 7.785 1.495 7.795 1.729 ;
        RECT 7.795 1.495 7.805 1.719 ;
        RECT 7.805 1.495 7.815 1.709 ;
        RECT 7.815 1.495 7.825 1.699 ;
        RECT 7.825 1.495 7.835 1.689 ;
        RECT 7.835 1.495 7.845 1.679 ;
        RECT 7.845 1.495 7.855 1.669 ;
        RECT 7.855 1.495 7.861 1.665 ;
        RECT 7.595 1.685 7.605 1.919 ;
        RECT 7.605 1.675 7.615 1.909 ;
        RECT 7.615 1.665 7.625 1.899 ;
        RECT 7.625 1.655 7.635 1.889 ;
        RECT 7.635 1.645 7.645 1.879 ;
        RECT 7.645 1.635 7.655 1.869 ;
        RECT 7.655 1.625 7.665 1.859 ;
        RECT 7.665 1.615 7.675 1.849 ;
        RECT 7.675 1.605 7.685 1.839 ;
        RECT 7.685 1.595 7.695 1.829 ;
        RECT 7.695 1.585 7.705 1.819 ;
        RECT 7.705 1.575 7.715 1.809 ;
        RECT 7.425 1.855 7.435 2.139 ;
        RECT 7.435 1.845 7.445 2.139 ;
        RECT 7.445 1.835 7.455 2.139 ;
        RECT 7.455 1.825 7.465 2.139 ;
        RECT 7.465 1.815 7.475 2.139 ;
        RECT 7.475 1.805 7.485 2.139 ;
        RECT 7.485 1.795 7.495 2.139 ;
        RECT 7.495 1.785 7.505 2.139 ;
        RECT 7.505 1.775 7.515 2.139 ;
        RECT 7.515 1.765 7.525 2.139 ;
        RECT 7.525 1.755 7.535 2.139 ;
        RECT 7.535 1.745 7.545 2.139 ;
        RECT 7.545 1.735 7.555 2.139 ;
        RECT 7.555 1.725 7.565 2.139 ;
        RECT 7.565 1.715 7.575 2.139 ;
        RECT 7.575 1.705 7.585 2.139 ;
        RECT 7.585 1.695 7.595 2.139 ;
        RECT 6.950 1.970 6.960 2.204 ;
        RECT 6.960 1.970 6.970 2.194 ;
        RECT 6.970 1.970 6.980 2.184 ;
        RECT 6.980 1.970 6.990 2.174 ;
        RECT 6.990 1.970 7.000 2.164 ;
        RECT 7.000 1.970 7.010 2.154 ;
        RECT 7.010 1.970 7.020 2.144 ;
        RECT 7.020 1.970 7.026 2.140 ;
        RECT 6.870 2.045 6.880 2.215 ;
        RECT 6.880 2.035 6.890 2.215 ;
        RECT 6.890 2.025 6.900 2.215 ;
        RECT 6.900 2.015 6.910 2.215 ;
        RECT 6.910 2.005 6.920 2.215 ;
        RECT 6.920 1.995 6.930 2.215 ;
        RECT 6.930 1.985 6.940 2.215 ;
        RECT 6.940 1.975 6.946 2.215 ;
        RECT 0.690 1.030 0.860 2.100 ;
        RECT 0.690 1.930 1.335 2.100 ;
        RECT 1.165 1.930 1.335 2.625 ;
        RECT 1.645 2.455 1.815 2.785 ;
        RECT 1.165 2.455 1.815 2.625 ;
        RECT 1.645 2.615 3.060 2.785 ;
        RECT 3.355 2.975 4.110 3.145 ;
        RECT 4.415 2.745 7.355 2.915 ;
        RECT 8.325 2.545 8.495 2.840 ;
        RECT 7.505 2.670 8.495 2.840 ;
        RECT 8.325 2.545 9.565 2.715 ;
        RECT 9.395 2.545 9.565 3.085 ;
        RECT 9.395 2.915 9.705 3.085 ;
        RECT 7.430 2.670 7.440 2.904 ;
        RECT 7.440 2.670 7.450 2.894 ;
        RECT 7.450 2.670 7.460 2.884 ;
        RECT 7.460 2.670 7.470 2.874 ;
        RECT 7.470 2.670 7.480 2.864 ;
        RECT 7.480 2.670 7.490 2.854 ;
        RECT 7.490 2.670 7.500 2.844 ;
        RECT 7.500 2.670 7.506 2.840 ;
        RECT 7.355 2.745 7.365 2.915 ;
        RECT 7.365 2.735 7.375 2.915 ;
        RECT 7.375 2.725 7.385 2.915 ;
        RECT 7.385 2.715 7.395 2.915 ;
        RECT 7.395 2.705 7.405 2.915 ;
        RECT 7.405 2.695 7.415 2.915 ;
        RECT 7.415 2.685 7.425 2.915 ;
        RECT 7.425 2.675 7.431 2.915 ;
        RECT 4.340 2.745 4.350 2.979 ;
        RECT 4.350 2.745 4.360 2.969 ;
        RECT 4.360 2.745 4.370 2.959 ;
        RECT 4.370 2.745 4.380 2.949 ;
        RECT 4.380 2.745 4.390 2.939 ;
        RECT 4.390 2.745 4.400 2.929 ;
        RECT 4.400 2.745 4.410 2.919 ;
        RECT 4.410 2.745 4.416 2.915 ;
        RECT 4.185 2.900 4.195 3.134 ;
        RECT 4.195 2.890 4.205 3.124 ;
        RECT 4.205 2.880 4.215 3.114 ;
        RECT 4.215 2.870 4.225 3.104 ;
        RECT 4.225 2.860 4.235 3.094 ;
        RECT 4.235 2.850 4.245 3.084 ;
        RECT 4.245 2.840 4.255 3.074 ;
        RECT 4.255 2.830 4.265 3.064 ;
        RECT 4.265 2.820 4.275 3.054 ;
        RECT 4.275 2.810 4.285 3.044 ;
        RECT 4.285 2.800 4.295 3.034 ;
        RECT 4.295 2.790 4.305 3.024 ;
        RECT 4.305 2.780 4.315 3.014 ;
        RECT 4.315 2.770 4.325 3.004 ;
        RECT 4.325 2.760 4.335 2.994 ;
        RECT 4.335 2.750 4.341 2.990 ;
        RECT 4.110 2.975 4.120 3.145 ;
        RECT 4.120 2.965 4.130 3.145 ;
        RECT 4.130 2.955 4.140 3.145 ;
        RECT 4.140 2.945 4.150 3.145 ;
        RECT 4.150 2.935 4.160 3.145 ;
        RECT 4.160 2.925 4.170 3.145 ;
        RECT 4.170 2.915 4.180 3.145 ;
        RECT 4.180 2.905 4.186 3.145 ;
        RECT 3.185 2.675 3.195 3.145 ;
        RECT 3.195 2.685 3.205 3.145 ;
        RECT 3.205 2.695 3.215 3.145 ;
        RECT 3.215 2.705 3.225 3.145 ;
        RECT 3.225 2.715 3.235 3.145 ;
        RECT 3.235 2.725 3.245 3.145 ;
        RECT 3.245 2.735 3.255 3.145 ;
        RECT 3.255 2.745 3.265 3.145 ;
        RECT 3.265 2.755 3.275 3.145 ;
        RECT 3.275 2.765 3.285 3.145 ;
        RECT 3.285 2.775 3.295 3.145 ;
        RECT 3.295 2.785 3.305 3.145 ;
        RECT 3.305 2.795 3.315 3.145 ;
        RECT 3.315 2.805 3.325 3.145 ;
        RECT 3.325 2.815 3.335 3.145 ;
        RECT 3.335 2.825 3.345 3.145 ;
        RECT 3.345 2.835 3.355 3.145 ;
        RECT 3.135 2.625 3.145 2.859 ;
        RECT 3.145 2.635 3.155 2.869 ;
        RECT 3.155 2.645 3.165 2.879 ;
        RECT 3.165 2.655 3.175 2.889 ;
        RECT 3.175 2.665 3.185 2.899 ;
        RECT 3.060 2.615 3.070 2.785 ;
        RECT 3.070 2.615 3.080 2.795 ;
        RECT 3.080 2.615 3.090 2.805 ;
        RECT 3.090 2.615 3.100 2.815 ;
        RECT 3.100 2.615 3.110 2.825 ;
        RECT 3.110 2.615 3.120 2.835 ;
        RECT 3.120 2.615 3.130 2.845 ;
        RECT 3.130 2.615 3.136 2.855 ;
        RECT 10.265 2.195 10.435 2.505 ;
        RECT 8.125 2.195 10.435 2.365 ;
        RECT 10.265 2.335 10.565 2.505 ;
        RECT 8.560 0.965 9.535 1.135 ;
        RECT 9.365 0.965 9.535 1.485 ;
        RECT 10.295 1.180 10.465 1.485 ;
        RECT 9.365 1.315 10.465 1.485 ;
        RECT 10.295 1.180 10.595 1.350 ;
        RECT 1.795 1.945 2.430 2.115 ;
        RECT 2.260 0.995 2.430 2.400 ;
        RECT 2.165 1.945 2.430 2.400 ;
        RECT 2.165 2.230 3.305 2.400 ;
        RECT 3.530 1.785 3.675 1.955 ;
        RECT 3.645 2.625 3.960 2.795 ;
        RECT 3.475 0.515 4.185 0.685 ;
        RECT 4.265 2.395 7.130 2.565 ;
        RECT 7.205 2.320 7.225 2.565 ;
        RECT 7.300 2.320 7.775 2.490 ;
        RECT 7.935 1.845 7.945 2.490 ;
        RECT 9.365 1.675 9.535 2.015 ;
        RECT 8.010 1.845 9.535 2.015 ;
        RECT 9.365 1.675 10.720 1.845 ;
        RECT 11.305 2.115 11.365 2.285 ;
        RECT 11.065 1.885 11.075 2.285 ;
        RECT 11.075 1.895 11.085 2.285 ;
        RECT 11.085 1.905 11.095 2.285 ;
        RECT 11.095 1.915 11.105 2.285 ;
        RECT 11.105 1.925 11.115 2.285 ;
        RECT 11.115 1.935 11.125 2.285 ;
        RECT 11.125 1.945 11.135 2.285 ;
        RECT 11.135 1.955 11.145 2.285 ;
        RECT 11.145 1.965 11.155 2.285 ;
        RECT 11.155 1.975 11.165 2.285 ;
        RECT 11.165 1.985 11.175 2.285 ;
        RECT 11.175 1.995 11.185 2.285 ;
        RECT 11.185 2.005 11.195 2.285 ;
        RECT 11.195 2.015 11.205 2.285 ;
        RECT 11.205 2.025 11.215 2.285 ;
        RECT 11.215 2.035 11.225 2.285 ;
        RECT 11.225 2.045 11.235 2.285 ;
        RECT 11.235 2.055 11.245 2.285 ;
        RECT 11.245 2.065 11.255 2.285 ;
        RECT 11.255 2.075 11.265 2.285 ;
        RECT 11.265 2.085 11.275 2.285 ;
        RECT 11.275 2.095 11.285 2.285 ;
        RECT 11.285 2.105 11.295 2.285 ;
        RECT 11.295 2.115 11.305 2.285 ;
        RECT 10.865 1.685 10.875 1.989 ;
        RECT 10.875 1.695 10.885 1.999 ;
        RECT 10.885 1.705 10.895 2.009 ;
        RECT 10.895 1.715 10.905 2.019 ;
        RECT 10.905 1.725 10.915 2.029 ;
        RECT 10.915 1.735 10.925 2.039 ;
        RECT 10.925 1.745 10.935 2.049 ;
        RECT 10.935 1.755 10.945 2.059 ;
        RECT 10.945 1.765 10.955 2.069 ;
        RECT 10.955 1.775 10.965 2.079 ;
        RECT 10.965 1.785 10.975 2.089 ;
        RECT 10.975 1.795 10.985 2.099 ;
        RECT 10.985 1.805 10.995 2.109 ;
        RECT 10.995 1.815 11.005 2.119 ;
        RECT 11.005 1.825 11.015 2.129 ;
        RECT 11.015 1.835 11.025 2.139 ;
        RECT 11.025 1.845 11.035 2.149 ;
        RECT 11.035 1.855 11.045 2.159 ;
        RECT 11.045 1.865 11.055 2.169 ;
        RECT 11.055 1.875 11.065 2.179 ;
        RECT 10.720 1.675 10.730 1.845 ;
        RECT 10.730 1.675 10.740 1.855 ;
        RECT 10.740 1.675 10.750 1.865 ;
        RECT 10.750 1.675 10.760 1.875 ;
        RECT 10.760 1.675 10.770 1.885 ;
        RECT 10.770 1.675 10.780 1.895 ;
        RECT 10.780 1.675 10.790 1.905 ;
        RECT 10.790 1.675 10.800 1.915 ;
        RECT 10.800 1.675 10.810 1.925 ;
        RECT 10.810 1.675 10.820 1.935 ;
        RECT 10.820 1.675 10.830 1.945 ;
        RECT 10.830 1.675 10.840 1.955 ;
        RECT 10.840 1.675 10.850 1.965 ;
        RECT 10.850 1.675 10.860 1.975 ;
        RECT 10.860 1.675 10.866 1.985 ;
        RECT 7.945 1.845 7.955 2.069 ;
        RECT 7.955 1.845 7.965 2.059 ;
        RECT 7.965 1.845 7.975 2.049 ;
        RECT 7.975 1.845 7.985 2.039 ;
        RECT 7.985 1.845 7.995 2.029 ;
        RECT 7.995 1.845 8.005 2.019 ;
        RECT 8.005 1.845 8.011 2.015 ;
        RECT 7.775 2.005 7.785 2.489 ;
        RECT 7.785 1.995 7.795 2.489 ;
        RECT 7.795 1.985 7.805 2.489 ;
        RECT 7.805 1.975 7.815 2.489 ;
        RECT 7.815 1.965 7.825 2.489 ;
        RECT 7.825 1.955 7.835 2.489 ;
        RECT 7.835 1.945 7.845 2.489 ;
        RECT 7.845 1.935 7.855 2.489 ;
        RECT 7.855 1.925 7.865 2.489 ;
        RECT 7.865 1.915 7.875 2.489 ;
        RECT 7.875 1.905 7.885 2.489 ;
        RECT 7.885 1.895 7.895 2.489 ;
        RECT 7.895 1.885 7.905 2.489 ;
        RECT 7.905 1.875 7.915 2.489 ;
        RECT 7.915 1.865 7.925 2.489 ;
        RECT 7.925 1.855 7.935 2.489 ;
        RECT 7.225 2.320 7.235 2.554 ;
        RECT 7.235 2.320 7.245 2.544 ;
        RECT 7.245 2.320 7.255 2.534 ;
        RECT 7.255 2.320 7.265 2.524 ;
        RECT 7.265 2.320 7.275 2.514 ;
        RECT 7.275 2.320 7.285 2.504 ;
        RECT 7.285 2.320 7.295 2.494 ;
        RECT 7.295 2.320 7.301 2.490 ;
        RECT 7.130 2.395 7.140 2.565 ;
        RECT 7.140 2.385 7.150 2.565 ;
        RECT 7.150 2.375 7.160 2.565 ;
        RECT 7.160 2.365 7.170 2.565 ;
        RECT 7.170 2.355 7.180 2.565 ;
        RECT 7.180 2.345 7.190 2.565 ;
        RECT 7.190 2.335 7.200 2.565 ;
        RECT 7.200 2.325 7.206 2.565 ;
        RECT 4.190 2.395 4.200 2.629 ;
        RECT 4.200 2.395 4.210 2.619 ;
        RECT 4.210 2.395 4.220 2.609 ;
        RECT 4.220 2.395 4.230 2.599 ;
        RECT 4.230 2.395 4.240 2.589 ;
        RECT 4.240 2.395 4.250 2.579 ;
        RECT 4.250 2.395 4.260 2.569 ;
        RECT 4.260 2.395 4.266 2.565 ;
        RECT 4.035 2.550 4.045 2.784 ;
        RECT 4.045 2.540 4.055 2.774 ;
        RECT 4.055 2.530 4.065 2.764 ;
        RECT 4.065 2.520 4.075 2.754 ;
        RECT 4.075 2.510 4.085 2.744 ;
        RECT 4.085 2.500 4.095 2.734 ;
        RECT 4.095 2.490 4.105 2.724 ;
        RECT 4.105 2.480 4.115 2.714 ;
        RECT 4.115 2.470 4.125 2.704 ;
        RECT 4.125 2.460 4.135 2.694 ;
        RECT 4.135 2.450 4.145 2.684 ;
        RECT 4.145 2.440 4.155 2.674 ;
        RECT 4.155 2.430 4.165 2.664 ;
        RECT 4.165 2.420 4.175 2.654 ;
        RECT 4.175 2.410 4.185 2.644 ;
        RECT 4.185 2.400 4.191 2.640 ;
        RECT 3.960 2.625 3.970 2.795 ;
        RECT 3.970 2.615 3.980 2.795 ;
        RECT 3.980 2.605 3.990 2.795 ;
        RECT 3.990 2.595 4.000 2.795 ;
        RECT 4.000 2.585 4.010 2.795 ;
        RECT 4.010 2.575 4.020 2.795 ;
        RECT 4.020 2.565 4.030 2.795 ;
        RECT 4.030 2.555 4.036 2.795 ;
        RECT 3.570 2.560 3.580 2.794 ;
        RECT 3.580 2.570 3.590 2.794 ;
        RECT 3.590 2.580 3.600 2.794 ;
        RECT 3.600 2.590 3.610 2.794 ;
        RECT 3.610 2.600 3.620 2.794 ;
        RECT 3.620 2.610 3.630 2.794 ;
        RECT 3.630 2.620 3.640 2.794 ;
        RECT 3.640 2.625 3.646 2.795 ;
        RECT 3.530 2.520 3.540 2.754 ;
        RECT 3.540 2.530 3.550 2.764 ;
        RECT 3.550 2.540 3.560 2.774 ;
        RECT 3.560 2.550 3.570 2.784 ;
        RECT 3.475 1.405 3.485 2.699 ;
        RECT 3.485 1.415 3.495 2.709 ;
        RECT 3.495 1.425 3.505 2.719 ;
        RECT 3.505 1.435 3.515 2.729 ;
        RECT 3.515 1.445 3.525 2.739 ;
        RECT 3.525 1.450 3.531 2.750 ;
        RECT 3.360 0.515 3.370 2.585 ;
        RECT 3.370 0.515 3.380 2.595 ;
        RECT 3.380 0.515 3.390 2.605 ;
        RECT 3.390 0.515 3.400 2.615 ;
        RECT 3.400 0.515 3.410 2.625 ;
        RECT 3.410 0.515 3.420 2.635 ;
        RECT 3.420 0.515 3.430 2.645 ;
        RECT 3.430 0.515 3.440 2.655 ;
        RECT 3.440 0.515 3.450 2.665 ;
        RECT 3.450 0.515 3.460 2.675 ;
        RECT 3.460 0.515 3.470 2.685 ;
        RECT 3.470 0.515 3.476 2.695 ;
        RECT 3.305 0.515 3.315 1.469 ;
        RECT 3.315 0.515 3.325 1.479 ;
        RECT 3.325 0.515 3.335 1.489 ;
        RECT 3.335 0.515 3.345 1.499 ;
        RECT 3.345 0.515 3.355 1.509 ;
        RECT 3.355 0.515 3.361 1.519 ;
        RECT 3.305 2.230 3.315 2.530 ;
        RECT 3.315 2.230 3.325 2.540 ;
        RECT 3.325 2.230 3.335 2.550 ;
        RECT 3.335 2.230 3.345 2.560 ;
        RECT 3.345 2.230 3.355 2.570 ;
        RECT 3.355 2.230 3.361 2.580 ;
        RECT 12.385 1.395 12.555 2.215 ;
        RECT 12.255 2.045 12.555 2.215 ;
        RECT 12.595 1.125 12.765 1.565 ;
        RECT 11.655 1.395 12.765 1.565 ;
        RECT 12.595 1.125 13.075 1.295 ;
        RECT 6.425 1.495 7.155 1.665 ;
        RECT 8.210 0.615 8.380 1.315 ;
        RECT 7.580 1.145 8.380 1.315 ;
        RECT 8.210 0.615 9.860 0.785 ;
        RECT 10.070 0.480 10.820 0.650 ;
        RECT 10.885 0.480 10.895 0.715 ;
        RECT 10.960 0.545 11.565 0.715 ;
        RECT 11.395 0.545 11.565 1.140 ;
        RECT 12.245 0.755 12.415 1.140 ;
        RECT 11.395 0.970 12.415 1.140 ;
        RECT 13.280 0.755 13.450 2.215 ;
        RECT 12.245 0.755 13.985 0.925 ;
        RECT 13.280 2.045 13.985 2.215 ;
        RECT 10.895 0.490 10.905 0.714 ;
        RECT 10.905 0.500 10.915 0.714 ;
        RECT 10.915 0.510 10.925 0.714 ;
        RECT 10.925 0.520 10.935 0.714 ;
        RECT 10.935 0.530 10.945 0.714 ;
        RECT 10.945 0.540 10.955 0.714 ;
        RECT 10.955 0.545 10.961 0.715 ;
        RECT 10.820 0.480 10.830 0.650 ;
        RECT 10.830 0.480 10.840 0.660 ;
        RECT 10.840 0.480 10.850 0.670 ;
        RECT 10.850 0.480 10.860 0.680 ;
        RECT 10.860 0.480 10.870 0.690 ;
        RECT 10.870 0.480 10.880 0.700 ;
        RECT 10.880 0.480 10.886 0.710 ;
        RECT 9.995 0.480 10.005 0.714 ;
        RECT 10.005 0.480 10.015 0.704 ;
        RECT 10.015 0.480 10.025 0.694 ;
        RECT 10.025 0.480 10.035 0.684 ;
        RECT 10.035 0.480 10.045 0.674 ;
        RECT 10.045 0.480 10.055 0.664 ;
        RECT 10.055 0.480 10.065 0.654 ;
        RECT 10.065 0.480 10.071 0.650 ;
        RECT 9.935 0.540 9.945 0.774 ;
        RECT 9.945 0.530 9.955 0.764 ;
        RECT 9.955 0.520 9.965 0.754 ;
        RECT 9.965 0.510 9.975 0.744 ;
        RECT 9.975 0.500 9.985 0.734 ;
        RECT 9.985 0.490 9.995 0.724 ;
        RECT 9.860 0.615 9.870 0.785 ;
        RECT 9.870 0.605 9.880 0.785 ;
        RECT 9.880 0.595 9.890 0.785 ;
        RECT 9.890 0.585 9.900 0.785 ;
        RECT 9.900 0.575 9.910 0.785 ;
        RECT 9.910 0.565 9.920 0.785 ;
        RECT 9.920 0.555 9.930 0.785 ;
        RECT 9.930 0.545 9.936 0.785 ;
        RECT 7.505 1.145 7.515 1.379 ;
        RECT 7.515 1.145 7.525 1.369 ;
        RECT 7.525 1.145 7.535 1.359 ;
        RECT 7.535 1.145 7.545 1.349 ;
        RECT 7.545 1.145 7.555 1.339 ;
        RECT 7.555 1.145 7.565 1.329 ;
        RECT 7.565 1.145 7.575 1.319 ;
        RECT 7.575 1.145 7.581 1.315 ;
        RECT 7.230 1.420 7.240 1.654 ;
        RECT 7.240 1.410 7.250 1.644 ;
        RECT 7.250 1.400 7.260 1.634 ;
        RECT 7.260 1.390 7.270 1.624 ;
        RECT 7.270 1.380 7.280 1.614 ;
        RECT 7.280 1.370 7.290 1.604 ;
        RECT 7.290 1.360 7.300 1.594 ;
        RECT 7.300 1.350 7.310 1.584 ;
        RECT 7.310 1.340 7.320 1.574 ;
        RECT 7.320 1.330 7.330 1.564 ;
        RECT 7.330 1.320 7.340 1.554 ;
        RECT 7.340 1.310 7.350 1.544 ;
        RECT 7.350 1.300 7.360 1.534 ;
        RECT 7.360 1.290 7.370 1.524 ;
        RECT 7.370 1.280 7.380 1.514 ;
        RECT 7.380 1.270 7.390 1.504 ;
        RECT 7.390 1.260 7.400 1.494 ;
        RECT 7.400 1.250 7.410 1.484 ;
        RECT 7.410 1.240 7.420 1.474 ;
        RECT 7.420 1.230 7.430 1.464 ;
        RECT 7.430 1.220 7.440 1.454 ;
        RECT 7.440 1.210 7.450 1.444 ;
        RECT 7.450 1.200 7.460 1.434 ;
        RECT 7.460 1.190 7.470 1.424 ;
        RECT 7.470 1.180 7.480 1.414 ;
        RECT 7.480 1.170 7.490 1.404 ;
        RECT 7.490 1.160 7.500 1.394 ;
        RECT 7.500 1.150 7.506 1.390 ;
        RECT 7.155 1.495 7.165 1.665 ;
        RECT 7.165 1.485 7.175 1.665 ;
        RECT 7.175 1.475 7.185 1.665 ;
        RECT 7.185 1.465 7.195 1.665 ;
        RECT 7.195 1.455 7.205 1.665 ;
        RECT 7.205 1.445 7.215 1.665 ;
        RECT 7.215 1.435 7.225 1.665 ;
        RECT 7.225 1.425 7.231 1.665 ;
        RECT 9.745 0.965 10.010 1.135 ;
        RECT 9.915 2.545 10.085 2.855 ;
        RECT 9.745 2.545 10.085 2.715 ;
        RECT 10.220 0.830 10.670 1.000 ;
        RECT 10.815 0.895 11.035 1.415 ;
        RECT 10.835 2.465 11.135 2.855 ;
        RECT 9.915 2.685 11.135 2.855 ;
        RECT 11.110 0.895 11.145 1.490 ;
        RECT 11.235 1.320 11.295 1.490 ;
        RECT 10.835 2.465 11.545 2.645 ;
        RECT 12.485 2.465 12.785 2.705 ;
        RECT 14.375 1.585 14.555 2.645 ;
        RECT 11.715 2.465 14.555 2.645 ;
        RECT 14.375 1.585 15.215 1.755 ;
        RECT 11.545 1.805 11.555 2.645 ;
        RECT 11.555 1.815 11.565 2.645 ;
        RECT 11.565 1.825 11.575 2.645 ;
        RECT 11.575 1.835 11.585 2.645 ;
        RECT 11.585 1.845 11.595 2.645 ;
        RECT 11.595 1.855 11.605 2.645 ;
        RECT 11.605 1.865 11.615 2.645 ;
        RECT 11.615 1.875 11.625 2.645 ;
        RECT 11.625 1.885 11.635 2.645 ;
        RECT 11.635 1.895 11.645 2.645 ;
        RECT 11.645 1.905 11.655 2.645 ;
        RECT 11.655 1.915 11.665 2.645 ;
        RECT 11.665 1.925 11.675 2.645 ;
        RECT 11.675 1.935 11.685 2.645 ;
        RECT 11.685 1.945 11.695 2.645 ;
        RECT 11.695 1.955 11.705 2.645 ;
        RECT 11.705 1.965 11.715 2.645 ;
        RECT 11.465 1.725 11.475 1.959 ;
        RECT 11.475 1.735 11.485 1.969 ;
        RECT 11.485 1.745 11.495 1.979 ;
        RECT 11.495 1.755 11.505 1.989 ;
        RECT 11.505 1.765 11.515 1.999 ;
        RECT 11.515 1.775 11.525 2.009 ;
        RECT 11.525 1.785 11.535 2.019 ;
        RECT 11.535 1.795 11.545 2.029 ;
        RECT 11.295 1.320 11.305 1.790 ;
        RECT 11.305 1.320 11.315 1.800 ;
        RECT 11.315 1.320 11.325 1.810 ;
        RECT 11.325 1.320 11.335 1.820 ;
        RECT 11.335 1.320 11.345 1.830 ;
        RECT 11.345 1.320 11.355 1.840 ;
        RECT 11.355 1.320 11.365 1.850 ;
        RECT 11.365 1.320 11.375 1.860 ;
        RECT 11.375 1.320 11.385 1.870 ;
        RECT 11.385 1.320 11.395 1.880 ;
        RECT 11.395 1.320 11.405 1.890 ;
        RECT 11.405 1.320 11.415 1.900 ;
        RECT 11.415 1.320 11.425 1.910 ;
        RECT 11.425 1.320 11.435 1.920 ;
        RECT 11.435 1.320 11.445 1.930 ;
        RECT 11.445 1.320 11.455 1.940 ;
        RECT 11.455 1.320 11.465 1.950 ;
        RECT 11.145 1.240 11.155 1.490 ;
        RECT 11.155 1.250 11.165 1.490 ;
        RECT 11.165 1.260 11.175 1.490 ;
        RECT 11.175 1.270 11.185 1.490 ;
        RECT 11.185 1.280 11.195 1.490 ;
        RECT 11.195 1.290 11.205 1.490 ;
        RECT 11.205 1.300 11.215 1.490 ;
        RECT 11.215 1.310 11.225 1.490 ;
        RECT 11.225 1.320 11.235 1.490 ;
        RECT 11.035 0.895 11.045 1.415 ;
        RECT 11.045 0.895 11.055 1.425 ;
        RECT 11.055 0.895 11.065 1.435 ;
        RECT 11.065 0.895 11.075 1.445 ;
        RECT 11.075 0.895 11.085 1.455 ;
        RECT 11.085 0.895 11.095 1.465 ;
        RECT 11.095 0.895 11.105 1.475 ;
        RECT 11.105 0.895 11.111 1.485 ;
        RECT 10.810 0.895 10.816 1.139 ;
        RECT 10.745 0.840 10.755 1.074 ;
        RECT 10.755 0.850 10.765 1.084 ;
        RECT 10.765 0.860 10.775 1.094 ;
        RECT 10.775 0.870 10.785 1.104 ;
        RECT 10.785 0.880 10.795 1.114 ;
        RECT 10.795 0.890 10.805 1.124 ;
        RECT 10.805 0.895 10.811 1.135 ;
        RECT 10.670 0.830 10.680 1.000 ;
        RECT 10.680 0.830 10.690 1.010 ;
        RECT 10.690 0.830 10.700 1.020 ;
        RECT 10.700 0.830 10.710 1.030 ;
        RECT 10.710 0.830 10.720 1.040 ;
        RECT 10.720 0.830 10.730 1.050 ;
        RECT 10.730 0.830 10.740 1.060 ;
        RECT 10.740 0.830 10.746 1.070 ;
        RECT 10.145 0.830 10.155 1.064 ;
        RECT 10.155 0.830 10.165 1.054 ;
        RECT 10.165 0.830 10.175 1.044 ;
        RECT 10.175 0.830 10.185 1.034 ;
        RECT 10.185 0.830 10.195 1.024 ;
        RECT 10.195 0.830 10.205 1.014 ;
        RECT 10.205 0.830 10.215 1.004 ;
        RECT 10.215 0.830 10.221 1.000 ;
        RECT 10.085 0.890 10.095 1.124 ;
        RECT 10.095 0.880 10.105 1.114 ;
        RECT 10.105 0.870 10.115 1.104 ;
        RECT 10.115 0.860 10.125 1.094 ;
        RECT 10.125 0.850 10.135 1.084 ;
        RECT 10.135 0.840 10.145 1.074 ;
        RECT 10.010 0.965 10.020 1.135 ;
        RECT 10.020 0.955 10.030 1.135 ;
        RECT 10.030 0.945 10.040 1.135 ;
        RECT 10.040 0.935 10.050 1.135 ;
        RECT 10.050 0.925 10.060 1.135 ;
        RECT 10.060 0.915 10.070 1.135 ;
        RECT 10.070 0.905 10.080 1.135 ;
        RECT 10.080 0.895 10.086 1.135 ;
  END 
END FFDSRHQHD3XHT

MACRO FFDSRHQHD2XHT
  CLASS  CORE ;
  FOREIGN FFDSRHQHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.760 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.710 0.720 13.935 2.960 ;
        RECT 13.710 1.610 14.250 2.095 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.495 2.560 2.050 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 12.620 1.260 13.130 1.785 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.995 ;
        RECT 2.175 -0.300 2.475 1.230 ;
        RECT 4.035 -0.300 4.335 0.990 ;
        RECT 7.115 -0.300 7.415 0.435 ;
        RECT 8.215 -0.300 8.515 0.435 ;
        RECT 10.645 -0.300 10.945 0.715 ;
        RECT 13.125 -0.300 13.425 1.055 ;
        RECT 14.165 -0.300 14.465 1.055 ;
        RECT 0.000 -0.300 14.760 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.870 1.260 1.130 1.795 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 11.125 2.905 11.860 3.185 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 1.980 0.340 3.990 ;
        RECT 2.145 3.215 2.445 3.990 ;
        RECT 3.915 3.095 4.215 3.990 ;
        RECT 5.980 3.235 6.280 3.990 ;
        RECT 6.825 3.025 7.125 3.990 ;
        RECT 7.825 3.025 8.125 3.990 ;
        RECT 10.645 2.845 10.945 3.990 ;
        RECT 12.055 2.885 12.355 3.990 ;
        RECT 13.125 2.975 13.425 3.990 ;
        RECT 14.165 2.295 14.465 3.990 ;
        RECT 0.000 3.390 14.760 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.000 1.975 1.170 2.215 ;
        RECT 0.870 2.045 1.170 2.215 ;
        RECT 1.145 0.825 1.480 0.995 ;
        RECT 1.000 1.975 1.480 2.145 ;
        RECT 1.310 0.825 1.480 2.145 ;
        RECT 1.310 1.610 1.540 1.910 ;
        RECT 3.115 2.165 3.285 2.335 ;
        RECT 3.130 0.995 3.300 1.495 ;
        RECT 3.130 1.325 3.415 1.495 ;
        RECT 3.315 1.325 3.415 2.335 ;
        RECT 3.485 1.325 4.150 1.495 ;
        RECT 4.490 1.675 5.045 1.845 ;
        RECT 4.320 1.430 4.330 1.844 ;
        RECT 4.330 1.440 4.340 1.844 ;
        RECT 4.340 1.450 4.350 1.844 ;
        RECT 4.350 1.460 4.360 1.844 ;
        RECT 4.360 1.470 4.370 1.844 ;
        RECT 4.370 1.480 4.380 1.844 ;
        RECT 4.380 1.490 4.390 1.844 ;
        RECT 4.390 1.500 4.400 1.844 ;
        RECT 4.400 1.510 4.410 1.844 ;
        RECT 4.410 1.520 4.420 1.844 ;
        RECT 4.420 1.530 4.430 1.844 ;
        RECT 4.430 1.540 4.440 1.844 ;
        RECT 4.440 1.550 4.450 1.844 ;
        RECT 4.450 1.560 4.460 1.844 ;
        RECT 4.460 1.570 4.470 1.844 ;
        RECT 4.470 1.580 4.480 1.844 ;
        RECT 4.480 1.590 4.490 1.844 ;
        RECT 4.225 1.335 4.235 1.569 ;
        RECT 4.235 1.345 4.245 1.579 ;
        RECT 4.245 1.355 4.255 1.589 ;
        RECT 4.255 1.365 4.265 1.599 ;
        RECT 4.265 1.375 4.275 1.609 ;
        RECT 4.275 1.385 4.285 1.619 ;
        RECT 4.285 1.395 4.295 1.629 ;
        RECT 4.295 1.405 4.305 1.639 ;
        RECT 4.305 1.415 4.315 1.649 ;
        RECT 4.315 1.420 4.321 1.660 ;
        RECT 4.150 1.325 4.160 1.495 ;
        RECT 4.160 1.325 4.170 1.505 ;
        RECT 4.170 1.325 4.180 1.515 ;
        RECT 4.180 1.325 4.190 1.525 ;
        RECT 4.190 1.325 4.200 1.535 ;
        RECT 4.200 1.325 4.210 1.545 ;
        RECT 4.210 1.325 4.220 1.555 ;
        RECT 4.220 1.325 4.226 1.565 ;
        RECT 3.415 1.325 3.425 2.325 ;
        RECT 3.425 1.325 3.435 2.315 ;
        RECT 3.435 1.325 3.445 2.305 ;
        RECT 3.445 1.325 3.455 2.295 ;
        RECT 3.455 1.325 3.465 2.285 ;
        RECT 3.465 1.325 3.475 2.275 ;
        RECT 3.475 1.325 3.485 2.265 ;
        RECT 3.285 2.165 3.295 2.335 ;
        RECT 3.295 2.155 3.305 2.335 ;
        RECT 3.305 2.145 3.315 2.335 ;
        RECT 4.455 1.125 4.645 1.295 ;
        RECT 4.965 1.325 5.120 1.495 ;
        RECT 5.550 1.675 5.895 1.845 ;
        RECT 5.470 1.605 5.480 1.845 ;
        RECT 5.480 1.615 5.490 1.845 ;
        RECT 5.490 1.625 5.500 1.845 ;
        RECT 5.500 1.635 5.510 1.845 ;
        RECT 5.510 1.645 5.520 1.845 ;
        RECT 5.520 1.655 5.530 1.845 ;
        RECT 5.530 1.665 5.540 1.845 ;
        RECT 5.540 1.675 5.550 1.845 ;
        RECT 5.200 1.335 5.210 1.575 ;
        RECT 5.210 1.345 5.220 1.585 ;
        RECT 5.220 1.355 5.230 1.595 ;
        RECT 5.230 1.365 5.240 1.605 ;
        RECT 5.240 1.375 5.250 1.615 ;
        RECT 5.250 1.385 5.260 1.625 ;
        RECT 5.260 1.395 5.270 1.635 ;
        RECT 5.270 1.405 5.280 1.645 ;
        RECT 5.280 1.415 5.290 1.655 ;
        RECT 5.290 1.425 5.300 1.665 ;
        RECT 5.300 1.435 5.310 1.675 ;
        RECT 5.310 1.445 5.320 1.685 ;
        RECT 5.320 1.455 5.330 1.695 ;
        RECT 5.330 1.465 5.340 1.705 ;
        RECT 5.340 1.475 5.350 1.715 ;
        RECT 5.350 1.485 5.360 1.725 ;
        RECT 5.360 1.495 5.370 1.735 ;
        RECT 5.370 1.505 5.380 1.745 ;
        RECT 5.380 1.515 5.390 1.755 ;
        RECT 5.390 1.525 5.400 1.765 ;
        RECT 5.400 1.535 5.410 1.775 ;
        RECT 5.410 1.545 5.420 1.785 ;
        RECT 5.420 1.555 5.430 1.795 ;
        RECT 5.430 1.565 5.440 1.805 ;
        RECT 5.440 1.575 5.450 1.815 ;
        RECT 5.450 1.585 5.460 1.825 ;
        RECT 5.460 1.595 5.470 1.835 ;
        RECT 5.120 1.325 5.130 1.495 ;
        RECT 5.130 1.325 5.140 1.505 ;
        RECT 5.140 1.325 5.150 1.515 ;
        RECT 5.150 1.325 5.160 1.525 ;
        RECT 5.160 1.325 5.170 1.535 ;
        RECT 5.170 1.325 5.180 1.545 ;
        RECT 5.180 1.325 5.190 1.555 ;
        RECT 5.190 1.325 5.200 1.565 ;
        RECT 4.845 1.215 4.855 1.495 ;
        RECT 4.855 1.225 4.865 1.495 ;
        RECT 4.865 1.235 4.875 1.495 ;
        RECT 4.875 1.245 4.885 1.495 ;
        RECT 4.885 1.255 4.895 1.495 ;
        RECT 4.895 1.265 4.905 1.495 ;
        RECT 4.905 1.275 4.915 1.495 ;
        RECT 4.915 1.285 4.925 1.495 ;
        RECT 4.925 1.295 4.935 1.495 ;
        RECT 4.935 1.305 4.945 1.495 ;
        RECT 4.945 1.315 4.955 1.495 ;
        RECT 4.955 1.325 4.965 1.495 ;
        RECT 4.765 1.135 4.775 1.415 ;
        RECT 4.775 1.145 4.785 1.425 ;
        RECT 4.785 1.155 4.795 1.435 ;
        RECT 4.795 1.165 4.805 1.445 ;
        RECT 4.805 1.175 4.815 1.455 ;
        RECT 4.815 1.185 4.825 1.465 ;
        RECT 4.825 1.195 4.835 1.475 ;
        RECT 4.835 1.205 4.845 1.485 ;
        RECT 4.645 1.125 4.655 1.295 ;
        RECT 4.655 1.125 4.665 1.305 ;
        RECT 4.665 1.125 4.675 1.315 ;
        RECT 4.675 1.125 4.685 1.325 ;
        RECT 4.685 1.125 4.695 1.335 ;
        RECT 4.695 1.125 4.705 1.345 ;
        RECT 4.705 1.125 4.715 1.355 ;
        RECT 4.715 1.125 4.725 1.365 ;
        RECT 4.725 1.125 4.735 1.375 ;
        RECT 4.735 1.125 4.745 1.385 ;
        RECT 4.745 1.125 4.755 1.395 ;
        RECT 4.755 1.125 4.765 1.405 ;
        RECT 4.735 0.540 5.035 0.775 ;
        RECT 4.735 0.540 6.075 0.710 ;
        RECT 5.775 0.540 6.075 1.145 ;
        RECT 5.775 0.975 6.805 1.145 ;
        RECT 6.505 0.975 6.805 1.295 ;
        RECT 3.775 1.675 4.075 2.215 ;
        RECT 6.085 1.325 6.255 2.215 ;
        RECT 5.700 1.325 6.255 1.495 ;
        RECT 6.085 1.495 6.325 2.215 ;
        RECT 3.770 2.045 6.325 2.215 ;
        RECT 6.085 1.495 7.835 1.665 ;
        RECT 5.625 1.260 5.635 1.494 ;
        RECT 5.635 1.270 5.645 1.494 ;
        RECT 5.645 1.280 5.655 1.494 ;
        RECT 5.655 1.290 5.665 1.494 ;
        RECT 5.665 1.300 5.675 1.494 ;
        RECT 5.675 1.310 5.685 1.494 ;
        RECT 5.685 1.320 5.695 1.494 ;
        RECT 5.695 1.325 5.701 1.495 ;
        RECT 5.490 1.125 5.500 1.359 ;
        RECT 5.500 1.135 5.510 1.369 ;
        RECT 5.510 1.145 5.520 1.379 ;
        RECT 5.520 1.155 5.530 1.389 ;
        RECT 5.530 1.165 5.540 1.399 ;
        RECT 5.540 1.175 5.550 1.409 ;
        RECT 5.550 1.185 5.560 1.419 ;
        RECT 5.560 1.195 5.570 1.429 ;
        RECT 5.570 1.205 5.580 1.439 ;
        RECT 5.580 1.215 5.590 1.449 ;
        RECT 5.590 1.225 5.600 1.459 ;
        RECT 5.600 1.235 5.610 1.469 ;
        RECT 5.610 1.245 5.620 1.479 ;
        RECT 5.620 1.250 5.626 1.490 ;
        RECT 5.320 0.890 5.330 1.190 ;
        RECT 5.330 0.890 5.340 1.200 ;
        RECT 5.340 0.890 5.350 1.210 ;
        RECT 5.350 0.890 5.360 1.220 ;
        RECT 5.360 0.890 5.370 1.230 ;
        RECT 5.370 0.890 5.380 1.240 ;
        RECT 5.380 0.890 5.390 1.250 ;
        RECT 5.390 0.890 5.400 1.260 ;
        RECT 5.400 0.890 5.410 1.270 ;
        RECT 5.410 0.890 5.420 1.280 ;
        RECT 5.420 0.890 5.430 1.290 ;
        RECT 5.430 0.890 5.440 1.300 ;
        RECT 5.440 0.890 5.450 1.310 ;
        RECT 5.450 0.890 5.460 1.320 ;
        RECT 5.460 0.890 5.470 1.330 ;
        RECT 5.470 0.890 5.480 1.340 ;
        RECT 5.480 0.890 5.490 1.350 ;
        RECT 0.170 0.720 0.340 1.790 ;
        RECT 0.170 1.620 0.690 1.790 ;
        RECT 0.520 1.620 0.690 2.665 ;
        RECT 0.520 2.495 1.230 2.665 ;
        RECT 1.060 2.495 1.230 3.035 ;
        RECT 1.060 2.865 3.640 3.035 ;
        RECT 3.835 2.745 6.560 2.915 ;
        RECT 6.630 2.675 6.645 2.915 ;
        RECT 6.715 2.675 8.200 2.845 ;
        RECT 8.450 2.850 8.655 3.085 ;
        RECT 8.355 2.765 8.365 3.085 ;
        RECT 8.365 2.775 8.375 3.085 ;
        RECT 8.375 2.785 8.385 3.085 ;
        RECT 8.385 2.795 8.395 3.085 ;
        RECT 8.395 2.805 8.405 3.085 ;
        RECT 8.405 2.815 8.415 3.085 ;
        RECT 8.415 2.825 8.425 3.085 ;
        RECT 8.425 2.835 8.435 3.085 ;
        RECT 8.435 2.845 8.445 3.085 ;
        RECT 8.445 2.850 8.451 3.084 ;
        RECT 8.275 2.685 8.285 2.919 ;
        RECT 8.285 2.695 8.295 2.929 ;
        RECT 8.295 2.705 8.305 2.939 ;
        RECT 8.305 2.715 8.315 2.949 ;
        RECT 8.315 2.725 8.325 2.959 ;
        RECT 8.325 2.735 8.335 2.969 ;
        RECT 8.335 2.745 8.345 2.979 ;
        RECT 8.345 2.755 8.355 2.989 ;
        RECT 8.200 2.675 8.210 2.845 ;
        RECT 8.210 2.675 8.220 2.855 ;
        RECT 8.220 2.675 8.230 2.865 ;
        RECT 8.230 2.675 8.240 2.875 ;
        RECT 8.240 2.675 8.250 2.885 ;
        RECT 8.250 2.675 8.260 2.895 ;
        RECT 8.260 2.675 8.270 2.905 ;
        RECT 8.270 2.675 8.276 2.915 ;
        RECT 6.645 2.675 6.655 2.905 ;
        RECT 6.655 2.675 6.665 2.895 ;
        RECT 6.665 2.675 6.675 2.885 ;
        RECT 6.675 2.675 6.685 2.875 ;
        RECT 6.685 2.675 6.695 2.865 ;
        RECT 6.695 2.675 6.705 2.855 ;
        RECT 6.705 2.675 6.715 2.845 ;
        RECT 6.560 2.745 6.570 2.915 ;
        RECT 6.570 2.735 6.580 2.915 ;
        RECT 6.580 2.725 6.590 2.915 ;
        RECT 6.590 2.715 6.600 2.915 ;
        RECT 6.600 2.705 6.610 2.915 ;
        RECT 6.610 2.695 6.620 2.915 ;
        RECT 6.620 2.685 6.630 2.915 ;
        RECT 3.760 2.745 3.770 2.979 ;
        RECT 3.770 2.745 3.780 2.969 ;
        RECT 3.780 2.745 3.790 2.959 ;
        RECT 3.790 2.745 3.800 2.949 ;
        RECT 3.800 2.745 3.810 2.939 ;
        RECT 3.810 2.745 3.820 2.929 ;
        RECT 3.820 2.745 3.830 2.919 ;
        RECT 3.830 2.745 3.836 2.915 ;
        RECT 3.715 2.790 3.725 3.024 ;
        RECT 3.725 2.780 3.735 3.014 ;
        RECT 3.735 2.770 3.745 3.004 ;
        RECT 3.745 2.760 3.755 2.994 ;
        RECT 3.755 2.750 3.761 2.990 ;
        RECT 3.640 2.865 3.650 3.035 ;
        RECT 3.650 2.855 3.660 3.035 ;
        RECT 3.660 2.845 3.670 3.035 ;
        RECT 3.670 2.835 3.680 3.035 ;
        RECT 3.680 2.825 3.690 3.035 ;
        RECT 3.690 2.815 3.700 3.035 ;
        RECT 3.700 2.805 3.710 3.035 ;
        RECT 3.710 2.795 3.716 3.035 ;
        RECT 7.375 2.210 8.235 2.380 ;
        RECT 8.555 2.455 9.390 2.625 ;
        RECT 9.220 2.455 9.390 2.755 ;
        RECT 8.480 2.390 8.490 2.624 ;
        RECT 8.490 2.400 8.500 2.624 ;
        RECT 8.500 2.410 8.510 2.624 ;
        RECT 8.510 2.420 8.520 2.624 ;
        RECT 8.520 2.430 8.530 2.624 ;
        RECT 8.530 2.440 8.540 2.624 ;
        RECT 8.540 2.450 8.550 2.624 ;
        RECT 8.550 2.455 8.556 2.625 ;
        RECT 8.310 2.220 8.320 2.454 ;
        RECT 8.320 2.230 8.330 2.464 ;
        RECT 8.330 2.240 8.340 2.474 ;
        RECT 8.340 2.250 8.350 2.484 ;
        RECT 8.350 2.260 8.360 2.494 ;
        RECT 8.360 2.270 8.370 2.504 ;
        RECT 8.370 2.280 8.380 2.514 ;
        RECT 8.380 2.290 8.390 2.524 ;
        RECT 8.390 2.300 8.400 2.534 ;
        RECT 8.400 2.310 8.410 2.544 ;
        RECT 8.410 2.320 8.420 2.554 ;
        RECT 8.420 2.330 8.430 2.564 ;
        RECT 8.430 2.340 8.440 2.574 ;
        RECT 8.440 2.350 8.450 2.584 ;
        RECT 8.450 2.360 8.460 2.594 ;
        RECT 8.460 2.370 8.470 2.604 ;
        RECT 8.470 2.380 8.480 2.614 ;
        RECT 8.235 2.210 8.245 2.380 ;
        RECT 8.245 2.210 8.255 2.390 ;
        RECT 8.255 2.210 8.265 2.400 ;
        RECT 8.265 2.210 8.275 2.410 ;
        RECT 8.275 2.210 8.285 2.420 ;
        RECT 8.285 2.210 8.295 2.430 ;
        RECT 8.295 2.210 8.305 2.440 ;
        RECT 8.305 2.210 8.311 2.450 ;
        RECT 7.665 1.125 8.405 1.295 ;
        RECT 8.235 1.125 8.405 1.485 ;
        RECT 9.155 1.180 9.455 1.485 ;
        RECT 8.235 1.315 9.455 1.485 ;
        RECT 1.720 0.995 1.890 2.685 ;
        RECT 1.440 2.350 1.890 2.685 ;
        RECT 2.765 0.525 2.935 2.685 ;
        RECT 2.765 1.795 3.135 1.965 ;
        RECT 1.440 2.515 3.490 2.685 ;
        RECT 2.765 0.525 3.595 0.695 ;
        RECT 3.685 2.395 6.405 2.565 ;
        RECT 6.475 2.325 6.480 2.565 ;
        RECT 7.025 1.845 7.195 2.495 ;
        RECT 6.550 2.325 7.195 2.495 ;
        RECT 8.045 1.675 8.215 2.015 ;
        RECT 7.025 1.845 8.215 2.015 ;
        RECT 8.045 1.675 9.610 1.845 ;
        RECT 10.195 2.115 10.255 2.285 ;
        RECT 9.955 1.885 9.965 2.285 ;
        RECT 9.965 1.895 9.975 2.285 ;
        RECT 9.975 1.905 9.985 2.285 ;
        RECT 9.985 1.915 9.995 2.285 ;
        RECT 9.995 1.925 10.005 2.285 ;
        RECT 10.005 1.935 10.015 2.285 ;
        RECT 10.015 1.945 10.025 2.285 ;
        RECT 10.025 1.955 10.035 2.285 ;
        RECT 10.035 1.965 10.045 2.285 ;
        RECT 10.045 1.975 10.055 2.285 ;
        RECT 10.055 1.985 10.065 2.285 ;
        RECT 10.065 1.995 10.075 2.285 ;
        RECT 10.075 2.005 10.085 2.285 ;
        RECT 10.085 2.015 10.095 2.285 ;
        RECT 10.095 2.025 10.105 2.285 ;
        RECT 10.105 2.035 10.115 2.285 ;
        RECT 10.115 2.045 10.125 2.285 ;
        RECT 10.125 2.055 10.135 2.285 ;
        RECT 10.135 2.065 10.145 2.285 ;
        RECT 10.145 2.075 10.155 2.285 ;
        RECT 10.155 2.085 10.165 2.285 ;
        RECT 10.165 2.095 10.175 2.285 ;
        RECT 10.175 2.105 10.185 2.285 ;
        RECT 10.185 2.115 10.195 2.285 ;
        RECT 9.755 1.685 9.765 1.989 ;
        RECT 9.765 1.695 9.775 1.999 ;
        RECT 9.775 1.705 9.785 2.009 ;
        RECT 9.785 1.715 9.795 2.019 ;
        RECT 9.795 1.725 9.805 2.029 ;
        RECT 9.805 1.735 9.815 2.039 ;
        RECT 9.815 1.745 9.825 2.049 ;
        RECT 9.825 1.755 9.835 2.059 ;
        RECT 9.835 1.765 9.845 2.069 ;
        RECT 9.845 1.775 9.855 2.079 ;
        RECT 9.855 1.785 9.865 2.089 ;
        RECT 9.865 1.795 9.875 2.099 ;
        RECT 9.875 1.805 9.885 2.109 ;
        RECT 9.885 1.815 9.895 2.119 ;
        RECT 9.895 1.825 9.905 2.129 ;
        RECT 9.905 1.835 9.915 2.139 ;
        RECT 9.915 1.845 9.925 2.149 ;
        RECT 9.925 1.855 9.935 2.159 ;
        RECT 9.935 1.865 9.945 2.169 ;
        RECT 9.945 1.875 9.955 2.179 ;
        RECT 9.610 1.675 9.620 1.845 ;
        RECT 9.620 1.675 9.630 1.855 ;
        RECT 9.630 1.675 9.640 1.865 ;
        RECT 9.640 1.675 9.650 1.875 ;
        RECT 9.650 1.675 9.660 1.885 ;
        RECT 9.660 1.675 9.670 1.895 ;
        RECT 9.670 1.675 9.680 1.905 ;
        RECT 9.680 1.675 9.690 1.915 ;
        RECT 9.690 1.675 9.700 1.925 ;
        RECT 9.700 1.675 9.710 1.935 ;
        RECT 9.710 1.675 9.720 1.945 ;
        RECT 9.720 1.675 9.730 1.955 ;
        RECT 9.730 1.675 9.740 1.965 ;
        RECT 9.740 1.675 9.750 1.975 ;
        RECT 9.750 1.675 9.756 1.985 ;
        RECT 6.480 2.325 6.490 2.555 ;
        RECT 6.490 2.325 6.500 2.545 ;
        RECT 6.500 2.325 6.510 2.535 ;
        RECT 6.510 2.325 6.520 2.525 ;
        RECT 6.520 2.325 6.530 2.515 ;
        RECT 6.530 2.325 6.540 2.505 ;
        RECT 6.540 2.325 6.550 2.495 ;
        RECT 6.405 2.395 6.415 2.565 ;
        RECT 6.415 2.385 6.425 2.565 ;
        RECT 6.425 2.375 6.435 2.565 ;
        RECT 6.435 2.365 6.445 2.565 ;
        RECT 6.445 2.355 6.455 2.565 ;
        RECT 6.455 2.345 6.465 2.565 ;
        RECT 6.465 2.335 6.475 2.565 ;
        RECT 3.610 2.395 3.620 2.629 ;
        RECT 3.620 2.395 3.630 2.619 ;
        RECT 3.630 2.395 3.640 2.609 ;
        RECT 3.640 2.395 3.650 2.599 ;
        RECT 3.650 2.395 3.660 2.589 ;
        RECT 3.660 2.395 3.670 2.579 ;
        RECT 3.670 2.395 3.680 2.569 ;
        RECT 3.680 2.395 3.686 2.565 ;
        RECT 3.565 2.440 3.575 2.674 ;
        RECT 3.575 2.430 3.585 2.664 ;
        RECT 3.585 2.420 3.595 2.654 ;
        RECT 3.595 2.410 3.605 2.644 ;
        RECT 3.605 2.400 3.611 2.640 ;
        RECT 3.490 2.515 3.500 2.685 ;
        RECT 3.500 2.505 3.510 2.685 ;
        RECT 3.510 2.495 3.520 2.685 ;
        RECT 3.520 2.485 3.530 2.685 ;
        RECT 3.530 2.475 3.540 2.685 ;
        RECT 3.540 2.465 3.550 2.685 ;
        RECT 3.550 2.455 3.560 2.685 ;
        RECT 3.560 2.445 3.566 2.685 ;
        RECT 11.265 1.400 11.435 2.215 ;
        RECT 11.135 2.045 11.435 2.215 ;
        RECT 11.475 1.125 11.645 1.570 ;
        RECT 10.535 1.400 11.645 1.570 ;
        RECT 11.475 1.125 11.955 1.295 ;
        RECT 6.255 0.615 8.720 0.785 ;
        RECT 8.930 0.480 9.680 0.650 ;
        RECT 9.745 0.480 9.755 0.715 ;
        RECT 9.820 0.545 10.445 0.715 ;
        RECT 10.275 0.545 10.445 1.140 ;
        RECT 11.125 0.775 11.295 1.140 ;
        RECT 10.275 0.970 11.295 1.140 ;
        RECT 12.135 0.775 12.305 2.215 ;
        RECT 11.125 0.775 12.875 0.945 ;
        RECT 12.135 2.045 12.875 2.215 ;
        RECT 9.755 0.490 9.765 0.714 ;
        RECT 9.765 0.500 9.775 0.714 ;
        RECT 9.775 0.510 9.785 0.714 ;
        RECT 9.785 0.520 9.795 0.714 ;
        RECT 9.795 0.530 9.805 0.714 ;
        RECT 9.805 0.540 9.815 0.714 ;
        RECT 9.815 0.545 9.821 0.715 ;
        RECT 9.680 0.480 9.690 0.650 ;
        RECT 9.690 0.480 9.700 0.660 ;
        RECT 9.700 0.480 9.710 0.670 ;
        RECT 9.710 0.480 9.720 0.680 ;
        RECT 9.720 0.480 9.730 0.690 ;
        RECT 9.730 0.480 9.740 0.700 ;
        RECT 9.740 0.480 9.746 0.710 ;
        RECT 8.855 0.480 8.865 0.714 ;
        RECT 8.865 0.480 8.875 0.704 ;
        RECT 8.875 0.480 8.885 0.694 ;
        RECT 8.885 0.480 8.895 0.684 ;
        RECT 8.895 0.480 8.905 0.674 ;
        RECT 8.905 0.480 8.915 0.664 ;
        RECT 8.915 0.480 8.925 0.654 ;
        RECT 8.925 0.480 8.931 0.650 ;
        RECT 8.795 0.540 8.805 0.774 ;
        RECT 8.805 0.530 8.815 0.764 ;
        RECT 8.815 0.520 8.825 0.754 ;
        RECT 8.825 0.510 8.835 0.744 ;
        RECT 8.835 0.500 8.845 0.734 ;
        RECT 8.845 0.490 8.855 0.724 ;
        RECT 8.720 0.615 8.730 0.785 ;
        RECT 8.730 0.605 8.740 0.785 ;
        RECT 8.740 0.595 8.750 0.785 ;
        RECT 8.750 0.585 8.760 0.785 ;
        RECT 8.760 0.575 8.770 0.785 ;
        RECT 8.770 0.565 8.780 0.785 ;
        RECT 8.780 0.555 8.790 0.785 ;
        RECT 8.790 0.545 8.796 0.785 ;
        RECT 8.605 0.965 8.870 1.135 ;
        RECT 8.635 2.025 8.935 2.275 ;
        RECT 8.635 2.025 9.390 2.195 ;
        RECT 9.080 0.830 9.530 1.000 ;
        RECT 9.595 0.830 9.605 1.065 ;
        RECT 9.670 0.895 9.925 1.065 ;
        RECT 9.705 0.895 9.925 1.415 ;
        RECT 10.000 0.895 10.005 1.490 ;
        RECT 9.775 2.465 10.065 2.675 ;
        RECT 10.125 1.320 10.185 1.490 ;
        RECT 9.775 2.465 10.435 2.635 ;
        RECT 11.365 2.465 11.665 2.705 ;
        RECT 13.360 1.510 13.530 2.635 ;
        RECT 10.605 2.465 13.530 2.635 ;
        RECT 10.435 1.805 10.445 2.635 ;
        RECT 10.445 1.815 10.455 2.635 ;
        RECT 10.455 1.825 10.465 2.635 ;
        RECT 10.465 1.835 10.475 2.635 ;
        RECT 10.475 1.845 10.485 2.635 ;
        RECT 10.485 1.855 10.495 2.635 ;
        RECT 10.495 1.865 10.505 2.635 ;
        RECT 10.505 1.875 10.515 2.635 ;
        RECT 10.515 1.885 10.525 2.635 ;
        RECT 10.525 1.895 10.535 2.635 ;
        RECT 10.535 1.905 10.545 2.635 ;
        RECT 10.545 1.915 10.555 2.635 ;
        RECT 10.555 1.925 10.565 2.635 ;
        RECT 10.565 1.935 10.575 2.635 ;
        RECT 10.575 1.945 10.585 2.635 ;
        RECT 10.585 1.955 10.595 2.635 ;
        RECT 10.595 1.965 10.605 2.635 ;
        RECT 10.355 1.725 10.365 1.959 ;
        RECT 10.365 1.735 10.375 1.969 ;
        RECT 10.375 1.745 10.385 1.979 ;
        RECT 10.385 1.755 10.395 1.989 ;
        RECT 10.395 1.765 10.405 1.999 ;
        RECT 10.405 1.775 10.415 2.009 ;
        RECT 10.415 1.785 10.425 2.019 ;
        RECT 10.425 1.795 10.435 2.029 ;
        RECT 10.185 1.320 10.195 1.790 ;
        RECT 10.195 1.320 10.205 1.800 ;
        RECT 10.205 1.320 10.215 1.810 ;
        RECT 10.215 1.320 10.225 1.820 ;
        RECT 10.225 1.320 10.235 1.830 ;
        RECT 10.235 1.320 10.245 1.840 ;
        RECT 10.245 1.320 10.255 1.850 ;
        RECT 10.255 1.320 10.265 1.860 ;
        RECT 10.265 1.320 10.275 1.870 ;
        RECT 10.275 1.320 10.285 1.880 ;
        RECT 10.285 1.320 10.295 1.890 ;
        RECT 10.295 1.320 10.305 1.900 ;
        RECT 10.305 1.320 10.315 1.910 ;
        RECT 10.315 1.320 10.325 1.920 ;
        RECT 10.325 1.320 10.335 1.930 ;
        RECT 10.335 1.320 10.345 1.940 ;
        RECT 10.345 1.320 10.355 1.950 ;
        RECT 10.005 1.210 10.015 1.490 ;
        RECT 10.015 1.220 10.025 1.490 ;
        RECT 10.025 1.230 10.035 1.490 ;
        RECT 10.035 1.240 10.045 1.490 ;
        RECT 10.045 1.250 10.055 1.490 ;
        RECT 10.055 1.260 10.065 1.490 ;
        RECT 10.065 1.270 10.075 1.490 ;
        RECT 10.075 1.280 10.085 1.490 ;
        RECT 10.085 1.290 10.095 1.490 ;
        RECT 10.095 1.300 10.105 1.490 ;
        RECT 10.105 1.310 10.115 1.490 ;
        RECT 10.115 1.320 10.125 1.490 ;
        RECT 9.925 0.895 9.935 1.415 ;
        RECT 9.935 0.895 9.945 1.425 ;
        RECT 9.945 0.895 9.955 1.435 ;
        RECT 9.955 0.895 9.965 1.445 ;
        RECT 9.965 0.895 9.975 1.455 ;
        RECT 9.975 0.895 9.985 1.465 ;
        RECT 9.985 0.895 9.995 1.475 ;
        RECT 9.995 0.895 10.001 1.485 ;
        RECT 9.605 2.170 9.615 2.674 ;
        RECT 9.615 2.180 9.625 2.674 ;
        RECT 9.625 2.190 9.635 2.674 ;
        RECT 9.635 2.200 9.645 2.674 ;
        RECT 9.645 2.210 9.655 2.674 ;
        RECT 9.655 2.220 9.665 2.674 ;
        RECT 9.665 2.230 9.675 2.674 ;
        RECT 9.675 2.240 9.685 2.674 ;
        RECT 9.685 2.250 9.695 2.674 ;
        RECT 9.695 2.260 9.705 2.674 ;
        RECT 9.705 2.270 9.715 2.674 ;
        RECT 9.715 2.280 9.725 2.674 ;
        RECT 9.725 2.290 9.735 2.674 ;
        RECT 9.735 2.300 9.745 2.674 ;
        RECT 9.745 2.310 9.755 2.674 ;
        RECT 9.755 2.320 9.765 2.674 ;
        RECT 9.765 2.330 9.775 2.674 ;
        RECT 9.605 0.840 9.615 1.064 ;
        RECT 9.615 0.850 9.625 1.064 ;
        RECT 9.625 0.860 9.635 1.064 ;
        RECT 9.635 0.870 9.645 1.064 ;
        RECT 9.645 0.880 9.655 1.064 ;
        RECT 9.655 0.890 9.665 1.064 ;
        RECT 9.665 0.895 9.671 1.065 ;
        RECT 9.470 2.035 9.480 2.275 ;
        RECT 9.480 2.045 9.490 2.285 ;
        RECT 9.490 2.055 9.500 2.295 ;
        RECT 9.500 2.065 9.510 2.305 ;
        RECT 9.510 2.075 9.520 2.315 ;
        RECT 9.520 2.085 9.530 2.325 ;
        RECT 9.530 2.095 9.540 2.335 ;
        RECT 9.540 2.105 9.550 2.345 ;
        RECT 9.550 2.115 9.560 2.355 ;
        RECT 9.560 2.125 9.570 2.365 ;
        RECT 9.570 2.135 9.580 2.375 ;
        RECT 9.580 2.145 9.590 2.385 ;
        RECT 9.590 2.155 9.600 2.395 ;
        RECT 9.600 2.160 9.606 2.404 ;
        RECT 9.530 0.830 9.540 1.000 ;
        RECT 9.540 0.830 9.550 1.010 ;
        RECT 9.550 0.830 9.560 1.020 ;
        RECT 9.560 0.830 9.570 1.030 ;
        RECT 9.570 0.830 9.580 1.040 ;
        RECT 9.580 0.830 9.590 1.050 ;
        RECT 9.590 0.830 9.596 1.060 ;
        RECT 9.390 2.025 9.400 2.195 ;
        RECT 9.400 2.025 9.410 2.205 ;
        RECT 9.410 2.025 9.420 2.215 ;
        RECT 9.420 2.025 9.430 2.225 ;
        RECT 9.430 2.025 9.440 2.235 ;
        RECT 9.440 2.025 9.450 2.245 ;
        RECT 9.450 2.025 9.460 2.255 ;
        RECT 9.460 2.025 9.470 2.265 ;
        RECT 9.005 0.830 9.015 1.064 ;
        RECT 9.015 0.830 9.025 1.054 ;
        RECT 9.025 0.830 9.035 1.044 ;
        RECT 9.035 0.830 9.045 1.034 ;
        RECT 9.045 0.830 9.055 1.024 ;
        RECT 9.055 0.830 9.065 1.014 ;
        RECT 9.065 0.830 9.075 1.004 ;
        RECT 9.075 0.830 9.081 1.000 ;
        RECT 8.945 0.890 8.955 1.124 ;
        RECT 8.955 0.880 8.965 1.114 ;
        RECT 8.965 0.870 8.975 1.104 ;
        RECT 8.975 0.860 8.985 1.094 ;
        RECT 8.985 0.850 8.995 1.084 ;
        RECT 8.995 0.840 9.005 1.074 ;
        RECT 8.870 0.965 8.880 1.135 ;
        RECT 8.880 0.955 8.890 1.135 ;
        RECT 8.890 0.945 8.900 1.135 ;
        RECT 8.900 0.935 8.910 1.135 ;
        RECT 8.910 0.925 8.920 1.135 ;
        RECT 8.920 0.915 8.930 1.135 ;
        RECT 8.930 0.905 8.940 1.135 ;
        RECT 8.940 0.895 8.946 1.135 ;
  END 
END FFDSRHQHD2XHT

MACRO FFDSRHQHD1XHT
  CLASS  CORE ;
  FOREIGN FFDSRHQHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.480 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.760 1.980 11.240 2.430 ;
        RECT 11.005 0.720 11.240 1.360 ;
        RECT 11.030 0.720 11.240 3.210 ;
        RECT 11.005 1.980 11.240 3.210 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.490 2.560 2.050 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 9.940 1.200 10.215 1.735 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.995 ;
        RECT 2.175 -0.300 2.475 1.230 ;
        RECT 3.975 -0.300 4.215 0.580 ;
        RECT 6.160 -0.300 6.330 0.550 ;
        RECT 8.050 -0.300 8.350 0.795 ;
        RECT 10.420 -0.300 10.720 1.055 ;
        RECT 0.000 -0.300 11.480 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.870 1.260 1.130 1.800 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 8.230 1.330 8.755 1.540 ;
        RECT 8.425 1.330 8.755 1.800 ;
        RECT 6.545 2.625 6.621 2.805 ;
        RECT 6.555 2.625 6.621 2.815 ;
        RECT 6.565 2.625 6.621 2.825 ;
        RECT 6.640 3.020 7.826 3.189 ;
        RECT 5.810 2.625 5.980 3.110 ;
        RECT 6.575 2.625 6.621 2.835 ;
        RECT 6.575 2.825 6.820 2.835 ;
        RECT 6.585 2.625 6.621 2.845 ;
        RECT 6.585 2.825 6.820 2.845 ;
        RECT 6.595 2.625 6.621 2.855 ;
        RECT 6.595 2.825 6.820 2.855 ;
        RECT 6.605 2.625 6.621 2.865 ;
        RECT 6.605 2.825 6.820 2.865 ;
        RECT 6.615 2.625 6.621 2.875 ;
        RECT 6.615 2.825 6.820 2.875 ;
        RECT 6.620 2.625 6.621 2.879 ;
        RECT 5.810 2.625 6.621 2.795 ;
        RECT 6.620 2.635 6.630 2.879 ;
        RECT 6.620 2.825 6.820 2.879 ;
        RECT 5.810 2.635 6.630 2.795 ;
        RECT 6.630 2.645 6.640 2.889 ;
        RECT 6.630 2.825 6.820 2.889 ;
        RECT 5.810 2.645 6.640 2.795 ;
        RECT 6.640 2.655 6.650 3.189 ;
        RECT 5.810 2.655 6.650 2.795 ;
        RECT 6.640 2.665 6.660 3.189 ;
        RECT 5.810 2.665 6.660 2.795 ;
        RECT 6.640 2.675 6.670 3.189 ;
        RECT 5.810 2.675 6.670 2.795 ;
        RECT 6.640 2.685 6.680 3.189 ;
        RECT 5.810 2.685 6.680 2.795 ;
        RECT 6.640 2.695 6.690 3.189 ;
        RECT 5.810 2.695 6.690 2.795 ;
        RECT 6.640 2.705 6.700 3.189 ;
        RECT 5.810 2.705 6.700 2.795 ;
        RECT 6.640 2.715 6.710 3.189 ;
        RECT 5.810 2.715 6.710 2.795 ;
        RECT 6.640 2.725 6.720 3.189 ;
        RECT 5.810 2.725 6.720 2.795 ;
        RECT 6.640 2.735 6.730 3.189 ;
        RECT 5.810 2.735 6.730 2.795 ;
        RECT 6.640 2.745 6.740 3.189 ;
        RECT 5.810 2.745 6.740 2.795 ;
        RECT 6.640 2.755 6.750 3.189 ;
        RECT 5.810 2.755 6.750 2.795 ;
        RECT 6.640 2.765 6.760 3.189 ;
        RECT 5.810 2.765 6.760 2.795 ;
        RECT 6.640 2.775 6.770 3.189 ;
        RECT 5.810 2.775 6.770 2.795 ;
        RECT 6.640 2.785 6.780 3.189 ;
        RECT 5.810 2.785 6.780 2.795 ;
        RECT 6.640 2.795 6.790 3.189 ;
        RECT 6.545 2.795 6.790 2.805 ;
        RECT 6.640 2.805 6.800 3.189 ;
        RECT 6.555 2.805 6.800 2.815 ;
        RECT 6.640 2.815 6.810 3.189 ;
        RECT 6.565 2.815 6.810 2.825 ;
        RECT 6.640 2.825 6.820 3.189 ;
        RECT 7.800 2.950 7.826 3.190 ;
        RECT 7.800 2.950 8.830 3.055 ;
        RECT 7.810 2.940 7.826 3.190 ;
        RECT 7.790 2.960 8.830 3.055 ;
        RECT 7.820 2.930 7.826 3.190 ;
        RECT 7.780 2.970 8.830 3.055 ;
        RECT 7.825 2.925 7.826 3.190 ;
        RECT 6.820 3.020 7.826 3.190 ;
        RECT 7.825 2.925 7.835 3.179 ;
        RECT 7.770 2.980 8.830 3.055 ;
        RECT 6.640 3.020 7.835 3.179 ;
        RECT 7.835 2.915 7.845 3.169 ;
        RECT 7.760 2.990 8.830 3.055 ;
        RECT 6.640 3.020 7.845 3.169 ;
        RECT 7.845 2.905 7.855 3.159 ;
        RECT 7.750 3.000 8.830 3.055 ;
        RECT 6.640 3.020 7.855 3.159 ;
        RECT 7.855 2.895 7.865 3.149 ;
        RECT 7.740 3.010 8.830 3.055 ;
        RECT 6.640 3.020 7.865 3.149 ;
        RECT 7.865 2.885 7.875 3.139 ;
        RECT 6.640 3.020 7.875 3.139 ;
        RECT 7.865 2.885 7.885 3.129 ;
        RECT 6.640 3.020 7.885 3.129 ;
        RECT 7.865 2.885 7.895 3.119 ;
        RECT 6.640 3.020 7.895 3.119 ;
        RECT 7.865 2.885 7.905 3.109 ;
        RECT 6.640 3.020 7.905 3.109 ;
        RECT 7.865 2.885 7.915 3.099 ;
        RECT 6.640 3.020 7.915 3.099 ;
        RECT 7.865 2.885 7.925 3.089 ;
        RECT 6.640 3.020 7.925 3.089 ;
        RECT 7.865 2.885 7.935 3.079 ;
        RECT 6.640 3.020 7.935 3.079 ;
        RECT 7.865 2.885 7.945 3.069 ;
        RECT 6.640 3.020 7.945 3.069 ;
        RECT 7.865 2.885 7.955 3.059 ;
        RECT 6.640 3.020 7.955 3.059 ;
        RECT 7.865 2.885 8.830 3.055 ;
        RECT 8.530 2.885 8.830 3.185 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 1.980 0.340 3.990 ;
        RECT 2.205 3.215 2.505 3.990 ;
        RECT 3.915 3.155 4.215 3.990 ;
        RECT 6.160 2.975 6.460 3.990 ;
        RECT 8.050 3.255 8.350 3.990 ;
        RECT 9.480 2.745 9.780 3.990 ;
        RECT 10.420 2.970 10.720 3.990 ;
        RECT 0.000 3.390 11.480 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.000 1.980 1.170 2.215 ;
        RECT 0.870 2.045 1.170 2.215 ;
        RECT 1.145 0.825 1.480 0.995 ;
        RECT 1.000 1.980 1.480 2.150 ;
        RECT 1.310 0.825 1.480 2.150 ;
        RECT 1.310 1.610 1.540 1.910 ;
        RECT 3.115 2.165 3.285 2.335 ;
        RECT 3.130 0.995 3.300 1.495 ;
        RECT 3.130 1.325 3.415 1.495 ;
        RECT 3.315 1.325 3.415 2.335 ;
        RECT 3.485 1.325 4.150 1.495 ;
        RECT 4.425 1.675 5.035 1.845 ;
        RECT 4.255 1.360 4.265 1.844 ;
        RECT 4.265 1.370 4.275 1.844 ;
        RECT 4.275 1.380 4.285 1.844 ;
        RECT 4.285 1.390 4.295 1.844 ;
        RECT 4.295 1.400 4.305 1.844 ;
        RECT 4.305 1.410 4.315 1.844 ;
        RECT 4.315 1.420 4.325 1.844 ;
        RECT 4.325 1.430 4.335 1.844 ;
        RECT 4.335 1.440 4.345 1.844 ;
        RECT 4.345 1.450 4.355 1.844 ;
        RECT 4.355 1.460 4.365 1.844 ;
        RECT 4.365 1.470 4.375 1.844 ;
        RECT 4.375 1.480 4.385 1.844 ;
        RECT 4.385 1.490 4.395 1.844 ;
        RECT 4.395 1.500 4.405 1.844 ;
        RECT 4.405 1.510 4.415 1.844 ;
        RECT 4.415 1.520 4.425 1.844 ;
        RECT 4.230 1.335 4.240 1.575 ;
        RECT 4.240 1.345 4.250 1.585 ;
        RECT 4.250 1.350 4.256 1.594 ;
        RECT 4.150 1.325 4.160 1.495 ;
        RECT 4.160 1.325 4.170 1.505 ;
        RECT 4.170 1.325 4.180 1.515 ;
        RECT 4.180 1.325 4.190 1.525 ;
        RECT 4.190 1.325 4.200 1.535 ;
        RECT 4.200 1.325 4.210 1.545 ;
        RECT 4.210 1.325 4.220 1.555 ;
        RECT 4.220 1.325 4.230 1.565 ;
        RECT 3.415 1.325 3.425 2.325 ;
        RECT 3.425 1.325 3.435 2.315 ;
        RECT 3.435 1.325 3.445 2.305 ;
        RECT 3.445 1.325 3.455 2.295 ;
        RECT 3.455 1.325 3.465 2.285 ;
        RECT 3.465 1.325 3.475 2.275 ;
        RECT 3.475 1.325 3.485 2.265 ;
        RECT 3.285 2.165 3.295 2.335 ;
        RECT 3.295 2.155 3.305 2.335 ;
        RECT 3.305 2.145 3.315 2.335 ;
        RECT 0.170 1.060 0.340 1.790 ;
        RECT 0.170 1.620 0.690 1.790 ;
        RECT 0.520 1.620 0.690 2.565 ;
        RECT 0.520 2.395 1.230 2.565 ;
        RECT 1.060 2.395 1.230 3.035 ;
        RECT 1.060 2.865 3.645 3.035 ;
        RECT 3.705 2.805 3.720 3.035 ;
        RECT 3.780 2.805 4.425 2.975 ;
        RECT 4.750 3.040 5.565 3.210 ;
        RECT 4.660 2.960 4.670 3.210 ;
        RECT 4.670 2.970 4.680 3.210 ;
        RECT 4.680 2.980 4.690 3.210 ;
        RECT 4.690 2.990 4.700 3.210 ;
        RECT 4.700 3.000 4.710 3.210 ;
        RECT 4.710 3.010 4.720 3.210 ;
        RECT 4.720 3.020 4.730 3.210 ;
        RECT 4.730 3.030 4.740 3.210 ;
        RECT 4.740 3.040 4.750 3.210 ;
        RECT 4.515 2.815 4.525 3.065 ;
        RECT 4.525 2.825 4.535 3.075 ;
        RECT 4.535 2.835 4.545 3.085 ;
        RECT 4.545 2.845 4.555 3.095 ;
        RECT 4.555 2.855 4.565 3.105 ;
        RECT 4.565 2.865 4.575 3.115 ;
        RECT 4.575 2.875 4.585 3.125 ;
        RECT 4.585 2.885 4.595 3.135 ;
        RECT 4.595 2.895 4.605 3.145 ;
        RECT 4.605 2.905 4.615 3.155 ;
        RECT 4.615 2.915 4.625 3.165 ;
        RECT 4.625 2.925 4.635 3.175 ;
        RECT 4.635 2.935 4.645 3.185 ;
        RECT 4.645 2.945 4.655 3.195 ;
        RECT 4.655 2.950 4.661 3.204 ;
        RECT 4.425 2.805 4.435 2.975 ;
        RECT 4.435 2.805 4.445 2.985 ;
        RECT 4.445 2.805 4.455 2.995 ;
        RECT 4.455 2.805 4.465 3.005 ;
        RECT 4.465 2.805 4.475 3.015 ;
        RECT 4.475 2.805 4.485 3.025 ;
        RECT 4.485 2.805 4.495 3.035 ;
        RECT 4.495 2.805 4.505 3.045 ;
        RECT 4.505 2.805 4.515 3.055 ;
        RECT 3.720 2.805 3.730 3.025 ;
        RECT 3.730 2.805 3.740 3.015 ;
        RECT 3.740 2.805 3.750 3.005 ;
        RECT 3.750 2.805 3.760 2.995 ;
        RECT 3.760 2.805 3.770 2.985 ;
        RECT 3.770 2.805 3.780 2.975 ;
        RECT 3.645 2.865 3.655 3.035 ;
        RECT 3.655 2.855 3.665 3.035 ;
        RECT 3.665 2.845 3.675 3.035 ;
        RECT 3.675 2.835 3.685 3.035 ;
        RECT 3.685 2.825 3.695 3.035 ;
        RECT 3.695 2.815 3.705 3.035 ;
        RECT 3.775 1.685 4.075 2.225 ;
        RECT 3.775 2.055 5.090 2.225 ;
        RECT 4.915 2.055 5.090 2.275 ;
        RECT 5.060 1.165 5.230 1.335 ;
        RECT 5.395 1.165 5.400 2.095 ;
        RECT 6.430 1.600 6.600 2.095 ;
        RECT 5.395 1.925 6.600 2.095 ;
        RECT 5.230 1.165 5.240 2.249 ;
        RECT 5.240 1.165 5.250 2.239 ;
        RECT 5.250 1.165 5.260 2.229 ;
        RECT 5.260 1.165 5.270 2.219 ;
        RECT 5.270 1.165 5.280 2.209 ;
        RECT 5.280 1.165 5.290 2.199 ;
        RECT 5.290 1.165 5.300 2.189 ;
        RECT 5.300 1.165 5.310 2.179 ;
        RECT 5.310 1.165 5.320 2.169 ;
        RECT 5.320 1.165 5.330 2.159 ;
        RECT 5.330 1.165 5.340 2.149 ;
        RECT 5.340 1.165 5.350 2.139 ;
        RECT 5.350 1.165 5.360 2.129 ;
        RECT 5.360 1.165 5.370 2.119 ;
        RECT 5.370 1.165 5.380 2.109 ;
        RECT 5.380 1.165 5.390 2.099 ;
        RECT 5.390 1.165 5.396 2.095 ;
        RECT 5.215 1.930 5.225 2.264 ;
        RECT 5.225 1.920 5.231 2.260 ;
        RECT 5.090 2.055 5.100 2.275 ;
        RECT 5.100 2.045 5.110 2.275 ;
        RECT 5.110 2.035 5.120 2.275 ;
        RECT 5.120 2.025 5.130 2.275 ;
        RECT 5.130 2.015 5.140 2.275 ;
        RECT 5.140 2.005 5.150 2.275 ;
        RECT 5.150 1.995 5.160 2.275 ;
        RECT 5.160 1.985 5.170 2.275 ;
        RECT 5.170 1.975 5.180 2.275 ;
        RECT 5.180 1.965 5.190 2.275 ;
        RECT 5.190 1.955 5.200 2.275 ;
        RECT 5.200 1.945 5.210 2.275 ;
        RECT 5.210 1.935 5.216 2.275 ;
        RECT 1.720 0.995 1.890 2.685 ;
        RECT 1.440 2.350 1.890 2.685 ;
        RECT 2.765 0.525 2.935 2.685 ;
        RECT 2.765 1.795 3.135 1.965 ;
        RECT 1.440 2.515 3.490 2.685 ;
        RECT 3.550 2.455 3.565 2.685 ;
        RECT 2.765 0.525 3.595 0.695 ;
        RECT 3.625 2.455 4.650 2.625 ;
        RECT 4.660 2.455 4.810 2.635 ;
        RECT 4.820 2.465 5.375 2.635 ;
        RECT 5.700 2.275 6.735 2.445 ;
        RECT 6.950 1.265 7.150 1.435 ;
        RECT 7.185 2.535 7.355 2.825 ;
        RECT 7.075 2.535 7.355 2.705 ;
        RECT 7.185 2.655 7.660 2.825 ;
        RECT 6.995 2.465 7.005 2.705 ;
        RECT 7.005 2.475 7.015 2.705 ;
        RECT 7.015 2.485 7.025 2.705 ;
        RECT 7.025 2.495 7.035 2.705 ;
        RECT 7.035 2.505 7.045 2.705 ;
        RECT 7.045 2.515 7.055 2.705 ;
        RECT 7.055 2.525 7.065 2.705 ;
        RECT 7.065 2.535 7.075 2.705 ;
        RECT 6.950 2.420 6.960 2.660 ;
        RECT 6.960 2.430 6.970 2.670 ;
        RECT 6.970 2.440 6.980 2.680 ;
        RECT 6.980 2.450 6.990 2.690 ;
        RECT 6.990 2.455 6.996 2.699 ;
        RECT 6.780 1.265 6.790 2.489 ;
        RECT 6.790 1.265 6.800 2.499 ;
        RECT 6.800 1.265 6.810 2.509 ;
        RECT 6.810 1.265 6.820 2.519 ;
        RECT 6.820 1.265 6.830 2.529 ;
        RECT 6.830 1.265 6.840 2.539 ;
        RECT 6.840 1.265 6.850 2.549 ;
        RECT 6.850 1.265 6.860 2.559 ;
        RECT 6.860 1.265 6.870 2.569 ;
        RECT 6.870 1.265 6.880 2.579 ;
        RECT 6.880 1.265 6.890 2.589 ;
        RECT 6.890 1.265 6.900 2.599 ;
        RECT 6.900 1.265 6.910 2.609 ;
        RECT 6.910 1.265 6.920 2.619 ;
        RECT 6.920 1.265 6.930 2.629 ;
        RECT 6.930 1.265 6.940 2.639 ;
        RECT 6.940 1.265 6.950 2.649 ;
        RECT 6.735 2.275 6.745 2.445 ;
        RECT 6.745 2.275 6.755 2.455 ;
        RECT 6.755 2.275 6.765 2.465 ;
        RECT 6.765 2.275 6.775 2.475 ;
        RECT 6.775 2.275 6.781 2.485 ;
        RECT 5.565 2.275 5.575 2.569 ;
        RECT 5.575 2.275 5.585 2.559 ;
        RECT 5.585 2.275 5.595 2.549 ;
        RECT 5.595 2.275 5.605 2.539 ;
        RECT 5.605 2.275 5.615 2.529 ;
        RECT 5.615 2.275 5.625 2.519 ;
        RECT 5.625 2.275 5.635 2.509 ;
        RECT 5.635 2.275 5.645 2.499 ;
        RECT 5.645 2.275 5.655 2.489 ;
        RECT 5.655 2.275 5.665 2.479 ;
        RECT 5.665 2.275 5.675 2.469 ;
        RECT 5.675 2.275 5.685 2.459 ;
        RECT 5.685 2.275 5.695 2.449 ;
        RECT 5.695 2.275 5.701 2.445 ;
        RECT 5.510 2.330 5.520 2.624 ;
        RECT 5.520 2.320 5.530 2.614 ;
        RECT 5.530 2.310 5.540 2.604 ;
        RECT 5.540 2.300 5.550 2.594 ;
        RECT 5.550 2.290 5.560 2.584 ;
        RECT 5.560 2.280 5.566 2.580 ;
        RECT 5.375 2.465 5.385 2.635 ;
        RECT 5.385 2.455 5.395 2.635 ;
        RECT 5.395 2.445 5.405 2.635 ;
        RECT 5.405 2.435 5.415 2.635 ;
        RECT 5.415 2.425 5.425 2.635 ;
        RECT 5.425 2.415 5.435 2.635 ;
        RECT 5.435 2.405 5.445 2.635 ;
        RECT 5.445 2.395 5.455 2.635 ;
        RECT 5.455 2.385 5.465 2.635 ;
        RECT 5.465 2.375 5.475 2.635 ;
        RECT 5.475 2.365 5.485 2.635 ;
        RECT 5.485 2.355 5.495 2.635 ;
        RECT 5.495 2.345 5.505 2.635 ;
        RECT 5.505 2.335 5.511 2.635 ;
        RECT 4.810 2.465 4.820 2.635 ;
        RECT 4.650 2.455 4.660 2.625 ;
        RECT 3.565 2.455 3.575 2.675 ;
        RECT 3.575 2.455 3.585 2.665 ;
        RECT 3.585 2.455 3.595 2.655 ;
        RECT 3.595 2.455 3.605 2.645 ;
        RECT 3.605 2.455 3.615 2.635 ;
        RECT 3.615 2.455 3.625 2.625 ;
        RECT 3.490 2.515 3.500 2.685 ;
        RECT 3.500 2.505 3.510 2.685 ;
        RECT 3.510 2.495 3.520 2.685 ;
        RECT 3.520 2.485 3.530 2.685 ;
        RECT 3.530 2.475 3.540 2.685 ;
        RECT 3.540 2.465 3.550 2.685 ;
        RECT 9.165 1.125 9.335 2.215 ;
        RECT 8.305 2.045 9.335 2.215 ;
        RECT 9.070 1.125 9.370 1.295 ;
        RECT 8.135 1.885 8.145 2.215 ;
        RECT 8.145 1.895 8.155 2.215 ;
        RECT 8.155 1.905 8.165 2.215 ;
        RECT 8.165 1.915 8.175 2.215 ;
        RECT 8.175 1.925 8.185 2.215 ;
        RECT 8.185 1.935 8.195 2.215 ;
        RECT 8.195 1.945 8.205 2.215 ;
        RECT 8.205 1.955 8.215 2.215 ;
        RECT 8.215 1.965 8.225 2.215 ;
        RECT 8.225 1.975 8.235 2.215 ;
        RECT 8.235 1.985 8.245 2.215 ;
        RECT 8.245 1.995 8.255 2.215 ;
        RECT 8.255 2.005 8.265 2.215 ;
        RECT 8.265 2.015 8.275 2.215 ;
        RECT 8.275 2.025 8.285 2.215 ;
        RECT 8.285 2.035 8.295 2.215 ;
        RECT 8.295 2.045 8.305 2.215 ;
        RECT 8.090 1.840 8.100 2.170 ;
        RECT 8.100 1.850 8.110 2.180 ;
        RECT 8.110 1.860 8.120 2.190 ;
        RECT 8.120 1.870 8.130 2.200 ;
        RECT 8.130 1.875 8.136 2.209 ;
        RECT 7.790 1.675 7.800 1.869 ;
        RECT 7.800 1.675 7.810 1.879 ;
        RECT 7.810 1.675 7.820 1.889 ;
        RECT 7.820 1.675 7.830 1.899 ;
        RECT 7.830 1.675 7.840 1.909 ;
        RECT 7.840 1.675 7.850 1.919 ;
        RECT 7.850 1.675 7.860 1.929 ;
        RECT 7.860 1.675 7.870 1.939 ;
        RECT 7.870 1.675 7.880 1.949 ;
        RECT 7.880 1.675 7.890 1.959 ;
        RECT 7.890 1.675 7.900 1.969 ;
        RECT 7.900 1.675 7.910 1.979 ;
        RECT 7.910 1.675 7.920 1.989 ;
        RECT 7.920 1.675 7.930 1.999 ;
        RECT 7.930 1.675 7.940 2.009 ;
        RECT 7.940 1.675 7.950 2.019 ;
        RECT 7.950 1.675 7.960 2.029 ;
        RECT 7.960 1.675 7.970 2.039 ;
        RECT 7.970 1.675 7.980 2.049 ;
        RECT 7.980 1.675 7.990 2.059 ;
        RECT 7.990 1.675 8.000 2.069 ;
        RECT 8.000 1.675 8.010 2.079 ;
        RECT 8.010 1.675 8.020 2.089 ;
        RECT 8.020 1.675 8.030 2.099 ;
        RECT 8.030 1.675 8.040 2.109 ;
        RECT 8.040 1.675 8.050 2.119 ;
        RECT 8.050 1.675 8.060 2.129 ;
        RECT 8.060 1.675 8.070 2.139 ;
        RECT 8.070 1.675 8.080 2.149 ;
        RECT 8.080 1.675 8.090 2.159 ;
        RECT 4.645 0.730 4.815 1.400 ;
        RECT 6.760 0.545 6.930 0.900 ;
        RECT 4.645 0.730 6.930 0.900 ;
        RECT 6.760 0.545 7.850 0.715 ;
        RECT 7.680 0.545 7.850 1.145 ;
        RECT 8.685 0.745 8.855 1.145 ;
        RECT 7.680 0.975 8.855 1.145 ;
        RECT 9.550 0.745 9.720 2.215 ;
        RECT 8.685 0.745 10.170 0.945 ;
        RECT 9.550 2.045 10.170 2.215 ;
        RECT 7.110 0.895 7.500 1.065 ;
        RECT 7.330 0.895 7.500 2.335 ;
        RECT 7.130 2.165 7.680 2.335 ;
        RECT 8.720 2.395 9.020 2.705 ;
        RECT 8.000 2.395 10.275 2.565 ;
        RECT 10.580 1.610 10.830 1.780 ;
        RECT 10.410 1.610 10.420 2.534 ;
        RECT 10.420 1.610 10.430 2.524 ;
        RECT 10.430 1.610 10.440 2.514 ;
        RECT 10.440 1.610 10.450 2.504 ;
        RECT 10.450 1.610 10.460 2.494 ;
        RECT 10.460 1.610 10.470 2.484 ;
        RECT 10.470 1.610 10.480 2.474 ;
        RECT 10.480 1.610 10.490 2.464 ;
        RECT 10.490 1.610 10.500 2.454 ;
        RECT 10.500 1.610 10.510 2.444 ;
        RECT 10.510 1.610 10.520 2.434 ;
        RECT 10.520 1.610 10.530 2.424 ;
        RECT 10.530 1.610 10.540 2.414 ;
        RECT 10.540 1.610 10.550 2.404 ;
        RECT 10.550 1.610 10.560 2.394 ;
        RECT 10.560 1.610 10.570 2.384 ;
        RECT 10.570 1.610 10.580 2.374 ;
        RECT 10.390 2.280 10.400 2.554 ;
        RECT 10.400 2.270 10.410 2.544 ;
        RECT 10.275 2.395 10.285 2.565 ;
        RECT 10.285 2.385 10.295 2.565 ;
        RECT 10.295 2.375 10.305 2.565 ;
        RECT 10.305 2.365 10.315 2.565 ;
        RECT 10.315 2.355 10.325 2.565 ;
        RECT 10.325 2.345 10.335 2.565 ;
        RECT 10.335 2.335 10.345 2.565 ;
        RECT 10.345 2.325 10.355 2.565 ;
        RECT 10.355 2.315 10.365 2.565 ;
        RECT 10.365 2.305 10.375 2.565 ;
        RECT 10.375 2.295 10.385 2.565 ;
        RECT 10.385 2.285 10.391 2.565 ;
        RECT 7.910 2.315 7.920 2.565 ;
        RECT 7.920 2.325 7.930 2.565 ;
        RECT 7.930 2.335 7.940 2.565 ;
        RECT 7.940 2.345 7.950 2.565 ;
        RECT 7.950 2.355 7.960 2.565 ;
        RECT 7.960 2.365 7.970 2.565 ;
        RECT 7.970 2.375 7.980 2.565 ;
        RECT 7.980 2.385 7.990 2.565 ;
        RECT 7.990 2.395 8.000 2.565 ;
        RECT 7.770 2.175 7.780 2.425 ;
        RECT 7.780 2.185 7.790 2.435 ;
        RECT 7.790 2.195 7.800 2.445 ;
        RECT 7.800 2.205 7.810 2.455 ;
        RECT 7.810 2.215 7.820 2.465 ;
        RECT 7.820 2.225 7.830 2.475 ;
        RECT 7.830 2.235 7.840 2.485 ;
        RECT 7.840 2.245 7.850 2.495 ;
        RECT 7.850 2.255 7.860 2.505 ;
        RECT 7.860 2.265 7.870 2.515 ;
        RECT 7.870 2.275 7.880 2.525 ;
        RECT 7.880 2.285 7.890 2.535 ;
        RECT 7.890 2.295 7.900 2.545 ;
        RECT 7.900 2.305 7.910 2.555 ;
        RECT 7.680 2.165 7.690 2.335 ;
        RECT 7.690 2.165 7.700 2.345 ;
        RECT 7.700 2.165 7.710 2.355 ;
        RECT 7.710 2.165 7.720 2.365 ;
        RECT 7.720 2.165 7.730 2.375 ;
        RECT 7.730 2.165 7.740 2.385 ;
        RECT 7.740 2.165 7.750 2.395 ;
        RECT 7.750 2.165 7.760 2.405 ;
        RECT 7.760 2.165 7.770 2.415 ;
  END 
END FFDSRHQHD1XHT

MACRO FFDSRHDMXHT
  CLASS  CORE ;
  FOREIGN FFDSRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.890 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.545 1.060 11.790 2.855 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.440 1.125 11.015 1.295 ;
        RECT 10.845 1.125 11.015 2.430 ;
        RECT 10.505 2.080 11.015 2.430 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.675 1.710 2.070 2.365 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.365 1.435 3.850 2.030 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.660 -0.300 0.830 0.670 ;
        RECT 1.730 -0.300 2.030 0.605 ;
        RECT 3.435 -0.300 3.735 1.160 ;
        RECT 6.215 -0.300 6.385 1.345 ;
        RECT 8.050 -0.300 8.350 0.740 ;
        RECT 9.930 -0.300 10.230 0.720 ;
        RECT 10.960 -0.300 11.260 0.595 ;
        RECT 0.000 -0.300 11.890 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.185 1.670 0.725 2.015 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 9.530 1.565 9.955 2.020 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.575 2.745 0.875 3.990 ;
        RECT 1.615 2.905 1.915 3.990 ;
        RECT 3.645 3.025 4.625 3.990 ;
        RECT 6.165 2.995 6.465 3.990 ;
        RECT 8.100 2.315 8.610 3.990 ;
        RECT 9.930 2.975 10.230 3.990 ;
        RECT 10.960 2.975 11.260 3.990 ;
        RECT 0.000 3.390 11.890 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 0.860 1.295 ;
        RECT 0.105 2.195 0.905 2.365 ;
        RECT 1.135 0.710 1.505 0.880 ;
        RECT 1.655 0.785 2.115 0.955 ;
        RECT 2.400 0.575 3.130 0.745 ;
        RECT 2.880 1.455 3.050 2.145 ;
        RECT 2.960 0.575 3.130 1.625 ;
        RECT 2.880 1.455 3.130 1.625 ;
        RECT 2.325 0.575 2.335 0.809 ;
        RECT 2.335 0.575 2.345 0.799 ;
        RECT 2.345 0.575 2.355 0.789 ;
        RECT 2.355 0.575 2.365 0.779 ;
        RECT 2.365 0.575 2.375 0.769 ;
        RECT 2.375 0.575 2.385 0.759 ;
        RECT 2.385 0.575 2.395 0.749 ;
        RECT 2.395 0.575 2.401 0.745 ;
        RECT 2.190 0.710 2.200 0.944 ;
        RECT 2.200 0.700 2.210 0.934 ;
        RECT 2.210 0.690 2.220 0.924 ;
        RECT 2.220 0.680 2.230 0.914 ;
        RECT 2.230 0.670 2.240 0.904 ;
        RECT 2.240 0.660 2.250 0.894 ;
        RECT 2.250 0.650 2.260 0.884 ;
        RECT 2.260 0.640 2.270 0.874 ;
        RECT 2.270 0.630 2.280 0.864 ;
        RECT 2.280 0.620 2.290 0.854 ;
        RECT 2.290 0.610 2.300 0.844 ;
        RECT 2.300 0.600 2.310 0.834 ;
        RECT 2.310 0.590 2.320 0.824 ;
        RECT 2.320 0.580 2.326 0.820 ;
        RECT 2.115 0.785 2.125 0.955 ;
        RECT 2.125 0.775 2.135 0.955 ;
        RECT 2.135 0.765 2.145 0.955 ;
        RECT 2.145 0.755 2.155 0.955 ;
        RECT 2.155 0.745 2.165 0.955 ;
        RECT 2.165 0.735 2.175 0.955 ;
        RECT 2.175 0.725 2.185 0.955 ;
        RECT 2.185 0.715 2.191 0.955 ;
        RECT 1.580 0.720 1.590 0.954 ;
        RECT 1.590 0.730 1.600 0.954 ;
        RECT 1.600 0.740 1.610 0.954 ;
        RECT 1.610 0.750 1.620 0.954 ;
        RECT 1.620 0.760 1.630 0.954 ;
        RECT 1.630 0.770 1.640 0.954 ;
        RECT 1.640 0.780 1.650 0.954 ;
        RECT 1.650 0.785 1.656 0.955 ;
        RECT 1.505 0.710 1.515 0.880 ;
        RECT 1.515 0.710 1.525 0.890 ;
        RECT 1.525 0.710 1.535 0.900 ;
        RECT 1.535 0.710 1.545 0.910 ;
        RECT 1.545 0.710 1.555 0.920 ;
        RECT 1.555 0.710 1.565 0.930 ;
        RECT 1.565 0.710 1.575 0.940 ;
        RECT 1.575 0.710 1.581 0.950 ;
        RECT 1.050 0.710 1.060 0.954 ;
        RECT 1.060 0.710 1.070 0.944 ;
        RECT 1.070 0.710 1.080 0.934 ;
        RECT 1.080 0.710 1.090 0.924 ;
        RECT 1.090 0.710 1.100 0.914 ;
        RECT 1.100 0.710 1.110 0.904 ;
        RECT 1.110 0.710 1.120 0.894 ;
        RECT 1.120 0.710 1.130 0.884 ;
        RECT 1.130 0.710 1.136 0.880 ;
        RECT 1.030 1.450 1.040 2.364 ;
        RECT 1.040 1.460 1.050 2.364 ;
        RECT 1.050 1.470 1.060 2.364 ;
        RECT 1.060 1.480 1.070 2.364 ;
        RECT 1.070 1.485 1.076 2.365 ;
        RECT 1.030 0.730 1.040 0.974 ;
        RECT 1.040 0.720 1.050 0.964 ;
        RECT 0.905 0.855 0.915 2.365 ;
        RECT 0.915 0.845 0.925 2.365 ;
        RECT 0.925 0.835 0.935 2.365 ;
        RECT 0.935 0.825 0.945 2.365 ;
        RECT 0.945 0.815 0.955 2.365 ;
        RECT 0.955 0.805 0.965 2.365 ;
        RECT 0.965 0.795 0.975 2.365 ;
        RECT 0.975 0.785 0.985 2.365 ;
        RECT 0.985 0.775 0.995 2.365 ;
        RECT 0.995 0.765 1.005 2.365 ;
        RECT 1.005 0.755 1.015 2.365 ;
        RECT 1.015 0.745 1.025 2.365 ;
        RECT 1.025 0.735 1.031 2.365 ;
        RECT 0.860 0.900 0.870 1.514 ;
        RECT 0.870 0.890 0.880 1.524 ;
        RECT 0.880 0.880 0.890 1.534 ;
        RECT 0.890 0.870 0.900 1.544 ;
        RECT 0.900 0.860 0.906 1.554 ;
        RECT 4.020 0.925 4.200 1.225 ;
        RECT 4.030 0.925 4.200 1.775 ;
        RECT 4.050 1.475 4.220 2.145 ;
        RECT 4.030 1.475 4.815 1.775 ;
        RECT 2.445 1.045 2.615 2.495 ;
        RECT 2.550 0.925 2.720 1.225 ;
        RECT 2.445 1.045 2.720 1.225 ;
        RECT 4.995 1.680 5.165 2.495 ;
        RECT 2.445 2.325 5.165 2.495 ;
        RECT 5.240 1.550 5.410 1.850 ;
        RECT 4.995 1.680 5.410 1.850 ;
        RECT 4.465 0.990 5.685 1.160 ;
        RECT 5.515 0.990 5.685 1.345 ;
        RECT 5.355 2.045 5.655 2.215 ;
        RECT 5.355 2.045 5.665 2.205 ;
        RECT 5.355 2.045 5.675 2.195 ;
        RECT 5.355 2.045 5.685 2.185 ;
        RECT 5.355 2.045 5.695 2.175 ;
        RECT 5.355 2.045 5.705 2.165 ;
        RECT 5.355 2.045 5.715 2.155 ;
        RECT 5.355 2.045 5.725 2.145 ;
        RECT 5.355 2.045 5.735 2.135 ;
        RECT 5.355 2.045 5.745 2.125 ;
        RECT 5.355 2.045 5.755 2.115 ;
        RECT 5.590 1.535 5.761 2.109 ;
        RECT 4.095 0.560 6.035 0.730 ;
        RECT 5.865 0.560 6.035 1.705 ;
        RECT 5.590 1.535 6.520 1.705 ;
        RECT 1.210 1.060 1.425 1.360 ;
        RECT 1.255 1.060 1.425 2.715 ;
        RECT 2.095 2.545 2.265 2.845 ;
        RECT 1.255 2.545 2.265 2.715 ;
        RECT 2.325 2.675 2.625 2.925 ;
        RECT 5.345 2.395 5.515 2.845 ;
        RECT 2.095 2.675 5.515 2.845 ;
        RECT 5.345 2.395 5.735 2.565 ;
        RECT 5.910 2.295 6.700 2.465 ;
        RECT 6.875 2.395 7.445 2.565 ;
        RECT 7.275 2.395 7.445 2.695 ;
        RECT 6.800 2.330 6.810 2.564 ;
        RECT 6.810 2.340 6.820 2.564 ;
        RECT 6.820 2.350 6.830 2.564 ;
        RECT 6.830 2.360 6.840 2.564 ;
        RECT 6.840 2.370 6.850 2.564 ;
        RECT 6.850 2.380 6.860 2.564 ;
        RECT 6.860 2.390 6.870 2.564 ;
        RECT 6.870 2.395 6.876 2.565 ;
        RECT 6.775 2.305 6.785 2.539 ;
        RECT 6.785 2.315 6.795 2.549 ;
        RECT 6.795 2.320 6.801 2.560 ;
        RECT 6.700 2.295 6.710 2.465 ;
        RECT 6.710 2.295 6.720 2.475 ;
        RECT 6.720 2.295 6.730 2.485 ;
        RECT 6.730 2.295 6.740 2.495 ;
        RECT 6.740 2.295 6.750 2.505 ;
        RECT 6.750 2.295 6.760 2.515 ;
        RECT 6.760 2.295 6.770 2.525 ;
        RECT 6.770 2.295 6.776 2.535 ;
        RECT 5.835 2.295 5.845 2.529 ;
        RECT 5.845 2.295 5.855 2.519 ;
        RECT 5.855 2.295 5.865 2.509 ;
        RECT 5.865 2.295 5.875 2.499 ;
        RECT 5.875 2.295 5.885 2.489 ;
        RECT 5.885 2.295 5.895 2.479 ;
        RECT 5.895 2.295 5.905 2.469 ;
        RECT 5.905 2.295 5.911 2.465 ;
        RECT 5.810 2.320 5.820 2.554 ;
        RECT 5.820 2.310 5.830 2.544 ;
        RECT 5.830 2.300 5.836 2.540 ;
        RECT 5.735 2.395 5.745 2.565 ;
        RECT 5.745 2.385 5.755 2.565 ;
        RECT 5.755 2.375 5.765 2.565 ;
        RECT 5.765 2.365 5.775 2.565 ;
        RECT 5.775 2.355 5.785 2.565 ;
        RECT 5.785 2.345 5.795 2.565 ;
        RECT 5.795 2.335 5.805 2.565 ;
        RECT 5.805 2.325 5.811 2.565 ;
        RECT 5.255 3.040 5.815 3.210 ;
        RECT 6.085 2.645 6.545 2.815 ;
        RECT 6.860 2.745 7.030 3.045 ;
        RECT 6.720 2.745 7.030 2.915 ;
        RECT 7.350 1.205 7.575 1.375 ;
        RECT 7.625 1.205 7.650 3.045 ;
        RECT 6.860 2.875 7.650 3.045 ;
        RECT 7.650 1.215 7.660 3.045 ;
        RECT 7.660 1.225 7.670 3.045 ;
        RECT 7.670 1.235 7.680 3.045 ;
        RECT 7.680 1.245 7.690 3.045 ;
        RECT 7.690 1.255 7.700 3.045 ;
        RECT 7.700 1.265 7.710 3.045 ;
        RECT 7.710 1.275 7.720 3.045 ;
        RECT 7.720 1.285 7.730 3.045 ;
        RECT 7.730 1.295 7.740 3.045 ;
        RECT 7.740 1.305 7.750 3.045 ;
        RECT 7.750 1.315 7.760 3.045 ;
        RECT 7.760 1.325 7.770 3.045 ;
        RECT 7.770 1.335 7.780 3.045 ;
        RECT 7.780 1.345 7.790 3.045 ;
        RECT 7.790 1.350 7.796 3.044 ;
        RECT 7.575 1.205 7.585 1.375 ;
        RECT 7.585 1.205 7.595 1.385 ;
        RECT 7.595 1.205 7.605 1.395 ;
        RECT 7.605 1.205 7.615 1.405 ;
        RECT 7.615 1.205 7.625 1.415 ;
        RECT 6.645 2.680 6.655 2.914 ;
        RECT 6.655 2.690 6.665 2.914 ;
        RECT 6.665 2.700 6.675 2.914 ;
        RECT 6.675 2.710 6.685 2.914 ;
        RECT 6.685 2.720 6.695 2.914 ;
        RECT 6.695 2.730 6.705 2.914 ;
        RECT 6.705 2.740 6.715 2.914 ;
        RECT 6.715 2.745 6.721 2.915 ;
        RECT 6.620 2.655 6.630 2.889 ;
        RECT 6.630 2.665 6.640 2.899 ;
        RECT 6.640 2.670 6.646 2.910 ;
        RECT 6.545 2.645 6.555 2.815 ;
        RECT 6.555 2.645 6.565 2.825 ;
        RECT 6.565 2.645 6.575 2.835 ;
        RECT 6.575 2.645 6.585 2.845 ;
        RECT 6.585 2.645 6.595 2.855 ;
        RECT 6.595 2.645 6.605 2.865 ;
        RECT 6.605 2.645 6.615 2.875 ;
        RECT 6.615 2.645 6.621 2.885 ;
        RECT 6.010 2.645 6.020 2.879 ;
        RECT 6.020 2.645 6.030 2.869 ;
        RECT 6.030 2.645 6.040 2.859 ;
        RECT 6.040 2.645 6.050 2.849 ;
        RECT 6.050 2.645 6.060 2.839 ;
        RECT 6.060 2.645 6.070 2.829 ;
        RECT 6.070 2.645 6.080 2.819 ;
        RECT 6.080 2.645 6.086 2.815 ;
        RECT 5.985 2.670 5.995 2.904 ;
        RECT 5.995 2.660 6.005 2.894 ;
        RECT 6.005 2.650 6.011 2.890 ;
        RECT 5.815 2.840 5.825 3.210 ;
        RECT 5.825 2.830 5.835 3.210 ;
        RECT 5.835 2.820 5.845 3.210 ;
        RECT 5.845 2.810 5.855 3.210 ;
        RECT 5.855 2.800 5.865 3.210 ;
        RECT 5.865 2.790 5.875 3.210 ;
        RECT 5.875 2.780 5.885 3.210 ;
        RECT 5.885 2.770 5.895 3.210 ;
        RECT 5.895 2.760 5.905 3.210 ;
        RECT 5.905 2.750 5.915 3.210 ;
        RECT 5.915 2.740 5.925 3.210 ;
        RECT 5.925 2.730 5.935 3.210 ;
        RECT 5.935 2.720 5.945 3.210 ;
        RECT 5.945 2.710 5.955 3.210 ;
        RECT 5.955 2.700 5.965 3.210 ;
        RECT 5.965 2.690 5.975 3.210 ;
        RECT 5.975 2.680 5.985 3.210 ;
        RECT 8.570 0.760 8.740 1.280 ;
        RECT 8.440 1.110 8.740 1.280 ;
        RECT 8.570 0.760 9.650 0.930 ;
        RECT 9.480 0.760 9.650 1.280 ;
        RECT 9.480 1.110 9.780 1.280 ;
        RECT 8.325 1.460 8.495 1.760 ;
        RECT 8.325 1.460 9.310 1.630 ;
        RECT 8.960 1.110 9.260 1.630 ;
        RECT 9.140 1.460 9.310 2.425 ;
        RECT 10.155 1.650 10.325 2.425 ;
        RECT 9.140 2.255 10.325 2.425 ;
        RECT 10.495 1.540 10.665 1.840 ;
        RECT 10.155 1.650 10.665 1.840 ;
        RECT 6.965 0.835 7.135 2.215 ;
        RECT 6.965 2.045 7.265 2.215 ;
        RECT 6.965 0.835 7.730 1.005 ;
        RECT 8.145 1.940 8.960 2.110 ;
        RECT 8.790 1.940 8.960 2.795 ;
        RECT 9.200 2.625 9.500 2.855 ;
        RECT 11.195 1.525 11.365 2.795 ;
        RECT 8.790 2.625 11.365 2.795 ;
        RECT 7.975 1.015 7.985 2.109 ;
        RECT 7.985 1.025 7.995 2.109 ;
        RECT 7.995 1.035 8.005 2.109 ;
        RECT 8.005 1.045 8.015 2.109 ;
        RECT 8.015 1.055 8.025 2.109 ;
        RECT 8.025 1.065 8.035 2.109 ;
        RECT 8.035 1.075 8.045 2.109 ;
        RECT 8.045 1.085 8.055 2.109 ;
        RECT 8.055 1.095 8.065 2.109 ;
        RECT 8.065 1.105 8.075 2.109 ;
        RECT 8.075 1.115 8.085 2.109 ;
        RECT 8.085 1.125 8.095 2.109 ;
        RECT 8.095 1.135 8.105 2.109 ;
        RECT 8.105 1.145 8.115 2.109 ;
        RECT 8.115 1.155 8.125 2.109 ;
        RECT 8.125 1.165 8.135 2.109 ;
        RECT 8.135 1.175 8.145 2.109 ;
        RECT 7.805 0.845 7.815 1.079 ;
        RECT 7.815 0.855 7.825 1.089 ;
        RECT 7.825 0.865 7.835 1.099 ;
        RECT 7.835 0.875 7.845 1.109 ;
        RECT 7.845 0.885 7.855 1.119 ;
        RECT 7.855 0.895 7.865 1.129 ;
        RECT 7.865 0.905 7.875 1.139 ;
        RECT 7.875 0.915 7.885 1.149 ;
        RECT 7.885 0.925 7.895 1.159 ;
        RECT 7.895 0.935 7.905 1.169 ;
        RECT 7.905 0.945 7.915 1.179 ;
        RECT 7.915 0.955 7.925 1.189 ;
        RECT 7.925 0.965 7.935 1.199 ;
        RECT 7.935 0.975 7.945 1.209 ;
        RECT 7.945 0.985 7.955 1.219 ;
        RECT 7.955 0.995 7.965 1.229 ;
        RECT 7.965 1.005 7.975 1.239 ;
        RECT 7.730 0.835 7.740 1.005 ;
        RECT 7.740 0.835 7.750 1.015 ;
        RECT 7.750 0.835 7.760 1.025 ;
        RECT 7.760 0.835 7.770 1.035 ;
        RECT 7.770 0.835 7.780 1.045 ;
        RECT 7.780 0.835 7.790 1.055 ;
        RECT 7.790 0.835 7.800 1.065 ;
        RECT 7.800 0.835 7.806 1.075 ;
  END 
END FFDSRHDMXHT

MACRO FFDSRHDLXHT
  CLASS  CORE ;
  FOREIGN FFDSRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.890 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.545 1.060 11.790 2.860 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.440 1.125 11.015 1.295 ;
        RECT 10.845 1.125 11.015 2.430 ;
        RECT 10.505 2.080 11.015 2.430 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.675 1.710 2.060 2.365 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.365 1.435 3.850 2.030 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.770 -0.300 1.750 0.530 ;
        RECT 3.435 -0.300 3.735 1.160 ;
        RECT 6.270 -0.300 6.440 0.875 ;
        RECT 8.025 -0.300 8.325 0.725 ;
        RECT 9.965 -0.300 10.265 0.810 ;
        RECT 10.960 -0.300 11.260 0.745 ;
        RECT 0.000 -0.300 11.890 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.195 1.670 0.725 2.015 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 9.530 1.565 9.955 2.020 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.575 2.625 0.875 3.990 ;
        RECT 1.585 2.905 1.885 3.990 ;
        RECT 3.645 3.025 4.625 3.990 ;
        RECT 6.165 2.995 6.465 3.990 ;
        RECT 8.100 2.290 8.610 3.990 ;
        RECT 9.990 2.975 10.290 3.990 ;
        RECT 10.960 2.975 11.260 3.990 ;
        RECT 0.000 3.390 11.890 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 1.030 1.295 ;
        RECT 0.860 0.710 1.030 1.514 ;
        RECT 0.870 1.485 1.076 1.524 ;
        RECT 0.880 1.485 1.076 1.534 ;
        RECT 0.890 1.485 1.076 1.544 ;
        RECT 0.900 1.485 1.076 1.554 ;
        RECT 0.105 2.195 1.030 2.365 ;
        RECT 0.860 1.450 1.040 1.514 ;
        RECT 0.860 1.460 1.050 1.514 ;
        RECT 0.860 1.470 1.060 1.514 ;
        RECT 0.905 1.480 1.070 2.364 ;
        RECT 1.070 1.485 1.076 2.365 ;
        RECT 1.930 0.620 2.100 0.880 ;
        RECT 0.860 0.710 2.100 0.880 ;
        RECT 1.930 0.620 3.170 0.790 ;
        RECT 2.880 1.340 3.050 2.145 ;
        RECT 3.000 0.620 3.170 1.510 ;
        RECT 2.880 1.340 3.170 1.510 ;
        RECT 4.020 0.925 4.200 1.225 ;
        RECT 4.030 0.925 4.200 1.775 ;
        RECT 4.050 1.475 4.220 2.145 ;
        RECT 4.030 1.475 4.815 1.775 ;
        RECT 2.445 0.990 2.615 2.495 ;
        RECT 2.445 0.990 2.785 1.160 ;
        RECT 4.995 1.680 5.165 2.495 ;
        RECT 2.445 2.325 5.165 2.495 ;
        RECT 5.240 1.550 5.410 1.850 ;
        RECT 4.995 1.680 5.410 1.850 ;
        RECT 4.465 0.990 5.740 1.160 ;
        RECT 5.570 0.990 5.740 1.345 ;
        RECT 5.355 2.045 5.655 2.215 ;
        RECT 5.355 2.045 5.665 2.205 ;
        RECT 5.355 2.045 5.675 2.195 ;
        RECT 5.355 2.045 5.685 2.185 ;
        RECT 5.355 2.045 5.695 2.175 ;
        RECT 5.355 2.045 5.705 2.165 ;
        RECT 5.355 2.045 5.715 2.155 ;
        RECT 5.355 2.045 5.725 2.145 ;
        RECT 5.355 2.045 5.735 2.135 ;
        RECT 5.355 2.045 5.745 2.125 ;
        RECT 5.355 2.045 5.755 2.115 ;
        RECT 5.590 1.535 5.761 2.109 ;
        RECT 4.095 0.560 6.090 0.730 ;
        RECT 5.920 0.560 6.090 1.705 ;
        RECT 5.590 1.535 6.530 1.705 ;
        RECT 1.210 1.060 1.425 1.360 ;
        RECT 1.255 1.060 1.425 2.715 ;
        RECT 2.095 2.545 2.265 2.845 ;
        RECT 1.255 2.545 2.265 2.715 ;
        RECT 2.295 2.675 2.595 2.925 ;
        RECT 5.345 2.395 5.515 2.845 ;
        RECT 2.095 2.675 5.515 2.845 ;
        RECT 5.345 2.395 5.735 2.565 ;
        RECT 5.910 2.295 6.700 2.465 ;
        RECT 6.875 2.395 7.445 2.565 ;
        RECT 7.275 2.395 7.445 2.695 ;
        RECT 6.800 2.330 6.810 2.564 ;
        RECT 6.810 2.340 6.820 2.564 ;
        RECT 6.820 2.350 6.830 2.564 ;
        RECT 6.830 2.360 6.840 2.564 ;
        RECT 6.840 2.370 6.850 2.564 ;
        RECT 6.850 2.380 6.860 2.564 ;
        RECT 6.860 2.390 6.870 2.564 ;
        RECT 6.870 2.395 6.876 2.565 ;
        RECT 6.775 2.305 6.785 2.539 ;
        RECT 6.785 2.315 6.795 2.549 ;
        RECT 6.795 2.320 6.801 2.560 ;
        RECT 6.700 2.295 6.710 2.465 ;
        RECT 6.710 2.295 6.720 2.475 ;
        RECT 6.720 2.295 6.730 2.485 ;
        RECT 6.730 2.295 6.740 2.495 ;
        RECT 6.740 2.295 6.750 2.505 ;
        RECT 6.750 2.295 6.760 2.515 ;
        RECT 6.760 2.295 6.770 2.525 ;
        RECT 6.770 2.295 6.776 2.535 ;
        RECT 5.835 2.295 5.845 2.529 ;
        RECT 5.845 2.295 5.855 2.519 ;
        RECT 5.855 2.295 5.865 2.509 ;
        RECT 5.865 2.295 5.875 2.499 ;
        RECT 5.875 2.295 5.885 2.489 ;
        RECT 5.885 2.295 5.895 2.479 ;
        RECT 5.895 2.295 5.905 2.469 ;
        RECT 5.905 2.295 5.911 2.465 ;
        RECT 5.810 2.320 5.820 2.554 ;
        RECT 5.820 2.310 5.830 2.544 ;
        RECT 5.830 2.300 5.836 2.540 ;
        RECT 5.735 2.395 5.745 2.565 ;
        RECT 5.745 2.385 5.755 2.565 ;
        RECT 5.755 2.375 5.765 2.565 ;
        RECT 5.765 2.365 5.775 2.565 ;
        RECT 5.775 2.355 5.785 2.565 ;
        RECT 5.785 2.345 5.795 2.565 ;
        RECT 5.795 2.335 5.805 2.565 ;
        RECT 5.805 2.325 5.811 2.565 ;
        RECT 5.255 3.040 5.815 3.210 ;
        RECT 6.085 2.645 6.545 2.815 ;
        RECT 6.860 2.745 7.030 3.045 ;
        RECT 6.720 2.745 7.030 2.915 ;
        RECT 7.335 1.205 7.575 1.375 ;
        RECT 7.625 1.205 7.650 3.045 ;
        RECT 6.860 2.875 7.650 3.045 ;
        RECT 7.650 1.215 7.660 3.045 ;
        RECT 7.660 1.225 7.670 3.045 ;
        RECT 7.670 1.235 7.680 3.045 ;
        RECT 7.680 1.245 7.690 3.045 ;
        RECT 7.690 1.255 7.700 3.045 ;
        RECT 7.700 1.265 7.710 3.045 ;
        RECT 7.710 1.275 7.720 3.045 ;
        RECT 7.720 1.285 7.730 3.045 ;
        RECT 7.730 1.295 7.740 3.045 ;
        RECT 7.740 1.305 7.750 3.045 ;
        RECT 7.750 1.315 7.760 3.045 ;
        RECT 7.760 1.325 7.770 3.045 ;
        RECT 7.770 1.335 7.780 3.045 ;
        RECT 7.780 1.345 7.790 3.045 ;
        RECT 7.790 1.350 7.796 3.044 ;
        RECT 7.575 1.205 7.585 1.375 ;
        RECT 7.585 1.205 7.595 1.385 ;
        RECT 7.595 1.205 7.605 1.395 ;
        RECT 7.605 1.205 7.615 1.405 ;
        RECT 7.615 1.205 7.625 1.415 ;
        RECT 6.645 2.680 6.655 2.914 ;
        RECT 6.655 2.690 6.665 2.914 ;
        RECT 6.665 2.700 6.675 2.914 ;
        RECT 6.675 2.710 6.685 2.914 ;
        RECT 6.685 2.720 6.695 2.914 ;
        RECT 6.695 2.730 6.705 2.914 ;
        RECT 6.705 2.740 6.715 2.914 ;
        RECT 6.715 2.745 6.721 2.915 ;
        RECT 6.620 2.655 6.630 2.889 ;
        RECT 6.630 2.665 6.640 2.899 ;
        RECT 6.640 2.670 6.646 2.910 ;
        RECT 6.545 2.645 6.555 2.815 ;
        RECT 6.555 2.645 6.565 2.825 ;
        RECT 6.565 2.645 6.575 2.835 ;
        RECT 6.575 2.645 6.585 2.845 ;
        RECT 6.585 2.645 6.595 2.855 ;
        RECT 6.595 2.645 6.605 2.865 ;
        RECT 6.605 2.645 6.615 2.875 ;
        RECT 6.615 2.645 6.621 2.885 ;
        RECT 6.010 2.645 6.020 2.879 ;
        RECT 6.020 2.645 6.030 2.869 ;
        RECT 6.030 2.645 6.040 2.859 ;
        RECT 6.040 2.645 6.050 2.849 ;
        RECT 6.050 2.645 6.060 2.839 ;
        RECT 6.060 2.645 6.070 2.829 ;
        RECT 6.070 2.645 6.080 2.819 ;
        RECT 6.080 2.645 6.086 2.815 ;
        RECT 5.985 2.670 5.995 2.904 ;
        RECT 5.995 2.660 6.005 2.894 ;
        RECT 6.005 2.650 6.011 2.890 ;
        RECT 5.815 2.840 5.825 3.210 ;
        RECT 5.825 2.830 5.835 3.210 ;
        RECT 5.835 2.820 5.845 3.210 ;
        RECT 5.845 2.810 5.855 3.210 ;
        RECT 5.855 2.800 5.865 3.210 ;
        RECT 5.865 2.790 5.875 3.210 ;
        RECT 5.875 2.780 5.885 3.210 ;
        RECT 5.885 2.770 5.895 3.210 ;
        RECT 5.895 2.760 5.905 3.210 ;
        RECT 5.905 2.750 5.915 3.210 ;
        RECT 5.915 2.740 5.925 3.210 ;
        RECT 5.925 2.730 5.935 3.210 ;
        RECT 5.935 2.720 5.945 3.210 ;
        RECT 5.945 2.710 5.955 3.210 ;
        RECT 5.955 2.700 5.965 3.210 ;
        RECT 5.965 2.690 5.975 3.210 ;
        RECT 5.975 2.680 5.985 3.210 ;
        RECT 8.570 0.760 8.740 1.280 ;
        RECT 8.415 1.110 8.740 1.280 ;
        RECT 9.450 0.640 9.750 0.930 ;
        RECT 8.570 0.760 9.750 0.930 ;
        RECT 8.325 1.460 8.495 1.760 ;
        RECT 8.325 1.460 9.310 1.630 ;
        RECT 8.995 1.110 9.295 1.630 ;
        RECT 9.140 1.460 9.310 2.425 ;
        RECT 10.155 1.650 10.325 2.425 ;
        RECT 9.140 2.255 10.325 2.425 ;
        RECT 10.495 1.540 10.665 1.840 ;
        RECT 10.155 1.650 10.665 1.840 ;
        RECT 6.965 0.835 7.135 2.215 ;
        RECT 6.965 2.045 7.265 2.215 ;
        RECT 6.965 0.835 7.730 1.005 ;
        RECT 8.145 1.940 8.960 2.110 ;
        RECT 8.790 1.940 8.960 2.795 ;
        RECT 11.195 1.525 11.365 2.795 ;
        RECT 8.790 2.625 11.365 2.795 ;
        RECT 7.975 1.015 7.985 2.109 ;
        RECT 7.985 1.025 7.995 2.109 ;
        RECT 7.995 1.035 8.005 2.109 ;
        RECT 8.005 1.045 8.015 2.109 ;
        RECT 8.015 1.055 8.025 2.109 ;
        RECT 8.025 1.065 8.035 2.109 ;
        RECT 8.035 1.075 8.045 2.109 ;
        RECT 8.045 1.085 8.055 2.109 ;
        RECT 8.055 1.095 8.065 2.109 ;
        RECT 8.065 1.105 8.075 2.109 ;
        RECT 8.075 1.115 8.085 2.109 ;
        RECT 8.085 1.125 8.095 2.109 ;
        RECT 8.095 1.135 8.105 2.109 ;
        RECT 8.105 1.145 8.115 2.109 ;
        RECT 8.115 1.155 8.125 2.109 ;
        RECT 8.125 1.165 8.135 2.109 ;
        RECT 8.135 1.175 8.145 2.109 ;
        RECT 7.805 0.845 7.815 1.079 ;
        RECT 7.815 0.855 7.825 1.089 ;
        RECT 7.825 0.865 7.835 1.099 ;
        RECT 7.835 0.875 7.845 1.109 ;
        RECT 7.845 0.885 7.855 1.119 ;
        RECT 7.855 0.895 7.865 1.129 ;
        RECT 7.865 0.905 7.875 1.139 ;
        RECT 7.875 0.915 7.885 1.149 ;
        RECT 7.885 0.925 7.895 1.159 ;
        RECT 7.895 0.935 7.905 1.169 ;
        RECT 7.905 0.945 7.915 1.179 ;
        RECT 7.915 0.955 7.925 1.189 ;
        RECT 7.925 0.965 7.935 1.199 ;
        RECT 7.935 0.975 7.945 1.209 ;
        RECT 7.945 0.985 7.955 1.219 ;
        RECT 7.955 0.995 7.965 1.229 ;
        RECT 7.965 1.005 7.975 1.239 ;
        RECT 7.730 0.835 7.740 1.005 ;
        RECT 7.740 0.835 7.750 1.015 ;
        RECT 7.750 0.835 7.760 1.025 ;
        RECT 7.760 0.835 7.770 1.035 ;
        RECT 7.770 0.835 7.780 1.045 ;
        RECT 7.780 0.835 7.790 1.055 ;
        RECT 7.790 0.835 7.800 1.065 ;
        RECT 7.800 0.835 7.806 1.075 ;
  END 
END FFDSRHDLXHT

MACRO FFDSRHD2XHT
  CLASS  CORE ;
  FOREIGN FFDSRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.530 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 12.670 0.720 12.840 1.470 ;
        RECT 12.670 1.300 13.075 1.470 ;
        RECT 12.605 2.045 12.905 2.895 ;
        RECT 12.905 1.300 13.075 2.430 ;
        RECT 12.605 2.045 13.075 2.430 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.565 1.190 11.975 1.360 ;
        RECT 11.805 0.785 11.865 2.320 ;
        RECT 11.565 0.785 11.865 1.360 ;
        RECT 11.805 1.190 11.975 2.320 ;
        RECT 11.565 2.150 11.975 2.320 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.640 1.540 1.970 2.455 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.380 1.465 3.590 2.060 ;
        RECT 3.380 1.465 3.810 1.765 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.715 ;
        RECT 1.525 -0.300 1.825 0.805 ;
        RECT 3.335 -0.300 3.635 1.185 ;
        RECT 6.195 -0.300 6.495 0.955 ;
        RECT 8.375 -0.300 8.675 0.665 ;
        RECT 10.670 -0.300 11.310 1.055 ;
        RECT 12.150 -0.300 12.320 1.120 ;
        RECT 13.125 -0.300 13.425 1.055 ;
        RECT 0.000 -0.300 13.530 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.475 0.320 2.015 ;
        RECT 0.100 1.475 0.495 1.775 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 10.630 1.235 10.800 1.840 ;
        RECT 10.630 1.235 11.085 1.540 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 2.795 0.865 3.990 ;
        RECT 1.525 3.030 1.825 3.990 ;
        RECT 3.540 3.025 4.520 3.990 ;
        RECT 6.225 3.025 6.525 3.990 ;
        RECT 8.300 2.530 8.470 3.990 ;
        RECT 10.075 3.025 10.375 3.990 ;
        RECT 11.045 2.975 11.345 3.990 ;
        RECT 12.085 2.975 12.385 3.990 ;
        RECT 13.125 2.635 13.425 3.990 ;
        RECT 0.000 3.390 13.530 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.195 0.570 2.365 ;
        RECT 0.105 1.125 0.830 1.295 ;
        RECT 0.830 1.125 0.840 2.179 ;
        RECT 0.840 1.125 0.850 2.169 ;
        RECT 0.850 1.125 0.860 2.159 ;
        RECT 0.860 1.125 0.870 2.149 ;
        RECT 0.870 1.125 0.880 2.139 ;
        RECT 0.880 1.125 0.890 2.129 ;
        RECT 0.890 1.125 0.900 2.119 ;
        RECT 0.900 1.125 0.910 2.109 ;
        RECT 0.910 1.125 0.920 2.099 ;
        RECT 0.920 1.125 0.930 2.089 ;
        RECT 0.930 1.125 0.940 2.079 ;
        RECT 0.940 1.125 0.950 2.069 ;
        RECT 0.950 1.125 0.960 2.059 ;
        RECT 0.960 1.125 0.970 2.049 ;
        RECT 0.970 1.125 0.980 2.039 ;
        RECT 0.980 1.125 0.990 2.029 ;
        RECT 0.990 1.125 1.000 2.019 ;
        RECT 0.655 2.110 0.665 2.354 ;
        RECT 0.665 2.100 0.675 2.344 ;
        RECT 0.675 2.090 0.685 2.334 ;
        RECT 0.685 2.080 0.695 2.324 ;
        RECT 0.695 2.070 0.705 2.314 ;
        RECT 0.705 2.060 0.715 2.304 ;
        RECT 0.715 2.050 0.725 2.294 ;
        RECT 0.725 2.040 0.735 2.284 ;
        RECT 0.735 2.030 0.745 2.274 ;
        RECT 0.745 2.020 0.755 2.264 ;
        RECT 0.755 2.010 0.765 2.254 ;
        RECT 0.765 2.000 0.775 2.244 ;
        RECT 0.775 1.990 0.785 2.234 ;
        RECT 0.785 1.980 0.795 2.224 ;
        RECT 0.795 1.970 0.805 2.214 ;
        RECT 0.805 1.960 0.815 2.204 ;
        RECT 0.815 1.950 0.825 2.194 ;
        RECT 0.825 1.940 0.831 2.190 ;
        RECT 0.570 2.195 0.580 2.365 ;
        RECT 0.580 2.185 0.590 2.365 ;
        RECT 0.590 2.175 0.600 2.365 ;
        RECT 0.600 2.165 0.610 2.365 ;
        RECT 0.610 2.155 0.620 2.365 ;
        RECT 0.620 2.145 0.630 2.365 ;
        RECT 0.630 2.135 0.640 2.365 ;
        RECT 0.640 2.125 0.650 2.365 ;
        RECT 0.650 2.115 0.656 2.365 ;
        RECT 2.265 0.545 3.030 0.715 ;
        RECT 2.860 0.545 3.030 2.125 ;
        RECT 2.775 1.955 3.075 2.125 ;
        RECT 3.865 1.015 4.165 1.185 ;
        RECT 3.995 1.015 4.165 2.145 ;
        RECT 3.915 1.975 4.215 2.145 ;
        RECT 3.995 1.485 4.815 1.655 ;
        RECT 2.425 0.950 2.595 2.495 ;
        RECT 2.425 0.950 2.680 1.250 ;
        RECT 4.580 1.835 4.750 2.495 ;
        RECT 2.425 2.325 4.750 2.495 ;
        RECT 4.580 1.835 4.955 2.005 ;
        RECT 5.025 1.675 5.040 2.005 ;
        RECT 5.200 1.675 5.325 1.845 ;
        RECT 5.040 1.675 5.050 1.995 ;
        RECT 5.050 1.675 5.060 1.985 ;
        RECT 5.060 1.675 5.070 1.975 ;
        RECT 5.070 1.675 5.080 1.965 ;
        RECT 5.080 1.675 5.090 1.955 ;
        RECT 5.090 1.675 5.100 1.945 ;
        RECT 5.100 1.675 5.110 1.935 ;
        RECT 5.110 1.675 5.120 1.925 ;
        RECT 5.120 1.675 5.130 1.915 ;
        RECT 5.130 1.675 5.140 1.905 ;
        RECT 5.140 1.675 5.150 1.895 ;
        RECT 5.150 1.675 5.160 1.885 ;
        RECT 5.160 1.675 5.170 1.875 ;
        RECT 5.170 1.675 5.180 1.865 ;
        RECT 5.180 1.675 5.190 1.855 ;
        RECT 5.190 1.675 5.200 1.845 ;
        RECT 4.955 1.835 4.965 2.005 ;
        RECT 4.965 1.825 4.975 2.005 ;
        RECT 4.975 1.815 4.985 2.005 ;
        RECT 4.985 1.805 4.995 2.005 ;
        RECT 4.995 1.795 5.005 2.005 ;
        RECT 5.005 1.785 5.015 2.005 ;
        RECT 5.015 1.775 5.025 2.005 ;
        RECT 4.375 0.985 4.675 1.305 ;
        RECT 5.480 0.920 5.650 1.305 ;
        RECT 4.375 1.135 5.650 1.305 ;
        RECT 4.005 0.480 4.305 0.740 ;
        RECT 4.895 0.570 5.195 0.955 ;
        RECT 5.530 1.590 5.700 2.215 ;
        RECT 5.400 2.045 5.700 2.215 ;
        RECT 4.005 0.570 6.000 0.740 ;
        RECT 5.830 0.570 6.000 1.760 ;
        RECT 5.530 1.590 6.735 1.760 ;
        RECT 1.150 2.130 1.350 2.430 ;
        RECT 1.180 1.060 1.350 2.845 ;
        RECT 2.225 2.675 2.525 3.085 ;
        RECT 4.990 2.470 5.160 2.845 ;
        RECT 1.180 2.675 5.160 2.845 ;
        RECT 4.990 2.470 5.720 2.640 ;
        RECT 5.940 2.325 6.795 2.495 ;
        RECT 7.560 1.585 7.730 2.630 ;
        RECT 7.005 2.460 7.730 2.630 ;
        RECT 6.930 2.395 6.940 2.629 ;
        RECT 6.940 2.405 6.950 2.629 ;
        RECT 6.950 2.415 6.960 2.629 ;
        RECT 6.960 2.425 6.970 2.629 ;
        RECT 6.970 2.435 6.980 2.629 ;
        RECT 6.980 2.445 6.990 2.629 ;
        RECT 6.990 2.455 7.000 2.629 ;
        RECT 7.000 2.460 7.006 2.630 ;
        RECT 6.870 2.335 6.880 2.569 ;
        RECT 6.880 2.345 6.890 2.579 ;
        RECT 6.890 2.355 6.900 2.589 ;
        RECT 6.900 2.365 6.910 2.599 ;
        RECT 6.910 2.375 6.920 2.609 ;
        RECT 6.920 2.385 6.930 2.619 ;
        RECT 6.795 2.325 6.805 2.495 ;
        RECT 6.805 2.325 6.815 2.505 ;
        RECT 6.815 2.325 6.825 2.515 ;
        RECT 6.825 2.325 6.835 2.525 ;
        RECT 6.835 2.325 6.845 2.535 ;
        RECT 6.845 2.325 6.855 2.545 ;
        RECT 6.855 2.325 6.865 2.555 ;
        RECT 6.865 2.325 6.871 2.565 ;
        RECT 5.865 2.325 5.875 2.559 ;
        RECT 5.875 2.325 5.885 2.549 ;
        RECT 5.885 2.325 5.895 2.539 ;
        RECT 5.895 2.325 5.905 2.529 ;
        RECT 5.905 2.325 5.915 2.519 ;
        RECT 5.915 2.325 5.925 2.509 ;
        RECT 5.925 2.325 5.935 2.499 ;
        RECT 5.935 2.325 5.941 2.495 ;
        RECT 5.795 2.395 5.805 2.629 ;
        RECT 5.805 2.385 5.815 2.619 ;
        RECT 5.815 2.375 5.825 2.609 ;
        RECT 5.825 2.365 5.835 2.599 ;
        RECT 5.835 2.355 5.845 2.589 ;
        RECT 5.845 2.345 5.855 2.579 ;
        RECT 5.855 2.335 5.865 2.569 ;
        RECT 5.720 2.470 5.730 2.640 ;
        RECT 5.730 2.460 5.740 2.640 ;
        RECT 5.740 2.450 5.750 2.640 ;
        RECT 5.750 2.440 5.760 2.640 ;
        RECT 5.760 2.430 5.770 2.640 ;
        RECT 5.770 2.420 5.780 2.640 ;
        RECT 5.780 2.410 5.790 2.640 ;
        RECT 5.790 2.400 5.796 2.640 ;
        RECT 5.535 2.825 5.835 3.210 ;
        RECT 5.535 2.825 5.870 3.005 ;
        RECT 6.095 2.675 6.640 2.845 ;
        RECT 7.425 2.810 7.725 2.995 ;
        RECT 7.560 1.155 8.080 1.325 ;
        RECT 7.910 1.155 8.080 2.980 ;
        RECT 6.850 2.810 8.080 2.980 ;
        RECT 6.775 2.745 6.785 2.979 ;
        RECT 6.785 2.755 6.795 2.979 ;
        RECT 6.795 2.765 6.805 2.979 ;
        RECT 6.805 2.775 6.815 2.979 ;
        RECT 6.815 2.785 6.825 2.979 ;
        RECT 6.825 2.795 6.835 2.979 ;
        RECT 6.835 2.805 6.845 2.979 ;
        RECT 6.845 2.810 6.851 2.980 ;
        RECT 6.715 2.685 6.725 2.919 ;
        RECT 6.725 2.695 6.735 2.929 ;
        RECT 6.735 2.705 6.745 2.939 ;
        RECT 6.745 2.715 6.755 2.949 ;
        RECT 6.755 2.725 6.765 2.959 ;
        RECT 6.765 2.735 6.775 2.969 ;
        RECT 6.640 2.675 6.650 2.845 ;
        RECT 6.650 2.675 6.660 2.855 ;
        RECT 6.660 2.675 6.670 2.865 ;
        RECT 6.670 2.675 6.680 2.875 ;
        RECT 6.680 2.675 6.690 2.885 ;
        RECT 6.690 2.675 6.700 2.895 ;
        RECT 6.700 2.675 6.710 2.905 ;
        RECT 6.710 2.675 6.716 2.915 ;
        RECT 6.020 2.675 6.030 2.909 ;
        RECT 6.030 2.675 6.040 2.899 ;
        RECT 6.040 2.675 6.050 2.889 ;
        RECT 6.050 2.675 6.060 2.879 ;
        RECT 6.060 2.675 6.070 2.869 ;
        RECT 6.070 2.675 6.080 2.859 ;
        RECT 6.080 2.675 6.090 2.849 ;
        RECT 6.090 2.675 6.096 2.845 ;
        RECT 5.935 2.760 5.945 2.994 ;
        RECT 5.945 2.750 5.955 2.984 ;
        RECT 5.955 2.740 5.965 2.974 ;
        RECT 5.965 2.730 5.975 2.964 ;
        RECT 5.975 2.720 5.985 2.954 ;
        RECT 5.985 2.710 5.995 2.944 ;
        RECT 5.995 2.700 6.005 2.934 ;
        RECT 6.005 2.690 6.015 2.924 ;
        RECT 6.015 2.680 6.021 2.920 ;
        RECT 5.870 2.825 5.880 3.005 ;
        RECT 5.880 2.815 5.890 3.005 ;
        RECT 5.890 2.805 5.900 3.005 ;
        RECT 5.900 2.795 5.910 3.005 ;
        RECT 5.910 2.785 5.920 3.005 ;
        RECT 5.920 2.775 5.930 3.005 ;
        RECT 5.930 2.765 5.936 3.005 ;
        RECT 8.610 1.570 8.910 1.805 ;
        RECT 8.610 1.570 10.050 1.740 ;
        RECT 9.880 1.570 10.050 2.125 ;
        RECT 8.885 0.700 9.185 0.920 ;
        RECT 8.885 0.700 10.320 0.870 ;
        RECT 10.020 0.700 10.320 0.920 ;
        RECT 8.610 1.090 8.780 1.390 ;
        RECT 9.405 1.050 9.705 1.390 ;
        RECT 8.610 1.220 10.450 1.390 ;
        RECT 10.280 1.220 10.450 2.495 ;
        RECT 9.155 2.325 10.450 2.495 ;
        RECT 11.020 1.780 11.190 2.215 ;
        RECT 10.280 2.045 11.190 2.215 ;
        RECT 11.450 1.540 11.620 1.950 ;
        RECT 11.020 1.780 11.620 1.950 ;
        RECT 7.210 0.785 7.380 2.280 ;
        RECT 7.210 0.785 8.160 0.955 ;
        RECT 8.430 2.075 8.905 2.245 ;
        RECT 8.805 2.075 8.905 2.845 ;
        RECT 9.100 1.955 9.490 2.125 ;
        RECT 10.705 2.515 10.875 2.845 ;
        RECT 8.975 2.675 10.875 2.845 ;
        RECT 10.705 2.515 12.380 2.710 ;
        RECT 12.210 1.650 12.380 2.710 ;
        RECT 12.210 1.650 12.725 1.820 ;
        RECT 9.025 1.955 9.035 2.189 ;
        RECT 9.035 1.955 9.045 2.179 ;
        RECT 9.045 1.955 9.055 2.169 ;
        RECT 9.055 1.955 9.065 2.159 ;
        RECT 9.065 1.955 9.075 2.149 ;
        RECT 9.075 1.955 9.085 2.139 ;
        RECT 9.085 1.955 9.095 2.129 ;
        RECT 9.095 1.955 9.101 2.125 ;
        RECT 8.975 2.005 8.985 2.239 ;
        RECT 8.985 1.995 8.995 2.229 ;
        RECT 8.995 1.985 9.005 2.219 ;
        RECT 9.005 1.975 9.015 2.209 ;
        RECT 9.015 1.965 9.025 2.199 ;
        RECT 8.905 2.075 8.915 2.845 ;
        RECT 8.915 2.065 8.925 2.845 ;
        RECT 8.925 2.055 8.935 2.845 ;
        RECT 8.935 2.045 8.945 2.845 ;
        RECT 8.945 2.035 8.955 2.845 ;
        RECT 8.955 2.025 8.965 2.845 ;
        RECT 8.965 2.015 8.975 2.845 ;
        RECT 8.260 0.820 8.270 2.244 ;
        RECT 8.270 0.830 8.280 2.244 ;
        RECT 8.280 0.840 8.290 2.244 ;
        RECT 8.290 0.850 8.300 2.244 ;
        RECT 8.300 0.860 8.310 2.244 ;
        RECT 8.310 0.870 8.320 2.244 ;
        RECT 8.320 0.880 8.330 2.244 ;
        RECT 8.330 0.890 8.340 2.244 ;
        RECT 8.340 0.900 8.350 2.244 ;
        RECT 8.350 0.910 8.360 2.244 ;
        RECT 8.360 0.920 8.370 2.244 ;
        RECT 8.370 0.930 8.380 2.244 ;
        RECT 8.380 0.940 8.390 2.244 ;
        RECT 8.390 0.950 8.400 2.244 ;
        RECT 8.400 0.960 8.410 2.244 ;
        RECT 8.410 0.970 8.420 2.244 ;
        RECT 8.420 0.980 8.430 2.244 ;
        RECT 8.235 0.795 8.245 1.029 ;
        RECT 8.245 0.805 8.255 1.039 ;
        RECT 8.255 0.810 8.261 1.050 ;
        RECT 8.160 0.785 8.170 0.955 ;
        RECT 8.170 0.785 8.180 0.965 ;
        RECT 8.180 0.785 8.190 0.975 ;
        RECT 8.190 0.785 8.200 0.985 ;
        RECT 8.200 0.785 8.210 0.995 ;
        RECT 8.210 0.785 8.220 1.005 ;
        RECT 8.220 0.785 8.230 1.015 ;
        RECT 8.230 0.785 8.236 1.025 ;
  END 
END FFDSRHD2XHT

MACRO FFDSRHD1XHT
  CLASS  CORE ;
  FOREIGN FFDSRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.890 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.545 0.720 11.790 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.505 0.720 10.675 1.360 ;
        RECT 10.505 1.155 11.015 1.360 ;
        RECT 10.845 1.155 11.015 2.430 ;
        RECT 10.505 2.080 11.015 2.430 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.675 1.710 2.070 2.365 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.365 1.435 3.850 2.030 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.660 -0.300 0.830 0.670 ;
        RECT 1.730 -0.300 2.030 0.605 ;
        RECT 3.435 -0.300 3.735 1.160 ;
        RECT 6.230 -0.300 6.400 1.310 ;
        RECT 8.025 -0.300 8.325 0.770 ;
        RECT 9.930 -0.300 10.230 0.680 ;
        RECT 10.960 -0.300 11.260 0.715 ;
        RECT 0.000 -0.300 11.890 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.190 1.670 0.725 2.015 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 9.530 1.515 9.955 2.020 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.575 2.745 0.875 3.990 ;
        RECT 1.615 2.905 1.915 3.990 ;
        RECT 3.575 3.025 4.215 3.990 ;
        RECT 6.165 2.995 6.465 3.990 ;
        RECT 8.100 2.350 8.610 3.990 ;
        RECT 9.930 2.975 10.230 3.990 ;
        RECT 10.960 2.975 11.260 3.990 ;
        RECT 0.000 3.390 11.890 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 0.860 1.295 ;
        RECT 0.105 2.195 0.905 2.365 ;
        RECT 1.135 0.710 1.505 0.880 ;
        RECT 1.655 0.785 2.115 0.955 ;
        RECT 2.400 0.575 3.130 0.745 ;
        RECT 2.880 1.455 3.050 2.145 ;
        RECT 2.960 0.575 3.130 1.625 ;
        RECT 2.880 1.455 3.130 1.625 ;
        RECT 2.325 0.575 2.335 0.809 ;
        RECT 2.335 0.575 2.345 0.799 ;
        RECT 2.345 0.575 2.355 0.789 ;
        RECT 2.355 0.575 2.365 0.779 ;
        RECT 2.365 0.575 2.375 0.769 ;
        RECT 2.375 0.575 2.385 0.759 ;
        RECT 2.385 0.575 2.395 0.749 ;
        RECT 2.395 0.575 2.401 0.745 ;
        RECT 2.190 0.710 2.200 0.944 ;
        RECT 2.200 0.700 2.210 0.934 ;
        RECT 2.210 0.690 2.220 0.924 ;
        RECT 2.220 0.680 2.230 0.914 ;
        RECT 2.230 0.670 2.240 0.904 ;
        RECT 2.240 0.660 2.250 0.894 ;
        RECT 2.250 0.650 2.260 0.884 ;
        RECT 2.260 0.640 2.270 0.874 ;
        RECT 2.270 0.630 2.280 0.864 ;
        RECT 2.280 0.620 2.290 0.854 ;
        RECT 2.290 0.610 2.300 0.844 ;
        RECT 2.300 0.600 2.310 0.834 ;
        RECT 2.310 0.590 2.320 0.824 ;
        RECT 2.320 0.580 2.326 0.820 ;
        RECT 2.115 0.785 2.125 0.955 ;
        RECT 2.125 0.775 2.135 0.955 ;
        RECT 2.135 0.765 2.145 0.955 ;
        RECT 2.145 0.755 2.155 0.955 ;
        RECT 2.155 0.745 2.165 0.955 ;
        RECT 2.165 0.735 2.175 0.955 ;
        RECT 2.175 0.725 2.185 0.955 ;
        RECT 2.185 0.715 2.191 0.955 ;
        RECT 1.580 0.720 1.590 0.954 ;
        RECT 1.590 0.730 1.600 0.954 ;
        RECT 1.600 0.740 1.610 0.954 ;
        RECT 1.610 0.750 1.620 0.954 ;
        RECT 1.620 0.760 1.630 0.954 ;
        RECT 1.630 0.770 1.640 0.954 ;
        RECT 1.640 0.780 1.650 0.954 ;
        RECT 1.650 0.785 1.656 0.955 ;
        RECT 1.505 0.710 1.515 0.880 ;
        RECT 1.515 0.710 1.525 0.890 ;
        RECT 1.525 0.710 1.535 0.900 ;
        RECT 1.535 0.710 1.545 0.910 ;
        RECT 1.545 0.710 1.555 0.920 ;
        RECT 1.555 0.710 1.565 0.930 ;
        RECT 1.565 0.710 1.575 0.940 ;
        RECT 1.575 0.710 1.581 0.950 ;
        RECT 1.050 0.710 1.060 0.954 ;
        RECT 1.060 0.710 1.070 0.944 ;
        RECT 1.070 0.710 1.080 0.934 ;
        RECT 1.080 0.710 1.090 0.924 ;
        RECT 1.090 0.710 1.100 0.914 ;
        RECT 1.100 0.710 1.110 0.904 ;
        RECT 1.110 0.710 1.120 0.894 ;
        RECT 1.120 0.710 1.130 0.884 ;
        RECT 1.130 0.710 1.136 0.880 ;
        RECT 1.030 1.450 1.040 2.364 ;
        RECT 1.040 1.460 1.050 2.364 ;
        RECT 1.050 1.470 1.060 2.364 ;
        RECT 1.060 1.480 1.070 2.364 ;
        RECT 1.070 1.485 1.076 2.365 ;
        RECT 1.030 0.730 1.040 0.974 ;
        RECT 1.040 0.720 1.050 0.964 ;
        RECT 0.905 0.855 0.915 2.365 ;
        RECT 0.915 0.845 0.925 2.365 ;
        RECT 0.925 0.835 0.935 2.365 ;
        RECT 0.935 0.825 0.945 2.365 ;
        RECT 0.945 0.815 0.955 2.365 ;
        RECT 0.955 0.805 0.965 2.365 ;
        RECT 0.965 0.795 0.975 2.365 ;
        RECT 0.975 0.785 0.985 2.365 ;
        RECT 0.985 0.775 0.995 2.365 ;
        RECT 0.995 0.765 1.005 2.365 ;
        RECT 1.005 0.755 1.015 2.365 ;
        RECT 1.015 0.745 1.025 2.365 ;
        RECT 1.025 0.735 1.031 2.365 ;
        RECT 0.860 0.900 0.870 1.514 ;
        RECT 0.870 0.890 0.880 1.524 ;
        RECT 0.880 0.880 0.890 1.534 ;
        RECT 0.890 0.870 0.900 1.544 ;
        RECT 0.900 0.860 0.906 1.554 ;
        RECT 4.020 0.925 4.200 1.225 ;
        RECT 4.030 0.925 4.200 1.775 ;
        RECT 4.050 1.475 4.220 2.145 ;
        RECT 4.030 1.475 4.815 1.775 ;
        RECT 2.445 1.045 2.615 2.495 ;
        RECT 2.610 0.925 2.780 1.225 ;
        RECT 2.445 1.045 2.780 1.225 ;
        RECT 4.400 1.955 4.570 2.495 ;
        RECT 2.445 2.325 4.570 2.495 ;
        RECT 4.995 1.680 5.165 2.125 ;
        RECT 4.400 1.955 5.165 2.125 ;
        RECT 5.240 1.550 5.410 1.850 ;
        RECT 4.995 1.680 5.410 1.850 ;
        RECT 4.465 0.990 5.700 1.160 ;
        RECT 5.530 0.990 5.700 1.345 ;
        RECT 5.355 2.045 5.655 2.215 ;
        RECT 5.355 2.045 5.665 2.205 ;
        RECT 5.355 2.045 5.675 2.195 ;
        RECT 5.355 2.045 5.685 2.185 ;
        RECT 5.355 2.045 5.695 2.175 ;
        RECT 5.355 2.045 5.705 2.165 ;
        RECT 5.355 2.045 5.715 2.155 ;
        RECT 5.355 2.045 5.725 2.145 ;
        RECT 5.355 2.045 5.735 2.135 ;
        RECT 5.355 2.045 5.745 2.125 ;
        RECT 5.355 2.045 5.755 2.115 ;
        RECT 5.590 1.535 5.761 2.109 ;
        RECT 4.095 0.525 6.050 0.695 ;
        RECT 5.880 0.525 6.050 1.705 ;
        RECT 5.590 1.535 6.520 1.705 ;
        RECT 1.210 1.060 1.425 1.360 ;
        RECT 1.255 1.060 1.425 2.715 ;
        RECT 2.095 2.545 2.265 2.845 ;
        RECT 1.255 2.545 2.265 2.715 ;
        RECT 2.325 2.675 2.625 3.085 ;
        RECT 4.750 2.395 4.920 2.845 ;
        RECT 2.095 2.675 4.920 2.845 ;
        RECT 4.750 2.395 5.735 2.565 ;
        RECT 5.910 2.295 6.700 2.465 ;
        RECT 6.875 2.395 7.445 2.565 ;
        RECT 7.275 2.395 7.445 2.770 ;
        RECT 6.800 2.330 6.810 2.564 ;
        RECT 6.810 2.340 6.820 2.564 ;
        RECT 6.820 2.350 6.830 2.564 ;
        RECT 6.830 2.360 6.840 2.564 ;
        RECT 6.840 2.370 6.850 2.564 ;
        RECT 6.850 2.380 6.860 2.564 ;
        RECT 6.860 2.390 6.870 2.564 ;
        RECT 6.870 2.395 6.876 2.565 ;
        RECT 6.775 2.305 6.785 2.539 ;
        RECT 6.785 2.315 6.795 2.549 ;
        RECT 6.795 2.320 6.801 2.560 ;
        RECT 6.700 2.295 6.710 2.465 ;
        RECT 6.710 2.295 6.720 2.475 ;
        RECT 6.720 2.295 6.730 2.485 ;
        RECT 6.730 2.295 6.740 2.495 ;
        RECT 6.740 2.295 6.750 2.505 ;
        RECT 6.750 2.295 6.760 2.515 ;
        RECT 6.760 2.295 6.770 2.525 ;
        RECT 6.770 2.295 6.776 2.535 ;
        RECT 5.835 2.295 5.845 2.529 ;
        RECT 5.845 2.295 5.855 2.519 ;
        RECT 5.855 2.295 5.865 2.509 ;
        RECT 5.865 2.295 5.875 2.499 ;
        RECT 5.875 2.295 5.885 2.489 ;
        RECT 5.885 2.295 5.895 2.479 ;
        RECT 5.895 2.295 5.905 2.469 ;
        RECT 5.905 2.295 5.911 2.465 ;
        RECT 5.810 2.320 5.820 2.554 ;
        RECT 5.820 2.310 5.830 2.544 ;
        RECT 5.830 2.300 5.836 2.540 ;
        RECT 5.735 2.395 5.745 2.565 ;
        RECT 5.745 2.385 5.755 2.565 ;
        RECT 5.755 2.375 5.765 2.565 ;
        RECT 5.765 2.365 5.775 2.565 ;
        RECT 5.775 2.355 5.785 2.565 ;
        RECT 5.785 2.345 5.795 2.565 ;
        RECT 5.795 2.335 5.805 2.565 ;
        RECT 5.805 2.325 5.811 2.565 ;
        RECT 5.100 2.745 5.270 3.210 ;
        RECT 4.395 3.040 5.270 3.210 ;
        RECT 5.100 2.745 5.910 2.915 ;
        RECT 6.085 2.645 6.545 2.815 ;
        RECT 6.720 2.745 7.030 2.915 ;
        RECT 6.860 2.745 7.030 3.120 ;
        RECT 7.335 1.205 7.575 1.375 ;
        RECT 7.625 1.205 7.650 3.120 ;
        RECT 6.860 2.950 7.650 3.120 ;
        RECT 7.650 1.215 7.660 3.119 ;
        RECT 7.660 1.225 7.670 3.119 ;
        RECT 7.670 1.235 7.680 3.119 ;
        RECT 7.680 1.245 7.690 3.119 ;
        RECT 7.690 1.255 7.700 3.119 ;
        RECT 7.700 1.265 7.710 3.119 ;
        RECT 7.710 1.275 7.720 3.119 ;
        RECT 7.720 1.285 7.730 3.119 ;
        RECT 7.730 1.295 7.740 3.119 ;
        RECT 7.740 1.305 7.750 3.119 ;
        RECT 7.750 1.315 7.760 3.119 ;
        RECT 7.760 1.325 7.770 3.119 ;
        RECT 7.770 1.335 7.780 3.119 ;
        RECT 7.780 1.345 7.790 3.119 ;
        RECT 7.790 1.350 7.796 3.120 ;
        RECT 7.575 1.205 7.585 1.375 ;
        RECT 7.585 1.205 7.595 1.385 ;
        RECT 7.595 1.205 7.605 1.395 ;
        RECT 7.605 1.205 7.615 1.405 ;
        RECT 7.615 1.205 7.625 1.415 ;
        RECT 6.645 2.680 6.655 2.914 ;
        RECT 6.655 2.690 6.665 2.914 ;
        RECT 6.665 2.700 6.675 2.914 ;
        RECT 6.675 2.710 6.685 2.914 ;
        RECT 6.685 2.720 6.695 2.914 ;
        RECT 6.695 2.730 6.705 2.914 ;
        RECT 6.705 2.740 6.715 2.914 ;
        RECT 6.715 2.745 6.721 2.915 ;
        RECT 6.620 2.655 6.630 2.889 ;
        RECT 6.630 2.665 6.640 2.899 ;
        RECT 6.640 2.670 6.646 2.910 ;
        RECT 6.545 2.645 6.555 2.815 ;
        RECT 6.555 2.645 6.565 2.825 ;
        RECT 6.565 2.645 6.575 2.835 ;
        RECT 6.575 2.645 6.585 2.845 ;
        RECT 6.585 2.645 6.595 2.855 ;
        RECT 6.595 2.645 6.605 2.865 ;
        RECT 6.605 2.645 6.615 2.875 ;
        RECT 6.615 2.645 6.621 2.885 ;
        RECT 6.010 2.645 6.020 2.879 ;
        RECT 6.020 2.645 6.030 2.869 ;
        RECT 6.030 2.645 6.040 2.859 ;
        RECT 6.040 2.645 6.050 2.849 ;
        RECT 6.050 2.645 6.060 2.839 ;
        RECT 6.060 2.645 6.070 2.829 ;
        RECT 6.070 2.645 6.080 2.819 ;
        RECT 6.080 2.645 6.086 2.815 ;
        RECT 5.985 2.670 5.995 2.904 ;
        RECT 5.995 2.660 6.005 2.894 ;
        RECT 6.005 2.650 6.011 2.890 ;
        RECT 5.910 2.745 5.920 2.915 ;
        RECT 5.920 2.735 5.930 2.915 ;
        RECT 5.930 2.725 5.940 2.915 ;
        RECT 5.940 2.715 5.950 2.915 ;
        RECT 5.950 2.705 5.960 2.915 ;
        RECT 5.960 2.695 5.970 2.915 ;
        RECT 5.970 2.685 5.980 2.915 ;
        RECT 5.980 2.675 5.986 2.915 ;
        RECT 8.570 0.760 8.740 1.280 ;
        RECT 8.440 1.110 8.740 1.280 ;
        RECT 8.570 0.760 9.650 0.930 ;
        RECT 9.480 0.760 9.650 1.280 ;
        RECT 9.480 1.110 9.780 1.280 ;
        RECT 8.325 1.460 8.495 1.760 ;
        RECT 8.325 1.460 9.310 1.630 ;
        RECT 8.960 1.110 9.260 1.630 ;
        RECT 9.140 1.460 9.310 2.425 ;
        RECT 10.155 1.650 10.325 2.425 ;
        RECT 9.140 2.255 10.325 2.425 ;
        RECT 10.495 1.540 10.665 1.840 ;
        RECT 10.155 1.650 10.665 1.840 ;
        RECT 6.965 0.835 7.135 2.215 ;
        RECT 6.965 2.045 7.265 2.215 ;
        RECT 6.965 0.835 7.710 1.005 ;
        RECT 7.965 1.015 8.145 1.185 ;
        RECT 7.975 1.015 8.145 2.110 ;
        RECT 7.975 1.940 8.960 2.110 ;
        RECT 8.790 1.940 8.960 2.795 ;
        RECT 9.200 2.625 9.500 2.955 ;
        RECT 11.195 1.525 11.365 2.795 ;
        RECT 8.790 2.625 11.365 2.795 ;
        RECT 7.890 0.950 7.900 1.184 ;
        RECT 7.900 0.960 7.910 1.184 ;
        RECT 7.910 0.970 7.920 1.184 ;
        RECT 7.920 0.980 7.930 1.184 ;
        RECT 7.930 0.990 7.940 1.184 ;
        RECT 7.940 1.000 7.950 1.184 ;
        RECT 7.950 1.010 7.960 1.184 ;
        RECT 7.960 1.015 7.966 1.185 ;
        RECT 7.785 0.845 7.795 1.079 ;
        RECT 7.795 0.855 7.805 1.089 ;
        RECT 7.805 0.865 7.815 1.099 ;
        RECT 7.815 0.875 7.825 1.109 ;
        RECT 7.825 0.885 7.835 1.119 ;
        RECT 7.835 0.895 7.845 1.129 ;
        RECT 7.845 0.905 7.855 1.139 ;
        RECT 7.855 0.915 7.865 1.149 ;
        RECT 7.865 0.925 7.875 1.159 ;
        RECT 7.875 0.935 7.885 1.169 ;
        RECT 7.885 0.940 7.891 1.180 ;
        RECT 7.710 0.835 7.720 1.005 ;
        RECT 7.720 0.835 7.730 1.015 ;
        RECT 7.730 0.835 7.740 1.025 ;
        RECT 7.740 0.835 7.750 1.035 ;
        RECT 7.750 0.835 7.760 1.045 ;
        RECT 7.760 0.835 7.770 1.055 ;
        RECT 7.770 0.835 7.780 1.065 ;
        RECT 7.780 0.835 7.786 1.075 ;
  END 
END FFDSRHD1XHT

MACRO FFDSHDMXHT
  CLASS  CORE ;
  FOREIGN FFDSHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.430 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.090 1.060 9.330 1.360 ;
        RECT 9.120 1.060 9.330 2.470 ;
        RECT 9.090 1.980 9.330 2.470 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.050 1.060 8.220 1.360 ;
        RECT 8.050 1.190 8.510 1.360 ;
        RECT 8.300 1.190 8.510 2.240 ;
        RECT 7.985 2.070 8.510 2.240 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.560 1.495 1.950 2.050 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.615 -0.300 0.915 0.825 ;
        RECT 1.475 -0.300 1.775 0.800 ;
        RECT 3.375 -0.300 3.675 1.020 ;
        RECT 4.570 -0.300 4.870 0.595 ;
        RECT 6.620 -0.300 6.790 0.720 ;
        RECT 8.505 -0.300 8.805 0.595 ;
        RECT 0.000 -0.300 9.430 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.115 0.755 4.415 0.945 ;
        RECT 5.185 0.605 5.355 0.945 ;
        RECT 4.115 0.775 5.355 0.945 ;
        RECT 5.185 0.605 6.375 0.775 ;
        RECT 6.205 0.605 6.375 1.145 ;
        RECT 7.005 0.920 7.360 1.145 ;
        RECT 7.190 0.540 7.360 1.145 ;
        RECT 6.205 0.975 7.360 1.145 ;
        RECT 7.190 0.540 7.595 0.710 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.615 2.810 0.915 3.990 ;
        RECT 1.440 2.810 1.610 3.990 ;
        RECT 3.395 3.160 3.695 3.990 ;
        RECT 4.570 3.160 4.870 3.990 ;
        RECT 6.575 2.770 6.875 3.990 ;
        RECT 7.215 2.945 7.515 3.990 ;
        RECT 8.505 2.925 8.805 3.990 ;
        RECT 0.000 3.390 9.430 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.490 0.915 2.825 1.130 ;
        RECT 2.490 0.830 2.660 1.130 ;
        RECT 2.610 1.980 2.780 2.280 ;
        RECT 2.655 0.915 2.825 2.215 ;
        RECT 2.610 1.980 2.825 2.215 ;
        RECT 2.655 1.675 3.895 1.845 ;
        RECT 3.115 1.245 4.245 1.415 ;
        RECT 4.075 1.125 4.245 2.215 ;
        RECT 3.945 2.045 4.245 2.215 ;
        RECT 4.075 1.125 5.135 1.295 ;
        RECT 0.170 0.590 0.340 1.295 ;
        RECT 0.170 2.195 0.340 2.900 ;
        RECT 0.170 1.125 0.965 1.295 ;
        RECT 0.170 2.195 0.965 2.365 ;
        RECT 0.795 1.125 0.965 2.630 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 2.460 1.960 2.630 ;
        RECT 1.790 2.460 1.960 2.980 ;
        RECT 1.790 2.810 5.675 2.980 ;
        RECT 1.150 1.060 1.380 1.360 ;
        RECT 1.210 1.060 1.380 2.280 ;
        RECT 1.150 1.980 1.380 2.280 ;
        RECT 1.150 1.060 2.310 1.230 ;
        RECT 2.140 0.480 2.310 2.630 ;
        RECT 2.140 1.685 2.400 1.985 ;
        RECT 2.140 0.480 2.965 0.650 ;
        RECT 5.340 1.645 5.510 2.630 ;
        RECT 5.380 1.245 5.550 1.815 ;
        RECT 5.340 1.645 5.550 1.815 ;
        RECT 2.140 2.460 6.255 2.630 ;
        RECT 6.445 1.325 7.710 1.495 ;
        RECT 7.540 0.890 7.710 2.215 ;
        RECT 7.125 2.045 7.710 2.215 ;
        RECT 7.540 1.540 8.120 1.840 ;
        RECT 5.775 0.955 5.945 2.215 ;
        RECT 5.685 0.955 5.985 1.125 ;
        RECT 5.690 2.045 5.990 2.215 ;
        RECT 6.480 1.675 6.650 2.590 ;
        RECT 5.775 1.675 7.225 1.845 ;
        RECT 8.740 1.540 8.910 2.590 ;
        RECT 6.480 2.420 8.910 2.590 ;
        RECT 8.740 1.540 8.920 1.840 ;
  END 
END FFDSHDMXHT

MACRO FFDQRHD1XHT
  CLASS  CORE ;
  FOREIGN FFDQRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.840 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.500 0.720 9.740 1.360 ;
        RECT 9.530 0.720 9.740 2.960 ;
        RECT 9.500 1.980 9.740 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.600 1.270 1.990 1.865 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.430 1.610 5.885 2.010 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.745 ;
        RECT 1.535 -0.300 1.835 0.740 ;
        RECT 3.435 -0.300 3.735 1.020 ;
        RECT 4.455 -0.300 4.755 0.595 ;
        RECT 5.525 -0.300 5.695 0.810 ;
        RECT 7.465 -0.300 7.765 0.575 ;
        RECT 8.915 -0.300 9.215 1.055 ;
        RECT 0.000 -0.300 9.840 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.010 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 2.810 0.865 3.990 ;
        RECT 1.500 2.810 1.670 3.990 ;
        RECT 3.435 3.195 3.735 3.990 ;
        RECT 5.565 3.195 5.865 3.990 ;
        RECT 7.565 2.810 7.865 3.990 ;
        RECT 8.915 2.975 9.215 3.990 ;
        RECT 0.000 3.390 9.840 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.550 1.190 2.810 1.390 ;
        RECT 2.550 0.830 2.720 1.390 ;
        RECT 2.640 1.190 2.810 2.305 ;
        RECT 2.640 1.675 3.935 1.845 ;
        RECT 3.205 1.245 4.285 1.415 ;
        RECT 4.050 0.775 4.220 1.415 ;
        RECT 4.115 1.245 4.285 2.240 ;
        RECT 4.115 2.070 4.655 2.240 ;
        RECT 4.940 0.480 5.110 0.945 ;
        RECT 4.050 0.775 5.110 0.945 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.190 0.965 2.360 ;
        RECT 0.795 1.125 0.965 2.630 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 2.460 2.020 2.630 ;
        RECT 1.850 2.460 2.020 3.015 ;
        RECT 6.305 2.745 6.605 3.015 ;
        RECT 1.850 2.845 6.605 3.015 ;
        RECT 1.210 0.920 1.400 1.360 ;
        RECT 1.230 0.920 1.400 2.280 ;
        RECT 1.210 1.980 1.400 2.280 ;
        RECT 1.210 0.920 2.370 1.090 ;
        RECT 2.200 0.480 2.370 2.665 ;
        RECT 2.200 1.655 2.460 1.955 ;
        RECT 2.200 0.480 3.025 0.650 ;
        RECT 5.505 2.395 5.675 2.665 ;
        RECT 2.200 2.495 5.675 2.665 ;
        RECT 6.225 1.330 6.395 2.565 ;
        RECT 6.225 1.330 6.525 1.500 ;
        RECT 5.505 2.395 7.120 2.565 ;
        RECT 6.950 2.395 7.120 2.770 ;
        RECT 4.465 1.595 5.210 1.765 ;
        RECT 5.040 1.125 5.210 2.280 ;
        RECT 5.875 0.605 6.045 1.295 ;
        RECT 5.015 1.125 6.045 1.295 ;
        RECT 7.090 0.605 7.260 0.945 ;
        RECT 5.875 0.605 7.260 0.775 ;
        RECT 7.090 0.775 8.735 0.945 ;
        RECT 8.565 0.775 8.735 1.675 ;
        RECT 8.015 1.125 8.385 1.495 ;
        RECT 7.255 1.325 8.385 1.495 ;
        RECT 8.215 1.125 8.385 2.215 ;
        RECT 8.215 2.045 8.785 2.215 ;
        RECT 6.515 0.955 6.875 1.125 ;
        RECT 6.705 0.955 6.875 2.215 ;
        RECT 6.620 2.045 6.920 2.215 ;
        RECT 6.705 1.675 8.035 1.845 ;
        RECT 7.865 1.675 8.035 2.630 ;
        RECT 9.150 1.535 9.320 2.630 ;
        RECT 7.865 2.460 9.320 2.630 ;
  END 
END FFDQRHD1XHT

MACRO FFDRHQHDMXHT
  CLASS  CORE ;
  FOREIGN FFDRHQHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.320 1.060 10.560 1.360 ;
        RECT 10.350 1.060 10.560 2.435 ;
        RECT 10.320 1.980 10.560 2.435 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.420 1.270 2.810 1.970 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.250 1.525 6.705 2.140 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.995 ;
        RECT 2.355 -0.300 2.655 0.740 ;
        RECT 4.255 -0.300 4.555 1.020 ;
        RECT 5.275 -0.300 5.575 0.545 ;
        RECT 6.345 -0.300 6.515 0.810 ;
        RECT 8.285 -0.300 8.585 0.575 ;
        RECT 9.735 -0.300 10.035 1.145 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.830 1.525 1.340 1.950 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.385 2.830 1.685 3.990 ;
        RECT 2.320 2.830 2.490 3.990 ;
        RECT 4.315 3.195 4.615 3.990 ;
        RECT 6.345 3.195 6.645 3.990 ;
        RECT 8.385 2.810 8.685 3.990 ;
        RECT 9.705 2.810 10.005 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.175 1.125 1.785 1.295 ;
        RECT 1.615 1.125 1.785 2.300 ;
        RECT 0.925 2.130 1.785 2.300 ;
        RECT 1.615 1.525 1.850 1.825 ;
        RECT 3.370 1.190 3.630 1.390 ;
        RECT 3.370 0.830 3.540 1.390 ;
        RECT 3.460 1.190 3.630 2.305 ;
        RECT 3.460 1.675 4.755 1.845 ;
        RECT 4.025 1.245 5.105 1.415 ;
        RECT 4.870 0.775 5.040 1.415 ;
        RECT 4.935 1.245 5.105 2.240 ;
        RECT 4.935 2.070 5.535 2.240 ;
        RECT 5.760 0.480 5.930 0.945 ;
        RECT 4.870 0.775 5.930 0.945 ;
        RECT 0.170 1.060 0.340 2.150 ;
        RECT 0.170 1.980 0.610 2.150 ;
        RECT 0.440 1.980 0.610 2.650 ;
        RECT 0.440 2.480 2.840 2.650 ;
        RECT 2.670 2.480 2.840 3.015 ;
        RECT 7.125 2.745 7.295 3.015 ;
        RECT 2.670 2.845 7.295 3.015 ;
        RECT 7.125 2.745 7.425 2.915 ;
        RECT 1.775 0.615 2.175 0.785 ;
        RECT 1.995 0.615 2.175 1.090 ;
        RECT 2.050 0.920 2.220 2.280 ;
        RECT 2.030 1.980 2.220 2.280 ;
        RECT 1.995 0.920 3.190 1.090 ;
        RECT 3.020 0.480 3.190 2.665 ;
        RECT 3.020 1.655 3.280 1.955 ;
        RECT 3.020 0.480 3.845 0.650 ;
        RECT 6.325 2.395 6.495 2.665 ;
        RECT 3.020 2.495 6.495 2.665 ;
        RECT 7.045 1.330 7.215 2.565 ;
        RECT 7.045 1.330 7.345 1.500 ;
        RECT 6.325 2.395 7.940 2.565 ;
        RECT 7.770 2.395 7.940 2.795 ;
        RECT 5.285 1.595 6.030 1.765 ;
        RECT 5.860 1.125 6.030 2.280 ;
        RECT 6.695 0.605 6.865 1.295 ;
        RECT 5.835 1.125 6.865 1.295 ;
        RECT 7.910 0.605 8.080 0.945 ;
        RECT 6.695 0.605 8.080 0.775 ;
        RECT 7.910 0.775 9.555 0.945 ;
        RECT 9.385 0.775 9.555 1.815 ;
        RECT 8.835 1.125 9.205 1.495 ;
        RECT 8.075 1.325 9.205 1.495 ;
        RECT 9.035 1.125 9.205 2.215 ;
        RECT 9.035 2.045 9.605 2.215 ;
        RECT 7.335 0.955 7.695 1.125 ;
        RECT 7.525 0.955 7.695 2.215 ;
        RECT 7.440 2.045 7.740 2.215 ;
        RECT 7.525 1.675 8.855 1.845 ;
        RECT 8.685 1.675 8.855 2.630 ;
        RECT 9.970 1.520 10.140 2.630 ;
        RECT 8.685 2.460 10.140 2.630 ;
  END 
END FFDRHQHDMXHT

MACRO FFDRHQHD3XHT
  CLASS  CORE ;
  FOREIGN FFDRHQHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.170 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 13.790 1.980 13.960 2.960 ;
        RECT 13.790 0.720 14.030 1.405 ;
        RECT 13.790 1.235 15.070 1.405 ;
        RECT 13.790 1.980 15.070 2.150 ;
        RECT 14.830 0.720 15.070 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.940 1.270 3.330 1.980 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.575 1.515 8.240 1.950 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 0.595 ;
        RECT 1.205 -0.300 1.505 0.595 ;
        RECT 2.875 -0.300 3.175 0.740 ;
        RECT 4.775 -0.300 5.075 1.020 ;
        RECT 5.755 -0.300 6.055 0.470 ;
        RECT 6.830 -0.300 7.000 0.535 ;
        RECT 7.955 -0.300 8.255 0.945 ;
        RECT 9.825 -0.300 10.125 0.470 ;
        RECT 11.755 -0.300 12.055 0.575 ;
        RECT 13.205 -0.300 13.505 1.055 ;
        RECT 14.245 -0.300 14.545 1.055 ;
        RECT 0.000 -0.300 15.170 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 1.260 1.525 1.860 1.950 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.475 2.935 0.775 3.990 ;
        RECT 1.895 2.965 2.195 3.990 ;
        RECT 2.930 2.830 3.100 3.990 ;
        RECT 4.775 3.195 5.075 3.990 ;
        RECT 6.855 3.255 7.155 3.990 ;
        RECT 7.985 3.200 8.285 3.990 ;
        RECT 9.855 3.215 10.155 3.990 ;
        RECT 11.855 2.810 12.155 3.990 ;
        RECT 13.205 2.975 13.505 3.990 ;
        RECT 14.310 2.570 14.480 3.990 ;
        RECT 0.000 3.390 15.170 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.755 1.125 2.305 1.295 ;
        RECT 2.135 1.125 2.305 2.300 ;
        RECT 1.445 2.130 2.305 2.300 ;
        RECT 2.135 1.525 2.370 1.825 ;
        RECT 3.890 1.190 4.150 1.390 ;
        RECT 3.890 0.835 4.060 1.390 ;
        RECT 3.980 1.190 4.150 2.305 ;
        RECT 3.980 1.700 5.275 1.870 ;
        RECT 4.545 1.270 5.625 1.440 ;
        RECT 5.360 0.775 5.530 1.440 ;
        RECT 5.455 1.270 5.625 2.240 ;
        RECT 5.455 2.070 6.115 2.240 ;
        RECT 6.305 0.775 6.605 1.070 ;
        RECT 7.225 0.480 7.395 0.945 ;
        RECT 5.360 0.775 7.395 0.945 ;
        RECT 7.225 0.480 7.525 0.650 ;
        RECT 0.655 1.125 1.010 1.295 ;
        RECT 0.840 1.125 1.010 2.650 ;
        RECT 0.840 2.480 3.450 2.650 ;
        RECT 3.280 2.480 3.450 3.015 ;
        RECT 9.145 2.845 9.445 3.180 ;
        RECT 3.280 2.845 10.885 3.015 ;
        RECT 10.715 2.845 10.885 3.195 ;
        RECT 10.715 3.025 11.015 3.195 ;
        RECT 3.540 1.655 3.800 1.955 ;
        RECT 0.170 0.775 0.340 2.460 ;
        RECT 2.360 0.550 2.530 0.945 ;
        RECT 0.170 0.775 2.695 0.945 ;
        RECT 2.570 0.920 2.740 2.280 ;
        RECT 2.510 1.980 2.740 2.280 ;
        RECT 2.515 0.920 3.710 1.090 ;
        RECT 3.540 0.480 3.710 1.955 ;
        RECT 3.630 1.655 3.800 2.665 ;
        RECT 3.540 0.480 4.375 0.650 ;
        RECT 8.585 1.485 8.755 2.665 ;
        RECT 8.585 1.485 8.930 1.785 ;
        RECT 9.775 2.395 9.965 2.665 ;
        RECT 3.630 2.495 9.965 2.665 ;
        RECT 10.535 1.350 10.705 2.565 ;
        RECT 10.515 1.350 10.815 1.520 ;
        RECT 9.775 2.395 11.410 2.565 ;
        RECT 11.240 2.395 11.410 2.795 ;
        RECT 5.830 1.520 7.310 1.690 ;
        RECT 7.140 1.125 7.310 2.315 ;
        RECT 7.140 2.145 7.735 2.315 ;
        RECT 8.505 0.650 8.675 1.295 ;
        RECT 7.140 1.125 8.675 1.295 ;
        RECT 10.335 0.605 10.505 0.820 ;
        RECT 8.505 0.650 10.505 0.820 ;
        RECT 10.335 0.605 11.550 0.775 ;
        RECT 11.380 0.605 11.550 0.945 ;
        RECT 11.380 0.775 13.025 0.945 ;
        RECT 12.855 0.775 13.025 1.760 ;
        RECT 12.305 1.125 12.675 1.495 ;
        RECT 11.545 1.325 12.675 1.495 ;
        RECT 12.505 1.125 12.675 2.215 ;
        RECT 12.505 2.045 13.075 2.215 ;
        RECT 8.875 1.125 9.315 1.295 ;
        RECT 9.145 1.000 9.315 2.315 ;
        RECT 8.935 2.145 9.315 2.315 ;
        RECT 9.145 1.000 11.165 1.170 ;
        RECT 10.805 0.955 11.165 1.170 ;
        RECT 10.995 0.955 11.165 2.215 ;
        RECT 10.910 2.045 11.210 2.215 ;
        RECT 10.995 1.675 12.325 1.845 ;
        RECT 12.155 1.675 12.325 2.630 ;
        RECT 13.315 1.585 13.485 2.630 ;
        RECT 12.155 2.460 13.485 2.630 ;
        RECT 13.315 1.585 14.620 1.755 ;
  END 
END FFDRHQHD3XHT

MACRO FFDRHQHD2XHT
  CLASS  CORE ;
  FOREIGN FFDRHQHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.120 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 12.260 0.720 12.430 1.360 ;
        RECT 12.260 1.980 12.430 2.960 ;
        RECT 12.260 1.190 12.610 1.360 ;
        RECT 12.440 1.190 12.610 2.460 ;
        RECT 12.260 1.980 12.610 2.460 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.420 1.270 2.810 1.995 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.900 1.600 6.610 1.950 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.135 ;
        RECT 2.355 -0.300 2.655 0.740 ;
        RECT 4.255 -0.300 4.555 1.020 ;
        RECT 5.235 -0.300 5.535 0.470 ;
        RECT 6.135 -0.300 6.435 0.470 ;
        RECT 8.295 -0.300 8.595 0.470 ;
        RECT 10.225 -0.300 10.525 0.575 ;
        RECT 11.675 -0.300 11.975 1.055 ;
        RECT 12.780 -0.300 12.950 1.120 ;
        RECT 0.000 -0.300 13.120 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.830 1.525 1.340 1.950 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.375 2.830 1.675 3.990 ;
        RECT 2.410 2.830 2.580 3.990 ;
        RECT 4.255 3.195 4.555 3.990 ;
        RECT 6.095 3.255 6.395 3.990 ;
        RECT 8.395 3.195 8.695 3.990 ;
        RECT 10.325 2.810 10.625 3.990 ;
        RECT 11.675 2.975 11.975 3.990 ;
        RECT 12.780 2.570 12.950 3.990 ;
        RECT 0.000 3.390 13.120 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.175 1.125 1.785 1.295 ;
        RECT 1.615 1.125 1.785 2.300 ;
        RECT 0.925 2.130 1.785 2.300 ;
        RECT 1.615 1.525 1.850 1.825 ;
        RECT 3.370 1.190 3.630 1.390 ;
        RECT 3.370 0.835 3.540 1.390 ;
        RECT 3.460 1.190 3.630 2.305 ;
        RECT 3.460 1.700 4.755 1.870 ;
        RECT 4.025 1.270 5.105 1.440 ;
        RECT 4.840 0.835 5.010 1.440 ;
        RECT 4.935 1.270 5.105 2.240 ;
        RECT 4.935 2.070 5.475 2.240 ;
        RECT 4.840 0.835 6.085 1.005 ;
        RECT 5.785 0.650 6.085 1.070 ;
        RECT 6.615 0.480 6.785 0.820 ;
        RECT 5.785 0.650 6.785 0.820 ;
        RECT 6.615 0.480 7.370 0.650 ;
        RECT 0.170 0.720 0.340 2.150 ;
        RECT 0.170 1.980 0.610 2.150 ;
        RECT 0.440 1.980 0.610 2.650 ;
        RECT 0.440 2.480 2.930 2.650 ;
        RECT 2.760 2.480 2.930 3.015 ;
        RECT 7.465 2.845 7.765 3.180 ;
        RECT 2.760 2.845 9.355 3.015 ;
        RECT 9.185 2.845 9.355 3.195 ;
        RECT 9.185 3.025 9.485 3.195 ;
        RECT 3.020 1.655 3.280 1.955 ;
        RECT 1.775 0.615 2.175 0.785 ;
        RECT 1.995 0.615 2.175 1.090 ;
        RECT 2.050 0.920 2.220 2.280 ;
        RECT 2.030 1.980 2.220 2.280 ;
        RECT 1.995 0.920 3.190 1.090 ;
        RECT 3.020 0.480 3.190 1.955 ;
        RECT 3.110 1.655 3.280 2.665 ;
        RECT 3.020 0.480 3.855 0.650 ;
        RECT 7.560 1.550 7.905 1.720 ;
        RECT 7.735 1.550 7.905 2.665 ;
        RECT 9.005 1.350 9.175 2.665 ;
        RECT 3.110 2.495 9.175 2.665 ;
        RECT 8.985 1.350 9.285 1.520 ;
        RECT 9.005 2.395 9.880 2.565 ;
        RECT 9.710 2.395 9.880 2.795 ;
        RECT 5.285 1.250 5.455 1.735 ;
        RECT 5.285 1.250 6.860 1.420 ;
        RECT 6.555 2.145 6.860 2.315 ;
        RECT 7.615 0.650 7.785 1.000 ;
        RECT 7.200 0.830 7.785 1.000 ;
        RECT 8.805 0.605 8.975 0.820 ;
        RECT 7.615 0.650 8.975 0.820 ;
        RECT 8.805 0.605 10.020 0.775 ;
        RECT 9.850 0.605 10.020 0.945 ;
        RECT 9.850 0.775 11.495 0.945 ;
        RECT 11.325 0.775 11.495 1.670 ;
        RECT 7.105 0.830 7.115 1.084 ;
        RECT 7.115 0.830 7.125 1.074 ;
        RECT 7.125 0.830 7.135 1.064 ;
        RECT 7.135 0.830 7.145 1.054 ;
        RECT 7.145 0.830 7.155 1.044 ;
        RECT 7.155 0.830 7.165 1.034 ;
        RECT 7.165 0.830 7.175 1.024 ;
        RECT 7.175 0.830 7.185 1.014 ;
        RECT 7.185 0.830 7.195 1.004 ;
        RECT 7.195 0.830 7.201 1.000 ;
        RECT 7.030 0.905 7.040 1.159 ;
        RECT 7.040 0.895 7.050 1.149 ;
        RECT 7.050 0.885 7.060 1.139 ;
        RECT 7.060 0.875 7.070 1.129 ;
        RECT 7.070 0.865 7.080 1.119 ;
        RECT 7.080 0.855 7.090 1.109 ;
        RECT 7.090 0.845 7.100 1.099 ;
        RECT 7.100 0.835 7.106 1.095 ;
        RECT 6.860 1.075 6.870 2.315 ;
        RECT 6.870 1.065 6.880 2.315 ;
        RECT 6.880 1.055 6.890 2.315 ;
        RECT 6.890 1.045 6.900 2.315 ;
        RECT 6.900 1.035 6.910 2.315 ;
        RECT 6.910 1.025 6.920 2.315 ;
        RECT 6.920 1.015 6.930 2.315 ;
        RECT 6.930 1.005 6.940 2.315 ;
        RECT 6.940 0.995 6.950 2.315 ;
        RECT 6.950 0.985 6.960 2.315 ;
        RECT 6.960 0.975 6.970 2.315 ;
        RECT 6.970 0.965 6.980 2.315 ;
        RECT 6.980 0.955 6.990 2.315 ;
        RECT 6.990 0.945 7.000 2.315 ;
        RECT 7.000 0.935 7.010 2.315 ;
        RECT 7.010 0.925 7.020 2.315 ;
        RECT 7.020 0.915 7.030 2.315 ;
        RECT 10.775 1.125 11.145 1.495 ;
        RECT 10.015 1.325 11.145 1.495 ;
        RECT 10.975 1.125 11.145 2.215 ;
        RECT 10.975 2.045 11.545 2.215 ;
        RECT 7.270 1.215 7.380 2.315 ;
        RECT 7.260 1.225 8.405 1.350 ;
        RECT 7.280 1.205 7.380 2.315 ;
        RECT 7.250 1.235 8.405 1.350 ;
        RECT 7.290 1.195 7.380 2.315 ;
        RECT 7.240 1.245 8.405 1.350 ;
        RECT 7.300 1.185 7.380 2.315 ;
        RECT 7.230 1.255 8.405 1.350 ;
        RECT 7.210 1.275 7.380 2.315 ;
        RECT 7.210 1.275 7.390 1.404 ;
        RECT 7.210 1.275 7.400 1.394 ;
        RECT 7.210 1.275 7.410 1.384 ;
        RECT 7.210 1.275 7.420 1.374 ;
        RECT 7.210 1.275 7.430 1.364 ;
        RECT 7.210 1.275 7.440 1.354 ;
        RECT 7.210 2.145 7.510 2.315 ;
        RECT 7.305 1.180 8.405 1.350 ;
        RECT 7.220 1.265 8.405 1.350 ;
        RECT 8.235 1.000 8.405 1.350 ;
        RECT 9.275 0.955 9.635 1.170 ;
        RECT 8.235 1.000 9.635 1.170 ;
        RECT 9.465 0.955 9.635 2.215 ;
        RECT 9.380 2.045 9.680 2.215 ;
        RECT 9.465 1.675 10.795 1.845 ;
        RECT 10.625 1.675 10.795 2.630 ;
        RECT 11.910 1.585 12.080 2.630 ;
        RECT 10.625 2.460 12.080 2.630 ;
        RECT 11.910 1.585 12.260 1.755 ;
  END 
END FFDRHQHD2XHT

MACRO FFDSHDLXHT
  CLASS  CORE ;
  FOREIGN FFDSHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.430 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.090 1.060 9.330 1.360 ;
        RECT 9.120 1.060 9.330 2.280 ;
        RECT 9.090 1.980 9.330 2.280 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.050 1.060 8.220 1.360 ;
        RECT 8.050 1.190 8.510 1.360 ;
        RECT 8.300 1.190 8.510 2.240 ;
        RECT 7.985 2.070 8.510 2.240 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.620 1.495 2.010 2.050 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.825 ;
        RECT 1.535 -0.300 1.835 0.805 ;
        RECT 3.435 -0.300 3.735 1.020 ;
        RECT 4.570 -0.300 4.870 0.595 ;
        RECT 6.555 -0.300 6.855 0.655 ;
        RECT 8.505 -0.300 8.805 0.745 ;
        RECT 0.000 -0.300 9.430 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.175 0.755 4.475 0.945 ;
        RECT 5.185 0.605 5.355 0.945 ;
        RECT 4.175 0.775 5.355 0.945 ;
        RECT 5.185 0.605 6.375 0.775 ;
        RECT 6.205 0.605 6.375 1.145 ;
        RECT 7.005 0.920 7.360 1.145 ;
        RECT 7.190 0.540 7.360 1.145 ;
        RECT 6.205 0.975 7.360 1.145 ;
        RECT 7.190 0.540 7.565 0.710 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.575 2.810 0.875 3.990 ;
        RECT 1.495 2.810 1.665 3.990 ;
        RECT 3.425 3.160 3.725 3.990 ;
        RECT 4.570 3.160 4.870 3.990 ;
        RECT 6.575 2.770 6.875 3.990 ;
        RECT 7.155 2.875 7.455 3.990 ;
        RECT 8.505 2.770 8.805 3.990 ;
        RECT 0.000 3.390 9.430 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.550 0.915 2.885 1.130 ;
        RECT 2.550 0.830 2.720 1.130 ;
        RECT 2.715 0.915 2.885 2.280 ;
        RECT 2.660 1.980 2.885 2.280 ;
        RECT 2.715 1.675 3.955 1.845 ;
        RECT 3.175 1.245 4.305 1.415 ;
        RECT 4.135 1.245 4.305 2.215 ;
        RECT 4.005 2.045 4.305 2.215 ;
        RECT 4.140 1.125 5.135 1.295 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.195 0.965 2.365 ;
        RECT 0.795 1.125 0.965 2.630 ;
        RECT 0.795 1.525 1.070 1.825 ;
        RECT 0.795 2.460 2.020 2.630 ;
        RECT 1.850 2.460 2.020 2.980 ;
        RECT 1.850 2.810 5.675 2.980 ;
        RECT 1.190 1.060 1.420 1.360 ;
        RECT 1.250 1.060 1.420 2.280 ;
        RECT 1.210 1.980 1.420 2.280 ;
        RECT 1.190 1.060 2.370 1.230 ;
        RECT 2.200 0.480 2.370 2.630 ;
        RECT 2.200 1.685 2.460 1.985 ;
        RECT 2.200 0.480 3.025 0.650 ;
        RECT 5.340 1.645 5.510 2.630 ;
        RECT 5.380 1.245 5.550 1.815 ;
        RECT 5.340 1.645 5.550 1.815 ;
        RECT 2.200 2.460 6.255 2.630 ;
        RECT 6.415 1.325 7.710 1.495 ;
        RECT 7.540 0.890 7.710 2.215 ;
        RECT 7.155 2.045 7.710 2.215 ;
        RECT 7.540 1.540 8.120 1.840 ;
        RECT 5.775 0.955 5.945 2.215 ;
        RECT 5.685 0.955 5.985 1.125 ;
        RECT 5.690 2.045 5.990 2.215 ;
        RECT 6.480 1.675 6.650 2.590 ;
        RECT 5.775 1.675 7.195 1.845 ;
        RECT 8.740 1.545 8.910 2.590 ;
        RECT 6.480 2.420 8.910 2.590 ;
        RECT 8.740 1.545 8.920 1.845 ;
  END 
END FFDSHDLXHT

MACRO FFDSHD2XHT
  CLASS  CORE ;
  FOREIGN FFDSHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.070 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.210 0.720 10.380 2.960 ;
        RECT 10.210 1.650 10.560 2.015 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.120 0.720 9.340 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.560 1.265 1.950 1.965 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.745 ;
        RECT 1.495 -0.300 1.795 0.735 ;
        RECT 3.395 -0.300 3.695 0.895 ;
        RECT 4.915 -0.300 5.215 0.715 ;
        RECT 7.035 -0.300 7.335 0.740 ;
        RECT 8.585 -0.300 8.885 1.055 ;
        RECT 9.625 -0.300 9.925 1.055 ;
        RECT 10.665 -0.300 10.965 1.055 ;
        RECT 0.000 -0.300 11.070 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.665 1.130 4.835 1.790 ;
        RECT 5.050 0.960 5.230 1.330 ;
        RECT 4.665 1.130 5.230 1.330 ;
        RECT 5.050 0.960 5.565 1.130 ;
        RECT 5.395 0.605 5.565 1.130 ;
        RECT 5.395 0.605 6.725 0.775 ;
        RECT 6.555 0.605 6.725 1.145 ;
        RECT 7.415 0.920 7.960 1.145 ;
        RECT 6.555 0.975 7.960 1.145 ;
        RECT 7.790 0.920 7.960 1.735 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.545 2.810 0.845 3.990 ;
        RECT 1.495 3.095 1.795 3.990 ;
        RECT 3.455 3.095 3.755 3.990 ;
        RECT 4.570 3.095 5.210 3.990 ;
        RECT 6.965 2.790 7.265 3.990 ;
        RECT 8.075 2.790 8.375 3.990 ;
        RECT 8.585 2.975 8.885 3.990 ;
        RECT 9.625 2.975 9.925 3.990 ;
        RECT 10.665 2.295 10.965 3.990 ;
        RECT 0.000 3.390 11.070 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.510 0.915 2.845 1.130 ;
        RECT 2.510 0.830 2.680 1.130 ;
        RECT 2.675 0.915 2.845 2.215 ;
        RECT 2.595 2.045 2.895 2.215 ;
        RECT 2.675 1.675 3.935 1.845 ;
        RECT 3.135 1.245 4.485 1.415 ;
        RECT 4.315 0.725 4.485 2.215 ;
        RECT 4.315 0.725 4.675 0.895 ;
        RECT 5.195 1.610 5.365 2.215 ;
        RECT 4.005 2.045 5.365 2.215 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.195 0.965 2.365 ;
        RECT 0.795 1.125 0.965 2.630 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 2.460 2.055 2.630 ;
        RECT 1.885 2.460 2.055 2.915 ;
        RECT 2.905 2.745 3.205 2.995 ;
        RECT 1.885 2.745 6.010 2.915 ;
        RECT 5.830 2.745 6.010 3.185 ;
        RECT 5.830 3.015 6.450 3.185 ;
        RECT 1.160 0.915 1.380 1.360 ;
        RECT 1.210 0.915 1.380 2.280 ;
        RECT 1.160 1.980 1.380 2.280 ;
        RECT 1.160 0.915 2.330 1.085 ;
        RECT 2.160 0.480 2.330 1.985 ;
        RECT 2.235 1.685 2.405 2.565 ;
        RECT 2.160 1.685 2.420 1.985 ;
        RECT 2.160 0.480 2.995 0.650 ;
        RECT 5.675 1.290 5.845 2.565 ;
        RECT 2.235 2.395 6.540 2.565 ;
        RECT 6.370 2.395 6.540 2.770 ;
        RECT 8.140 1.060 8.310 2.215 ;
        RECT 7.525 2.045 8.310 2.215 ;
        RECT 8.140 1.615 8.940 1.785 ;
        RECT 6.035 0.955 6.335 1.125 ;
        RECT 6.120 0.955 6.335 2.215 ;
        RECT 6.100 2.045 6.400 2.215 ;
        RECT 7.175 1.590 7.345 2.610 ;
        RECT 6.120 1.590 7.545 1.760 ;
        RECT 8.570 2.440 8.815 2.630 ;
        RECT 7.175 2.440 8.815 2.610 ;
        RECT 9.860 1.545 10.030 2.630 ;
        RECT 8.570 2.460 10.030 2.630 ;
  END 
END FFDSHD2XHT

MACRO FFDSHD1XHT
  CLASS  CORE ;
  FOREIGN FFDSHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.430 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.090 0.720 9.330 1.360 ;
        RECT 9.120 0.720 9.330 2.960 ;
        RECT 9.090 1.980 9.330 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.050 0.720 8.220 1.360 ;
        RECT 8.050 1.190 8.510 1.360 ;
        RECT 8.300 1.190 8.510 2.240 ;
        RECT 7.985 2.070 8.510 2.240 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.560 1.495 1.950 2.050 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.745 ;
        RECT 1.475 -0.300 1.775 0.795 ;
        RECT 3.365 -0.300 3.665 1.020 ;
        RECT 4.570 -0.300 4.870 0.595 ;
        RECT 6.620 -0.300 6.790 0.640 ;
        RECT 8.505 -0.300 8.805 0.715 ;
        RECT 0.000 -0.300 9.430 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.105 0.705 4.405 0.945 ;
        RECT 5.185 0.605 5.355 0.945 ;
        RECT 4.105 0.775 5.355 0.945 ;
        RECT 5.185 0.605 6.375 0.775 ;
        RECT 6.205 0.605 6.375 1.145 ;
        RECT 7.005 0.920 7.360 1.145 ;
        RECT 7.190 0.535 7.360 1.145 ;
        RECT 6.205 0.975 7.360 1.145 ;
        RECT 7.190 0.535 7.595 0.705 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 2.810 0.835 3.990 ;
        RECT 1.440 2.810 1.610 3.990 ;
        RECT 3.395 3.160 3.695 3.990 ;
        RECT 4.570 3.160 4.870 3.990 ;
        RECT 6.575 2.770 6.875 3.990 ;
        RECT 7.215 3.005 7.515 3.990 ;
        RECT 8.505 2.975 8.805 3.990 ;
        RECT 0.000 3.390 9.430 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.490 0.915 2.825 1.130 ;
        RECT 2.490 0.830 2.660 1.130 ;
        RECT 2.610 1.980 2.780 2.280 ;
        RECT 2.655 0.915 2.825 2.215 ;
        RECT 2.610 1.980 2.825 2.215 ;
        RECT 2.655 1.675 3.895 1.845 ;
        RECT 3.115 1.245 4.245 1.415 ;
        RECT 4.075 1.125 4.245 2.215 ;
        RECT 3.945 2.045 4.245 2.215 ;
        RECT 4.075 1.125 5.135 1.295 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.195 0.965 2.365 ;
        RECT 0.795 1.125 0.965 2.630 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 2.460 1.960 2.630 ;
        RECT 1.790 2.460 1.960 2.980 ;
        RECT 1.790 2.810 5.675 2.980 ;
        RECT 1.150 1.060 1.380 1.360 ;
        RECT 1.210 1.060 1.380 2.280 ;
        RECT 1.150 1.980 1.380 2.280 ;
        RECT 1.150 1.060 2.310 1.230 ;
        RECT 2.140 0.480 2.310 2.630 ;
        RECT 2.140 1.685 2.400 1.985 ;
        RECT 2.140 0.480 2.965 0.650 ;
        RECT 5.340 1.645 5.510 2.630 ;
        RECT 5.380 1.245 5.550 1.815 ;
        RECT 5.340 1.645 5.550 1.815 ;
        RECT 2.140 2.460 6.190 2.630 ;
        RECT 6.020 2.460 6.190 2.770 ;
        RECT 6.445 1.325 7.710 1.495 ;
        RECT 7.540 0.890 7.710 2.215 ;
        RECT 7.125 2.045 7.710 2.215 ;
        RECT 7.540 1.540 8.120 1.840 ;
        RECT 5.775 0.955 5.945 2.215 ;
        RECT 5.685 0.955 5.985 1.125 ;
        RECT 5.690 2.045 5.990 2.215 ;
        RECT 6.480 1.675 6.650 2.590 ;
        RECT 5.775 1.675 7.225 1.845 ;
        RECT 8.740 1.530 8.910 2.590 ;
        RECT 6.480 2.420 8.910 2.590 ;
        RECT 8.740 1.530 8.920 1.830 ;
  END 
END FFDSHD1XHT

MACRO FFDRHQHD1XHT
  CLASS  CORE ;
  FOREIGN FFDRHQHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.320 0.720 10.560 1.360 ;
        RECT 10.350 0.720 10.560 2.960 ;
        RECT 10.320 1.980 10.560 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.420 1.270 2.810 1.935 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.250 1.515 6.705 2.010 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.995 ;
        RECT 2.355 -0.300 2.655 0.740 ;
        RECT 4.255 -0.300 4.555 1.020 ;
        RECT 5.275 -0.300 5.575 0.545 ;
        RECT 6.345 -0.300 6.515 0.810 ;
        RECT 8.285 -0.300 8.585 0.575 ;
        RECT 9.735 -0.300 10.035 1.055 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.830 1.525 1.340 1.950 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.385 2.830 1.685 3.990 ;
        RECT 2.320 2.830 2.490 3.990 ;
        RECT 4.315 3.195 4.615 3.990 ;
        RECT 6.345 3.195 6.645 3.990 ;
        RECT 8.385 2.810 8.685 3.990 ;
        RECT 9.735 2.975 10.035 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.175 1.125 1.785 1.295 ;
        RECT 1.615 1.125 1.785 2.300 ;
        RECT 0.925 2.130 1.785 2.300 ;
        RECT 1.615 1.525 1.850 1.825 ;
        RECT 3.370 1.190 3.630 1.390 ;
        RECT 3.370 0.835 3.540 1.390 ;
        RECT 3.460 1.190 3.630 2.305 ;
        RECT 3.460 1.675 4.755 1.845 ;
        RECT 4.025 1.245 5.105 1.415 ;
        RECT 4.870 0.775 5.040 1.415 ;
        RECT 4.935 1.245 5.105 2.240 ;
        RECT 4.935 2.070 5.535 2.240 ;
        RECT 5.760 0.480 5.930 0.945 ;
        RECT 4.870 0.775 5.930 0.945 ;
        RECT 0.170 1.060 0.340 2.150 ;
        RECT 0.170 1.980 0.610 2.150 ;
        RECT 0.440 1.980 0.610 2.650 ;
        RECT 0.440 2.480 2.840 2.650 ;
        RECT 2.670 2.480 2.840 3.015 ;
        RECT 2.670 2.845 7.085 3.015 ;
        RECT 6.915 2.845 7.085 3.195 ;
        RECT 6.915 3.025 7.385 3.195 ;
        RECT 1.775 0.615 2.175 0.785 ;
        RECT 1.995 0.615 2.175 1.090 ;
        RECT 2.050 0.920 2.220 2.280 ;
        RECT 2.030 1.980 2.220 2.280 ;
        RECT 1.995 0.920 3.190 1.090 ;
        RECT 3.020 0.480 3.190 2.665 ;
        RECT 3.020 1.655 3.280 1.955 ;
        RECT 3.020 0.480 3.845 0.650 ;
        RECT 6.325 2.395 6.495 2.665 ;
        RECT 3.020 2.495 6.495 2.665 ;
        RECT 7.045 1.330 7.215 2.565 ;
        RECT 7.045 1.330 7.345 1.500 ;
        RECT 6.325 2.395 7.940 2.565 ;
        RECT 7.770 2.395 7.940 2.795 ;
        RECT 5.285 1.595 6.030 1.765 ;
        RECT 5.860 1.125 6.030 2.280 ;
        RECT 6.695 0.605 6.865 1.295 ;
        RECT 5.835 1.125 6.865 1.295 ;
        RECT 7.910 0.605 8.080 0.945 ;
        RECT 6.695 0.605 8.080 0.775 ;
        RECT 7.910 0.775 9.555 0.945 ;
        RECT 9.385 0.775 9.555 1.715 ;
        RECT 8.835 1.125 9.205 1.495 ;
        RECT 8.075 1.325 9.205 1.495 ;
        RECT 9.035 1.125 9.205 2.215 ;
        RECT 9.035 2.045 9.605 2.215 ;
        RECT 7.335 0.955 7.695 1.125 ;
        RECT 7.525 0.955 7.695 2.215 ;
        RECT 7.470 2.045 7.770 2.215 ;
        RECT 7.525 1.675 8.855 1.845 ;
        RECT 8.685 1.675 8.855 2.630 ;
        RECT 9.970 1.515 10.140 2.630 ;
        RECT 8.685 2.460 10.140 2.630 ;
  END 
END FFDRHQHD1XHT

MACRO FFDRHDMXHT
  CLASS  CORE ;
  FOREIGN FFDRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.220 1.060 10.560 1.360 ;
        RECT 10.350 1.060 10.560 2.280 ;
        RECT 10.220 1.980 10.560 2.280 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.120 0.855 9.370 1.470 ;
        RECT 9.120 1.300 9.690 1.470 ;
        RECT 9.520 1.300 9.690 2.215 ;
        RECT 9.115 2.045 9.690 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.640 1.270 2.030 1.815 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.430 1.485 5.925 2.010 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.825 ;
        RECT 1.575 -0.300 1.875 0.740 ;
        RECT 3.505 -0.300 3.805 1.020 ;
        RECT 4.495 -0.300 4.795 0.595 ;
        RECT 5.565 -0.300 5.735 0.810 ;
        RECT 7.505 -0.300 7.805 0.575 ;
        RECT 8.635 -0.300 8.935 0.595 ;
        RECT 9.665 -0.300 9.965 0.595 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.590 2.010 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.635 2.810 0.935 3.990 ;
        RECT 1.540 2.810 1.710 3.990 ;
        RECT 3.535 3.195 3.835 3.990 ;
        RECT 5.605 3.195 5.905 3.990 ;
        RECT 7.605 2.810 7.905 3.990 ;
        RECT 9.605 2.925 9.905 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.590 1.190 2.850 1.390 ;
        RECT 2.590 0.830 2.760 1.390 ;
        RECT 2.680 1.190 2.850 2.305 ;
        RECT 2.680 1.675 3.975 1.845 ;
        RECT 3.245 1.245 4.325 1.415 ;
        RECT 4.120 0.775 4.290 1.415 ;
        RECT 4.155 1.245 4.325 2.215 ;
        RECT 4.155 2.045 4.755 2.215 ;
        RECT 4.980 0.480 5.150 0.945 ;
        RECT 4.120 0.775 5.150 0.945 ;
        RECT 0.105 1.125 1.005 1.295 ;
        RECT 0.105 2.190 1.005 2.360 ;
        RECT 0.835 1.125 1.005 2.630 ;
        RECT 0.835 1.525 1.070 1.825 ;
        RECT 0.835 2.460 2.060 2.630 ;
        RECT 1.890 2.460 2.060 3.015 ;
        RECT 5.900 2.745 6.070 3.015 ;
        RECT 1.890 2.845 6.070 3.015 ;
        RECT 5.900 2.745 6.620 2.915 ;
        RECT 1.250 0.920 1.440 1.360 ;
        RECT 1.270 0.920 1.440 2.280 ;
        RECT 1.250 1.980 1.440 2.280 ;
        RECT 1.250 0.920 2.410 1.090 ;
        RECT 2.240 0.480 2.410 2.665 ;
        RECT 2.240 1.655 2.500 1.955 ;
        RECT 2.240 0.480 3.065 0.650 ;
        RECT 5.545 2.395 5.715 2.665 ;
        RECT 2.240 2.495 5.715 2.665 ;
        RECT 6.285 1.330 6.455 2.565 ;
        RECT 6.265 1.330 6.565 1.500 ;
        RECT 5.545 2.395 7.225 2.565 ;
        RECT 6.925 2.395 7.225 2.595 ;
        RECT 4.505 1.585 5.250 1.755 ;
        RECT 5.080 1.125 5.250 2.280 ;
        RECT 5.915 0.605 6.085 1.295 ;
        RECT 5.055 1.125 6.085 1.295 ;
        RECT 7.130 0.605 7.300 0.945 ;
        RECT 5.915 0.605 7.300 0.775 ;
        RECT 7.130 0.775 8.775 0.945 ;
        RECT 8.605 0.775 8.775 1.515 ;
        RECT 8.055 1.125 8.425 1.495 ;
        RECT 7.295 1.325 8.425 1.495 ;
        RECT 8.255 1.125 8.425 1.865 ;
        RECT 8.590 1.695 8.760 2.280 ;
        RECT 9.040 1.675 9.340 1.865 ;
        RECT 8.255 1.695 9.340 1.865 ;
        RECT 6.555 0.955 6.915 1.125 ;
        RECT 6.745 0.955 6.915 2.215 ;
        RECT 6.660 2.045 6.960 2.215 ;
        RECT 6.745 1.675 8.075 1.845 ;
        RECT 7.905 1.675 8.075 2.630 ;
        RECT 9.870 1.515 10.040 2.630 ;
        RECT 7.905 2.460 10.040 2.630 ;
  END 
END FFDRHDMXHT

MACRO FFDRHDLXHT
  CLASS  CORE ;
  FOREIGN FFDRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.220 1.060 10.560 1.360 ;
        RECT 10.350 1.060 10.560 2.445 ;
        RECT 10.220 1.980 10.560 2.445 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.120 0.855 9.350 1.470 ;
        RECT 9.120 1.300 9.690 1.470 ;
        RECT 9.520 1.300 9.690 2.215 ;
        RECT 9.115 2.045 9.690 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.640 1.270 2.030 1.815 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.430 1.480 5.925 2.010 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.685 -0.300 0.985 0.865 ;
        RECT 1.575 -0.300 1.875 0.740 ;
        RECT 3.505 -0.300 3.805 1.020 ;
        RECT 4.495 -0.300 4.795 0.595 ;
        RECT 5.565 -0.300 5.735 0.810 ;
        RECT 7.505 -0.300 7.805 0.595 ;
        RECT 8.605 -0.300 8.905 0.595 ;
        RECT 9.665 -0.300 9.965 0.745 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.590 2.010 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.635 2.810 0.935 3.990 ;
        RECT 1.540 2.810 1.710 3.990 ;
        RECT 3.565 3.195 3.865 3.990 ;
        RECT 5.605 3.195 5.905 3.990 ;
        RECT 7.605 2.810 7.905 3.990 ;
        RECT 9.605 2.810 9.905 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.590 1.190 2.850 1.390 ;
        RECT 2.590 0.830 2.760 1.390 ;
        RECT 2.680 1.190 2.850 2.305 ;
        RECT 2.680 1.675 3.975 1.845 ;
        RECT 3.245 1.245 4.325 1.415 ;
        RECT 4.150 0.775 4.320 1.415 ;
        RECT 4.155 1.245 4.325 2.215 ;
        RECT 4.155 2.045 4.785 2.215 ;
        RECT 4.980 0.480 5.150 0.945 ;
        RECT 4.150 0.775 5.150 0.945 ;
        RECT 0.105 1.125 1.005 1.295 ;
        RECT 0.105 2.190 1.005 2.360 ;
        RECT 0.835 1.125 1.005 2.630 ;
        RECT 0.835 1.525 1.070 1.825 ;
        RECT 0.835 2.460 2.060 2.630 ;
        RECT 1.890 2.460 2.060 3.015 ;
        RECT 5.900 2.745 6.070 3.015 ;
        RECT 1.890 2.845 6.070 3.015 ;
        RECT 5.900 2.745 6.590 2.915 ;
        RECT 1.250 0.920 1.440 1.360 ;
        RECT 1.270 0.920 1.440 2.280 ;
        RECT 1.250 1.980 1.440 2.280 ;
        RECT 1.250 0.920 2.410 1.090 ;
        RECT 2.240 0.480 2.410 2.665 ;
        RECT 2.240 1.655 2.500 1.955 ;
        RECT 2.240 0.480 3.065 0.650 ;
        RECT 5.545 2.395 5.715 2.665 ;
        RECT 2.240 2.495 5.715 2.665 ;
        RECT 6.285 1.330 6.455 2.565 ;
        RECT 6.265 1.330 6.565 1.500 ;
        RECT 5.545 2.395 7.225 2.565 ;
        RECT 6.925 2.395 7.225 2.585 ;
        RECT 4.505 1.500 5.250 1.800 ;
        RECT 5.080 1.125 5.250 2.280 ;
        RECT 5.915 0.605 6.085 1.295 ;
        RECT 5.055 1.125 6.085 1.295 ;
        RECT 7.130 0.605 7.300 0.945 ;
        RECT 5.915 0.605 7.300 0.775 ;
        RECT 7.130 0.775 8.775 0.945 ;
        RECT 8.605 0.775 8.775 1.515 ;
        RECT 8.055 1.125 8.425 1.495 ;
        RECT 7.295 1.325 8.425 1.495 ;
        RECT 8.255 1.125 8.425 1.865 ;
        RECT 8.590 1.695 8.760 2.280 ;
        RECT 9.040 1.675 9.340 1.865 ;
        RECT 8.255 1.695 9.340 1.865 ;
        RECT 6.555 0.955 6.915 1.125 ;
        RECT 6.745 0.955 6.915 2.215 ;
        RECT 6.660 2.045 6.960 2.215 ;
        RECT 6.745 1.675 8.075 1.845 ;
        RECT 7.905 1.675 8.075 2.630 ;
        RECT 9.870 1.510 10.040 2.630 ;
        RECT 7.905 2.460 10.040 2.630 ;
  END 
END FFDRHDLXHT

MACRO FFDRHD2XHT
  CLASS  CORE ;
  FOREIGN FFDRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.480 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.620 0.720 10.790 2.960 ;
        RECT 10.620 1.605 10.970 2.015 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.530 0.720 9.750 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.580 1.270 1.965 1.805 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.480 1.610 6.070 1.910 ;
        RECT 5.840 1.610 6.070 2.130 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.745 ;
        RECT 1.515 -0.300 1.815 0.785 ;
        RECT 3.435 -0.300 3.735 1.020 ;
        RECT 4.505 -0.300 4.805 0.595 ;
        RECT 5.675 -0.300 5.845 0.780 ;
        RECT 7.510 -0.300 7.810 0.595 ;
        RECT 8.995 -0.300 9.295 1.055 ;
        RECT 10.035 -0.300 10.335 1.055 ;
        RECT 11.075 -0.300 11.375 1.055 ;
        RECT 0.000 -0.300 11.480 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.545 2.810 0.845 3.990 ;
        RECT 1.515 3.140 1.815 3.990 ;
        RECT 3.450 3.140 3.750 3.990 ;
        RECT 5.610 3.095 5.910 3.990 ;
        RECT 7.620 2.910 7.920 3.990 ;
        RECT 8.995 2.975 9.295 3.990 ;
        RECT 10.035 2.975 10.335 3.990 ;
        RECT 11.075 2.295 11.375 3.990 ;
        RECT 0.000 3.390 11.480 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.530 1.190 2.855 1.390 ;
        RECT 2.530 0.885 2.700 1.390 ;
        RECT 2.685 1.190 2.855 2.260 ;
        RECT 2.530 2.090 2.855 2.260 ;
        RECT 2.685 1.675 3.915 1.845 ;
        RECT 3.185 1.245 4.265 1.415 ;
        RECT 4.020 0.735 4.190 1.415 ;
        RECT 4.095 1.245 4.265 2.215 ;
        RECT 4.095 2.045 4.715 2.215 ;
        RECT 4.985 0.480 5.155 0.945 ;
        RECT 4.020 0.775 5.155 0.945 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.220 0.965 2.390 ;
        RECT 0.795 1.125 0.965 2.630 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 2.460 2.000 2.630 ;
        RECT 1.830 2.460 2.000 2.960 ;
        RECT 2.835 2.790 3.135 2.975 ;
        RECT 5.150 2.745 5.320 2.960 ;
        RECT 1.830 2.790 5.320 2.960 ;
        RECT 5.150 2.745 6.480 2.915 ;
        RECT 6.310 2.745 6.480 3.210 ;
        RECT 6.310 3.040 7.140 3.210 ;
        RECT 1.190 1.060 1.380 1.360 ;
        RECT 1.210 1.060 1.380 2.280 ;
        RECT 1.190 1.980 1.380 2.280 ;
        RECT 1.190 2.090 2.350 2.280 ;
        RECT 2.180 0.480 2.350 2.610 ;
        RECT 2.180 1.720 2.505 1.890 ;
        RECT 2.180 0.480 3.005 0.650 ;
        RECT 4.795 2.395 4.965 2.610 ;
        RECT 2.180 2.440 4.965 2.610 ;
        RECT 6.270 1.355 6.440 2.565 ;
        RECT 6.270 1.355 6.570 1.525 ;
        RECT 4.795 2.395 7.165 2.565 ;
        RECT 6.995 2.395 7.165 2.795 ;
        RECT 4.445 1.510 5.300 1.810 ;
        RECT 5.130 1.125 5.300 2.215 ;
        RECT 5.020 2.045 5.320 2.215 ;
        RECT 5.560 0.960 5.730 1.295 ;
        RECT 5.060 1.125 5.730 1.295 ;
        RECT 5.560 0.960 6.195 1.130 ;
        RECT 6.025 0.635 6.195 1.130 ;
        RECT 7.145 0.635 7.315 0.945 ;
        RECT 6.025 0.635 7.315 0.805 ;
        RECT 7.145 0.775 8.780 0.945 ;
        RECT 8.610 0.775 8.780 1.490 ;
        RECT 8.060 1.125 8.430 1.495 ;
        RECT 7.250 1.325 8.430 1.495 ;
        RECT 8.260 1.125 8.430 1.845 ;
        RECT 8.595 1.675 8.765 2.305 ;
        RECT 8.260 1.675 9.350 1.845 ;
        RECT 6.560 0.985 6.965 1.155 ;
        RECT 6.795 0.985 6.965 2.215 ;
        RECT 6.665 2.045 6.965 2.215 ;
        RECT 6.795 1.675 8.080 1.845 ;
        RECT 7.910 1.675 8.080 2.655 ;
        RECT 10.270 1.540 10.440 2.655 ;
        RECT 7.910 2.485 10.440 2.655 ;
  END 
END FFDRHD2XHT

MACRO FFDRHD1XHT
  CLASS  CORE ;
  FOREIGN FFDRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.180 0.720 10.560 1.360 ;
        RECT 10.350 0.720 10.560 2.960 ;
        RECT 10.180 1.980 10.560 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.120 1.300 9.650 1.345 ;
        RECT 9.125 0.720 9.330 1.470 ;
        RECT 9.120 0.720 9.330 1.345 ;
        RECT 9.125 1.300 9.650 1.470 ;
        RECT 9.480 1.300 9.650 2.215 ;
        RECT 9.075 2.045 9.650 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.685 1.270 1.990 1.950 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.430 1.485 5.885 2.010 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.745 ;
        RECT 1.535 -0.300 1.835 0.740 ;
        RECT 3.435 -0.300 3.735 1.020 ;
        RECT 4.455 -0.300 4.755 0.595 ;
        RECT 5.525 -0.300 5.695 0.810 ;
        RECT 7.465 -0.300 7.765 0.525 ;
        RECT 8.565 -0.300 8.865 0.480 ;
        RECT 9.595 -0.300 9.895 1.055 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.010 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 2.810 0.865 3.990 ;
        RECT 1.500 2.810 1.670 3.990 ;
        RECT 3.495 3.195 3.795 3.990 ;
        RECT 5.565 3.195 5.865 3.990 ;
        RECT 7.565 2.810 7.865 3.990 ;
        RECT 9.595 2.975 9.895 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.550 1.190 2.810 1.390 ;
        RECT 2.550 0.830 2.720 1.390 ;
        RECT 2.640 1.190 2.810 2.305 ;
        RECT 2.640 1.675 3.935 1.845 ;
        RECT 3.205 1.245 4.285 1.415 ;
        RECT 4.050 0.775 4.220 1.415 ;
        RECT 4.115 1.245 4.285 2.240 ;
        RECT 4.115 2.070 4.715 2.240 ;
        RECT 4.940 0.480 5.110 0.945 ;
        RECT 4.050 0.775 5.110 0.945 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.190 0.965 2.360 ;
        RECT 0.795 1.125 0.965 2.630 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 2.460 2.020 2.630 ;
        RECT 1.850 2.460 2.020 3.015 ;
        RECT 5.860 2.745 6.030 3.015 ;
        RECT 1.850 2.845 6.030 3.015 ;
        RECT 5.860 2.745 6.605 2.915 ;
        RECT 1.210 0.920 1.400 1.360 ;
        RECT 1.230 0.920 1.400 2.280 ;
        RECT 1.210 1.980 1.400 2.280 ;
        RECT 1.210 0.920 2.370 1.090 ;
        RECT 2.200 0.480 2.370 2.665 ;
        RECT 2.200 1.655 2.460 1.955 ;
        RECT 2.200 0.480 3.025 0.650 ;
        RECT 5.505 2.395 5.675 2.665 ;
        RECT 2.200 2.495 5.675 2.665 ;
        RECT 6.245 1.330 6.415 2.565 ;
        RECT 6.225 1.330 6.525 1.500 ;
        RECT 5.505 2.395 7.120 2.565 ;
        RECT 6.950 2.395 7.120 2.770 ;
        RECT 4.465 1.675 5.210 1.845 ;
        RECT 5.040 1.125 5.210 2.280 ;
        RECT 5.875 0.605 6.045 1.295 ;
        RECT 5.015 1.125 6.045 1.295 ;
        RECT 7.090 0.605 7.260 0.945 ;
        RECT 5.875 0.605 7.260 0.775 ;
        RECT 7.090 0.775 8.735 0.945 ;
        RECT 8.565 0.775 8.735 1.515 ;
        RECT 7.255 1.325 8.385 1.495 ;
        RECT 8.015 1.125 8.315 1.495 ;
        RECT 8.215 1.325 8.385 1.865 ;
        RECT 8.550 1.695 8.720 2.280 ;
        RECT 9.000 1.675 9.300 1.865 ;
        RECT 8.215 1.695 9.300 1.865 ;
        RECT 6.515 0.955 6.875 1.125 ;
        RECT 6.705 0.955 6.875 2.215 ;
        RECT 6.620 2.045 6.920 2.215 ;
        RECT 6.705 1.675 8.035 1.845 ;
        RECT 7.865 1.675 8.035 2.630 ;
        RECT 9.830 1.530 10.000 2.630 ;
        RECT 7.865 2.460 10.000 2.630 ;
  END 
END FFDRHD1XHT

MACRO FFDQSRHDMXHT
  CLASS  CORE ;
  FOREIGN FFDQSRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.070 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.730 1.045 10.970 2.480 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.265 2.070 1.845 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.380 1.410 3.850 2.030 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.505 -0.300 0.675 0.850 ;
        RECT 1.720 -0.300 2.020 0.565 ;
        RECT 3.500 -0.300 3.670 1.225 ;
        RECT 6.230 -0.300 6.400 1.360 ;
        RECT 8.125 -0.300 8.425 0.815 ;
        RECT 10.115 -0.300 10.415 0.730 ;
        RECT 0.000 -0.300 11.070 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.195 1.670 0.725 2.015 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 9.780 1.480 10.150 1.880 ;
        RECT 9.940 1.480 10.150 2.020 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.610 2.665 0.910 3.990 ;
        RECT 1.580 2.600 1.880 3.990 ;
        RECT 3.635 3.025 4.615 3.990 ;
        RECT 6.165 2.995 6.465 3.990 ;
        RECT 8.130 2.345 8.770 3.990 ;
        RECT 10.115 2.835 10.415 3.990 ;
        RECT 0.000 3.390 11.070 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 1.030 1.295 ;
        RECT 0.860 0.710 1.030 1.514 ;
        RECT 0.870 1.485 1.076 1.524 ;
        RECT 0.880 1.485 1.076 1.534 ;
        RECT 0.890 1.485 1.076 1.544 ;
        RECT 0.900 1.485 1.076 1.554 ;
        RECT 0.105 2.195 1.030 2.365 ;
        RECT 0.860 1.450 1.040 1.514 ;
        RECT 0.860 1.460 1.050 1.514 ;
        RECT 0.860 1.470 1.060 1.514 ;
        RECT 0.905 1.480 1.070 2.364 ;
        RECT 1.070 1.485 1.076 2.365 ;
        RECT 0.860 0.710 1.590 0.880 ;
        RECT 1.525 0.745 2.370 0.890 ;
        RECT 1.535 0.745 2.370 0.900 ;
        RECT 1.545 0.745 2.370 0.910 ;
        RECT 1.550 0.710 1.590 0.915 ;
        RECT 0.860 0.720 1.600 0.880 ;
        RECT 0.860 0.730 1.610 0.880 ;
        RECT 1.550 0.745 2.370 0.914 ;
        RECT 0.860 0.740 1.620 0.880 ;
        RECT 2.200 0.575 2.370 0.915 ;
        RECT 1.620 0.745 2.370 0.915 ;
        RECT 2.200 0.575 3.130 0.745 ;
        RECT 2.880 1.840 3.050 2.140 ;
        RECT 2.960 0.575 3.130 2.010 ;
        RECT 2.880 1.840 3.130 2.010 ;
        RECT 4.020 0.925 4.200 1.225 ;
        RECT 4.030 0.925 4.200 1.730 ;
        RECT 4.050 1.430 4.220 2.145 ;
        RECT 4.030 1.430 4.820 1.730 ;
        RECT 2.445 1.410 2.615 2.495 ;
        RECT 2.550 0.925 2.720 1.590 ;
        RECT 2.445 1.410 2.720 1.590 ;
        RECT 4.980 2.305 5.171 2.370 ;
        RECT 4.990 2.295 5.045 2.495 ;
        RECT 4.970 2.315 5.171 2.370 ;
        RECT 2.445 2.325 5.045 2.495 ;
        RECT 2.445 2.325 5.055 2.484 ;
        RECT 2.445 2.325 5.065 2.474 ;
        RECT 2.445 2.325 5.075 2.464 ;
        RECT 2.445 2.325 5.085 2.454 ;
        RECT 2.445 2.325 5.095 2.444 ;
        RECT 2.445 2.325 5.105 2.434 ;
        RECT 2.445 2.325 5.115 2.424 ;
        RECT 2.445 2.325 5.125 2.414 ;
        RECT 2.445 2.325 5.135 2.404 ;
        RECT 2.445 2.325 5.145 2.394 ;
        RECT 2.445 2.325 5.155 2.384 ;
        RECT 2.445 2.325 5.165 2.374 ;
        RECT 5.000 1.680 5.171 2.370 ;
        RECT 5.240 1.550 5.410 1.850 ;
        RECT 5.000 1.680 5.410 1.850 ;
        RECT 4.465 0.990 5.700 1.160 ;
        RECT 5.530 0.990 5.700 1.360 ;
        RECT 4.095 0.490 4.395 0.730 ;
        RECT 5.580 2.035 5.761 2.110 ;
        RECT 5.355 2.045 5.655 2.215 ;
        RECT 5.355 2.045 5.665 2.204 ;
        RECT 5.355 2.045 5.675 2.194 ;
        RECT 5.355 2.045 5.685 2.184 ;
        RECT 5.355 2.045 5.695 2.174 ;
        RECT 5.355 2.045 5.705 2.164 ;
        RECT 5.355 2.045 5.715 2.154 ;
        RECT 5.355 2.045 5.725 2.144 ;
        RECT 5.355 2.045 5.735 2.134 ;
        RECT 5.355 2.045 5.745 2.124 ;
        RECT 5.355 2.045 5.755 2.114 ;
        RECT 5.590 1.600 5.761 2.110 ;
        RECT 4.095 0.560 6.050 0.730 ;
        RECT 5.880 0.560 6.050 1.770 ;
        RECT 5.590 1.600 6.675 1.770 ;
        RECT 1.210 1.060 1.425 1.360 ;
        RECT 1.255 1.060 1.425 2.410 ;
        RECT 1.255 2.240 2.265 2.410 ;
        RECT 2.095 2.240 2.265 2.845 ;
        RECT 2.335 2.675 2.635 2.865 ;
        RECT 2.095 2.675 5.185 2.845 ;
        RECT 5.520 2.395 5.735 2.565 ;
        RECT 5.910 2.295 6.700 2.465 ;
        RECT 6.905 2.425 7.600 2.595 ;
        RECT 7.430 2.425 7.600 2.725 ;
        RECT 6.830 2.360 6.840 2.594 ;
        RECT 6.840 2.370 6.850 2.594 ;
        RECT 6.850 2.380 6.860 2.594 ;
        RECT 6.860 2.390 6.870 2.594 ;
        RECT 6.870 2.400 6.880 2.594 ;
        RECT 6.880 2.410 6.890 2.594 ;
        RECT 6.890 2.420 6.900 2.594 ;
        RECT 6.900 2.425 6.906 2.595 ;
        RECT 6.775 2.305 6.785 2.539 ;
        RECT 6.785 2.315 6.795 2.549 ;
        RECT 6.795 2.325 6.805 2.559 ;
        RECT 6.805 2.335 6.815 2.569 ;
        RECT 6.815 2.345 6.825 2.579 ;
        RECT 6.825 2.350 6.831 2.590 ;
        RECT 6.700 2.295 6.710 2.465 ;
        RECT 6.710 2.295 6.720 2.475 ;
        RECT 6.720 2.295 6.730 2.485 ;
        RECT 6.730 2.295 6.740 2.495 ;
        RECT 6.740 2.295 6.750 2.505 ;
        RECT 6.750 2.295 6.760 2.515 ;
        RECT 6.760 2.295 6.770 2.525 ;
        RECT 6.770 2.295 6.776 2.535 ;
        RECT 5.835 2.295 5.845 2.529 ;
        RECT 5.845 2.295 5.855 2.519 ;
        RECT 5.855 2.295 5.865 2.509 ;
        RECT 5.865 2.295 5.875 2.499 ;
        RECT 5.875 2.295 5.885 2.489 ;
        RECT 5.885 2.295 5.895 2.479 ;
        RECT 5.895 2.295 5.905 2.469 ;
        RECT 5.905 2.295 5.911 2.465 ;
        RECT 5.810 2.320 5.820 2.554 ;
        RECT 5.820 2.310 5.830 2.544 ;
        RECT 5.830 2.300 5.836 2.540 ;
        RECT 5.735 2.395 5.745 2.565 ;
        RECT 5.745 2.385 5.755 2.565 ;
        RECT 5.755 2.375 5.765 2.565 ;
        RECT 5.765 2.365 5.775 2.565 ;
        RECT 5.775 2.355 5.785 2.565 ;
        RECT 5.785 2.345 5.795 2.565 ;
        RECT 5.795 2.335 5.805 2.565 ;
        RECT 5.805 2.325 5.811 2.565 ;
        RECT 5.350 2.395 5.360 2.749 ;
        RECT 5.360 2.395 5.370 2.739 ;
        RECT 5.370 2.395 5.380 2.729 ;
        RECT 5.380 2.395 5.390 2.719 ;
        RECT 5.390 2.395 5.400 2.709 ;
        RECT 5.400 2.395 5.410 2.699 ;
        RECT 5.410 2.395 5.420 2.689 ;
        RECT 5.420 2.395 5.430 2.679 ;
        RECT 5.430 2.395 5.440 2.669 ;
        RECT 5.440 2.395 5.450 2.659 ;
        RECT 5.450 2.395 5.460 2.649 ;
        RECT 5.460 2.395 5.470 2.639 ;
        RECT 5.470 2.395 5.480 2.629 ;
        RECT 5.480 2.395 5.490 2.619 ;
        RECT 5.490 2.395 5.500 2.609 ;
        RECT 5.500 2.395 5.510 2.599 ;
        RECT 5.510 2.395 5.520 2.589 ;
        RECT 5.265 2.595 5.275 2.835 ;
        RECT 5.275 2.585 5.285 2.825 ;
        RECT 5.285 2.575 5.295 2.815 ;
        RECT 5.295 2.565 5.305 2.805 ;
        RECT 5.305 2.555 5.315 2.795 ;
        RECT 5.315 2.545 5.325 2.785 ;
        RECT 5.325 2.535 5.335 2.775 ;
        RECT 5.335 2.525 5.345 2.765 ;
        RECT 5.345 2.515 5.351 2.759 ;
        RECT 5.185 2.675 5.195 2.845 ;
        RECT 5.195 2.665 5.205 2.845 ;
        RECT 5.205 2.655 5.215 2.845 ;
        RECT 5.215 2.645 5.225 2.845 ;
        RECT 5.225 2.635 5.235 2.845 ;
        RECT 5.235 2.625 5.245 2.845 ;
        RECT 5.245 2.615 5.255 2.845 ;
        RECT 5.255 2.605 5.265 2.845 ;
        RECT 5.625 2.745 5.795 3.210 ;
        RECT 4.805 3.040 5.795 3.210 ;
        RECT 5.625 2.745 5.910 2.915 ;
        RECT 6.085 2.645 6.545 2.815 ;
        RECT 6.875 2.805 7.175 3.075 ;
        RECT 6.780 2.805 7.175 2.975 ;
        RECT 7.435 1.220 7.565 1.390 ;
        RECT 6.875 2.905 7.780 3.075 ;
        RECT 7.780 1.910 7.790 3.074 ;
        RECT 7.790 1.920 7.800 3.074 ;
        RECT 7.800 1.930 7.810 3.074 ;
        RECT 7.810 1.940 7.820 3.074 ;
        RECT 7.820 1.950 7.830 3.074 ;
        RECT 7.830 1.960 7.840 3.074 ;
        RECT 7.840 1.970 7.850 3.074 ;
        RECT 7.850 1.980 7.860 3.074 ;
        RECT 7.860 1.990 7.870 3.074 ;
        RECT 7.870 2.000 7.880 3.074 ;
        RECT 7.880 2.010 7.890 3.074 ;
        RECT 7.890 2.020 7.900 3.074 ;
        RECT 7.900 2.030 7.910 3.074 ;
        RECT 7.910 2.040 7.920 3.074 ;
        RECT 7.920 2.050 7.930 3.074 ;
        RECT 7.930 2.060 7.940 3.074 ;
        RECT 7.940 2.070 7.950 3.074 ;
        RECT 7.735 1.865 7.745 2.115 ;
        RECT 7.745 1.875 7.755 2.125 ;
        RECT 7.755 1.885 7.765 2.135 ;
        RECT 7.765 1.895 7.775 2.145 ;
        RECT 7.775 1.900 7.781 2.154 ;
        RECT 7.565 1.220 7.575 1.944 ;
        RECT 7.575 1.220 7.585 1.954 ;
        RECT 7.585 1.220 7.595 1.964 ;
        RECT 7.595 1.220 7.605 1.974 ;
        RECT 7.605 1.220 7.615 1.984 ;
        RECT 7.615 1.220 7.625 1.994 ;
        RECT 7.625 1.220 7.635 2.004 ;
        RECT 7.635 1.220 7.645 2.014 ;
        RECT 7.645 1.220 7.655 2.024 ;
        RECT 7.655 1.220 7.665 2.034 ;
        RECT 7.665 1.220 7.675 2.044 ;
        RECT 7.675 1.220 7.685 2.054 ;
        RECT 7.685 1.220 7.695 2.064 ;
        RECT 7.695 1.220 7.705 2.074 ;
        RECT 7.705 1.220 7.715 2.084 ;
        RECT 7.715 1.220 7.725 2.094 ;
        RECT 7.725 1.220 7.735 2.104 ;
        RECT 6.705 2.740 6.715 2.974 ;
        RECT 6.715 2.750 6.725 2.974 ;
        RECT 6.725 2.760 6.735 2.974 ;
        RECT 6.735 2.770 6.745 2.974 ;
        RECT 6.745 2.780 6.755 2.974 ;
        RECT 6.755 2.790 6.765 2.974 ;
        RECT 6.765 2.800 6.775 2.974 ;
        RECT 6.775 2.805 6.781 2.975 ;
        RECT 6.620 2.655 6.630 2.889 ;
        RECT 6.630 2.665 6.640 2.899 ;
        RECT 6.640 2.675 6.650 2.909 ;
        RECT 6.650 2.685 6.660 2.919 ;
        RECT 6.660 2.695 6.670 2.929 ;
        RECT 6.670 2.705 6.680 2.939 ;
        RECT 6.680 2.715 6.690 2.949 ;
        RECT 6.690 2.725 6.700 2.959 ;
        RECT 6.700 2.730 6.706 2.970 ;
        RECT 6.545 2.645 6.555 2.815 ;
        RECT 6.555 2.645 6.565 2.825 ;
        RECT 6.565 2.645 6.575 2.835 ;
        RECT 6.575 2.645 6.585 2.845 ;
        RECT 6.585 2.645 6.595 2.855 ;
        RECT 6.595 2.645 6.605 2.865 ;
        RECT 6.605 2.645 6.615 2.875 ;
        RECT 6.615 2.645 6.621 2.885 ;
        RECT 6.010 2.645 6.020 2.879 ;
        RECT 6.020 2.645 6.030 2.869 ;
        RECT 6.030 2.645 6.040 2.859 ;
        RECT 6.040 2.645 6.050 2.849 ;
        RECT 6.050 2.645 6.060 2.839 ;
        RECT 6.060 2.645 6.070 2.829 ;
        RECT 6.070 2.645 6.080 2.819 ;
        RECT 6.080 2.645 6.086 2.815 ;
        RECT 5.985 2.670 5.995 2.904 ;
        RECT 5.995 2.660 6.005 2.894 ;
        RECT 6.005 2.650 6.011 2.890 ;
        RECT 5.910 2.745 5.920 2.915 ;
        RECT 5.920 2.735 5.930 2.915 ;
        RECT 5.930 2.725 5.940 2.915 ;
        RECT 5.940 2.715 5.950 2.915 ;
        RECT 5.950 2.705 5.960 2.915 ;
        RECT 5.960 2.695 5.970 2.915 ;
        RECT 5.970 2.685 5.980 2.915 ;
        RECT 5.980 2.675 5.986 2.915 ;
        RECT 8.420 1.460 8.590 1.760 ;
        RECT 8.420 1.460 9.520 1.630 ;
        RECT 9.080 1.110 9.380 1.630 ;
        RECT 9.350 1.460 9.520 2.305 ;
        RECT 9.350 2.135 9.800 2.305 ;
        RECT 8.690 0.760 8.860 1.280 ;
        RECT 8.560 1.110 8.860 1.280 ;
        RECT 8.690 0.760 9.770 0.930 ;
        RECT 9.600 0.760 9.770 1.280 ;
        RECT 9.600 1.110 9.900 1.280 ;
        RECT 7.010 0.850 7.180 2.245 ;
        RECT 7.010 2.075 7.385 2.245 ;
        RECT 7.010 0.850 7.825 1.020 ;
        RECT 8.400 1.995 9.135 2.165 ;
        RECT 8.965 1.995 9.135 2.655 ;
        RECT 9.320 2.485 9.620 2.900 ;
        RECT 10.380 1.550 10.550 2.655 ;
        RECT 8.965 2.485 10.550 2.655 ;
        RECT 8.315 1.920 8.325 2.164 ;
        RECT 8.325 1.930 8.335 2.164 ;
        RECT 8.335 1.940 8.345 2.164 ;
        RECT 8.345 1.950 8.355 2.164 ;
        RECT 8.355 1.960 8.365 2.164 ;
        RECT 8.365 1.970 8.375 2.164 ;
        RECT 8.375 1.980 8.385 2.164 ;
        RECT 8.385 1.990 8.395 2.164 ;
        RECT 8.395 1.995 8.401 2.165 ;
        RECT 8.150 1.755 8.160 1.999 ;
        RECT 8.160 1.765 8.170 2.009 ;
        RECT 8.170 1.775 8.180 2.019 ;
        RECT 8.180 1.785 8.190 2.029 ;
        RECT 8.190 1.795 8.200 2.039 ;
        RECT 8.200 1.805 8.210 2.049 ;
        RECT 8.210 1.815 8.220 2.059 ;
        RECT 8.220 1.825 8.230 2.069 ;
        RECT 8.230 1.835 8.240 2.079 ;
        RECT 8.240 1.845 8.250 2.089 ;
        RECT 8.250 1.855 8.260 2.099 ;
        RECT 8.260 1.865 8.270 2.109 ;
        RECT 8.270 1.875 8.280 2.119 ;
        RECT 8.280 1.885 8.290 2.129 ;
        RECT 8.290 1.895 8.300 2.139 ;
        RECT 8.300 1.905 8.310 2.149 ;
        RECT 8.310 1.910 8.316 2.160 ;
        RECT 7.980 0.940 7.990 1.830 ;
        RECT 7.990 0.950 8.000 1.840 ;
        RECT 8.000 0.960 8.010 1.850 ;
        RECT 8.010 0.970 8.020 1.860 ;
        RECT 8.020 0.980 8.030 1.870 ;
        RECT 8.030 0.990 8.040 1.880 ;
        RECT 8.040 1.000 8.050 1.890 ;
        RECT 8.050 1.010 8.060 1.900 ;
        RECT 8.060 1.020 8.070 1.910 ;
        RECT 8.070 1.030 8.080 1.920 ;
        RECT 8.080 1.040 8.090 1.930 ;
        RECT 8.090 1.050 8.100 1.940 ;
        RECT 8.100 1.060 8.110 1.950 ;
        RECT 8.110 1.070 8.120 1.960 ;
        RECT 8.120 1.080 8.130 1.970 ;
        RECT 8.130 1.090 8.140 1.980 ;
        RECT 8.140 1.100 8.150 1.990 ;
        RECT 7.900 0.860 7.910 1.094 ;
        RECT 7.910 0.870 7.920 1.104 ;
        RECT 7.920 0.880 7.930 1.114 ;
        RECT 7.930 0.890 7.940 1.124 ;
        RECT 7.940 0.900 7.950 1.134 ;
        RECT 7.950 0.910 7.960 1.144 ;
        RECT 7.960 0.920 7.970 1.154 ;
        RECT 7.970 0.930 7.980 1.164 ;
        RECT 7.825 0.850 7.835 1.020 ;
        RECT 7.835 0.850 7.845 1.030 ;
        RECT 7.845 0.850 7.855 1.040 ;
        RECT 7.855 0.850 7.865 1.050 ;
        RECT 7.865 0.850 7.875 1.060 ;
        RECT 7.875 0.850 7.885 1.070 ;
        RECT 7.885 0.850 7.895 1.080 ;
        RECT 7.895 0.850 7.901 1.090 ;
  END 
END FFDQSRHDMXHT

MACRO FFDQSRHDLXHT
  CLASS  CORE ;
  FOREIGN FFDQSRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.070 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.730 1.045 10.970 2.470 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.265 2.095 1.880 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.380 1.410 3.860 2.030 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.505 -0.300 0.675 0.850 ;
        RECT 1.735 -0.300 2.035 0.565 ;
        RECT 3.520 -0.300 3.690 1.225 ;
        RECT 6.290 -0.300 6.460 0.930 ;
        RECT 8.155 -0.300 8.455 0.780 ;
        RECT 10.180 -0.300 10.350 0.875 ;
        RECT 0.000 -0.300 11.070 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.185 1.670 0.725 2.015 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 9.830 1.375 10.150 1.870 ;
        RECT 9.940 1.375 10.150 2.020 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.630 2.625 0.930 3.990 ;
        RECT 1.585 2.555 1.885 3.990 ;
        RECT 3.635 3.025 4.615 3.990 ;
        RECT 6.165 2.995 6.465 3.990 ;
        RECT 8.130 2.345 8.770 3.990 ;
        RECT 10.115 2.835 10.415 3.990 ;
        RECT 0.000 3.390 11.070 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 1.030 1.295 ;
        RECT 0.860 0.710 1.030 1.514 ;
        RECT 0.870 1.485 1.076 1.524 ;
        RECT 0.880 1.485 1.076 1.534 ;
        RECT 0.890 1.485 1.076 1.544 ;
        RECT 0.900 1.485 1.076 1.554 ;
        RECT 0.105 2.195 1.030 2.365 ;
        RECT 0.860 1.450 1.040 1.514 ;
        RECT 0.860 1.460 1.050 1.514 ;
        RECT 0.860 1.470 1.060 1.514 ;
        RECT 0.905 1.480 1.070 2.364 ;
        RECT 1.070 1.485 1.076 2.365 ;
        RECT 0.860 0.710 1.590 0.880 ;
        RECT 1.525 0.745 2.385 0.890 ;
        RECT 1.535 0.745 2.385 0.900 ;
        RECT 1.545 0.745 2.385 0.910 ;
        RECT 1.550 0.710 1.590 0.915 ;
        RECT 0.860 0.720 1.600 0.880 ;
        RECT 0.860 0.730 1.610 0.880 ;
        RECT 1.550 0.745 2.385 0.914 ;
        RECT 0.860 0.740 1.620 0.880 ;
        RECT 2.215 0.575 2.385 0.915 ;
        RECT 1.620 0.745 2.385 0.915 ;
        RECT 2.215 0.575 3.130 0.745 ;
        RECT 2.880 1.840 3.050 2.140 ;
        RECT 2.960 0.575 3.130 2.010 ;
        RECT 2.880 1.840 3.130 2.010 ;
        RECT 4.040 0.925 4.210 1.730 ;
        RECT 4.050 1.430 4.220 2.145 ;
        RECT 4.040 1.430 4.805 1.730 ;
        RECT 2.445 1.410 2.615 2.495 ;
        RECT 2.570 0.925 2.740 1.590 ;
        RECT 2.445 1.410 2.740 1.590 ;
        RECT 4.975 2.305 5.050 2.495 ;
        RECT 4.965 2.315 5.156 2.390 ;
        RECT 2.445 2.325 5.050 2.495 ;
        RECT 2.445 2.325 5.060 2.484 ;
        RECT 2.445 2.325 5.070 2.474 ;
        RECT 2.445 2.325 5.080 2.464 ;
        RECT 2.445 2.325 5.090 2.454 ;
        RECT 2.445 2.325 5.100 2.444 ;
        RECT 2.445 2.325 5.110 2.434 ;
        RECT 2.445 2.325 5.120 2.424 ;
        RECT 2.445 2.325 5.130 2.414 ;
        RECT 2.445 2.325 5.140 2.404 ;
        RECT 2.445 2.325 5.150 2.394 ;
        RECT 4.985 1.680 5.156 2.390 ;
        RECT 5.240 1.550 5.410 1.850 ;
        RECT 4.985 1.680 5.410 1.850 ;
        RECT 4.485 0.990 5.760 1.160 ;
        RECT 5.590 0.990 5.760 1.360 ;
        RECT 4.120 0.505 4.420 0.745 ;
        RECT 5.580 2.035 5.761 2.110 ;
        RECT 5.355 2.045 5.655 2.215 ;
        RECT 5.355 2.045 5.665 2.204 ;
        RECT 5.355 2.045 5.675 2.194 ;
        RECT 5.355 2.045 5.685 2.184 ;
        RECT 5.355 2.045 5.695 2.174 ;
        RECT 5.355 2.045 5.705 2.164 ;
        RECT 5.355 2.045 5.715 2.154 ;
        RECT 5.355 2.045 5.725 2.144 ;
        RECT 5.355 2.045 5.735 2.134 ;
        RECT 5.355 2.045 5.745 2.124 ;
        RECT 5.355 2.045 5.755 2.114 ;
        RECT 5.590 1.600 5.761 2.110 ;
        RECT 4.120 0.575 6.110 0.745 ;
        RECT 5.940 0.575 6.110 1.770 ;
        RECT 5.590 1.600 6.665 1.770 ;
        RECT 1.210 1.060 1.425 1.360 ;
        RECT 1.255 1.060 1.425 2.365 ;
        RECT 1.255 2.195 2.265 2.365 ;
        RECT 2.095 2.195 2.265 2.845 ;
        RECT 2.325 2.675 2.625 2.915 ;
        RECT 2.095 2.675 5.195 2.845 ;
        RECT 5.505 2.395 5.735 2.565 ;
        RECT 5.910 2.295 6.700 2.465 ;
        RECT 6.905 2.425 7.600 2.595 ;
        RECT 7.430 2.425 7.600 2.730 ;
        RECT 6.830 2.360 6.840 2.594 ;
        RECT 6.840 2.370 6.850 2.594 ;
        RECT 6.850 2.380 6.860 2.594 ;
        RECT 6.860 2.390 6.870 2.594 ;
        RECT 6.870 2.400 6.880 2.594 ;
        RECT 6.880 2.410 6.890 2.594 ;
        RECT 6.890 2.420 6.900 2.594 ;
        RECT 6.900 2.425 6.906 2.595 ;
        RECT 6.775 2.305 6.785 2.539 ;
        RECT 6.785 2.315 6.795 2.549 ;
        RECT 6.795 2.325 6.805 2.559 ;
        RECT 6.805 2.335 6.815 2.569 ;
        RECT 6.815 2.345 6.825 2.579 ;
        RECT 6.825 2.350 6.831 2.590 ;
        RECT 6.700 2.295 6.710 2.465 ;
        RECT 6.710 2.295 6.720 2.475 ;
        RECT 6.720 2.295 6.730 2.485 ;
        RECT 6.730 2.295 6.740 2.495 ;
        RECT 6.740 2.295 6.750 2.505 ;
        RECT 6.750 2.295 6.760 2.515 ;
        RECT 6.760 2.295 6.770 2.525 ;
        RECT 6.770 2.295 6.776 2.535 ;
        RECT 5.835 2.295 5.845 2.529 ;
        RECT 5.845 2.295 5.855 2.519 ;
        RECT 5.855 2.295 5.865 2.509 ;
        RECT 5.865 2.295 5.875 2.499 ;
        RECT 5.875 2.295 5.885 2.489 ;
        RECT 5.885 2.295 5.895 2.479 ;
        RECT 5.895 2.295 5.905 2.469 ;
        RECT 5.905 2.295 5.911 2.465 ;
        RECT 5.810 2.320 5.820 2.554 ;
        RECT 5.820 2.310 5.830 2.544 ;
        RECT 5.830 2.300 5.836 2.540 ;
        RECT 5.735 2.395 5.745 2.565 ;
        RECT 5.745 2.385 5.755 2.565 ;
        RECT 5.755 2.375 5.765 2.565 ;
        RECT 5.765 2.365 5.775 2.565 ;
        RECT 5.775 2.355 5.785 2.565 ;
        RECT 5.785 2.345 5.795 2.565 ;
        RECT 5.795 2.335 5.805 2.565 ;
        RECT 5.805 2.325 5.811 2.565 ;
        RECT 5.335 2.395 5.345 2.769 ;
        RECT 5.345 2.395 5.355 2.759 ;
        RECT 5.355 2.395 5.365 2.749 ;
        RECT 5.365 2.395 5.375 2.739 ;
        RECT 5.375 2.395 5.385 2.729 ;
        RECT 5.385 2.395 5.395 2.719 ;
        RECT 5.395 2.395 5.405 2.709 ;
        RECT 5.405 2.395 5.415 2.699 ;
        RECT 5.415 2.395 5.425 2.689 ;
        RECT 5.425 2.395 5.435 2.679 ;
        RECT 5.435 2.395 5.445 2.669 ;
        RECT 5.445 2.395 5.455 2.659 ;
        RECT 5.455 2.395 5.465 2.649 ;
        RECT 5.465 2.395 5.475 2.639 ;
        RECT 5.475 2.395 5.485 2.629 ;
        RECT 5.485 2.395 5.495 2.619 ;
        RECT 5.495 2.395 5.505 2.609 ;
        RECT 5.270 2.600 5.280 2.834 ;
        RECT 5.280 2.590 5.290 2.824 ;
        RECT 5.290 2.580 5.300 2.814 ;
        RECT 5.300 2.570 5.310 2.804 ;
        RECT 5.310 2.560 5.320 2.794 ;
        RECT 5.320 2.550 5.330 2.784 ;
        RECT 5.330 2.540 5.336 2.780 ;
        RECT 5.195 2.675 5.205 2.845 ;
        RECT 5.205 2.665 5.215 2.845 ;
        RECT 5.215 2.655 5.225 2.845 ;
        RECT 5.225 2.645 5.235 2.845 ;
        RECT 5.235 2.635 5.245 2.845 ;
        RECT 5.245 2.625 5.255 2.845 ;
        RECT 5.255 2.615 5.265 2.845 ;
        RECT 5.265 2.605 5.271 2.845 ;
        RECT 5.625 2.745 5.795 3.210 ;
        RECT 4.805 3.040 5.795 3.210 ;
        RECT 5.625 2.745 5.910 2.915 ;
        RECT 6.085 2.645 6.545 2.815 ;
        RECT 7.005 2.805 7.175 3.080 ;
        RECT 6.780 2.805 7.175 2.975 ;
        RECT 7.435 1.220 7.605 1.390 ;
        RECT 7.005 2.910 7.780 3.080 ;
        RECT 7.780 1.315 7.790 3.079 ;
        RECT 7.790 1.325 7.800 3.079 ;
        RECT 7.800 1.335 7.810 3.079 ;
        RECT 7.810 1.345 7.820 3.079 ;
        RECT 7.820 1.355 7.830 3.079 ;
        RECT 7.830 1.365 7.840 3.079 ;
        RECT 7.840 1.375 7.850 3.079 ;
        RECT 7.850 1.385 7.860 3.079 ;
        RECT 7.860 1.395 7.870 3.079 ;
        RECT 7.870 1.405 7.880 3.079 ;
        RECT 7.880 1.415 7.890 3.079 ;
        RECT 7.890 1.425 7.900 3.079 ;
        RECT 7.900 1.435 7.910 3.079 ;
        RECT 7.910 1.445 7.920 3.079 ;
        RECT 7.920 1.455 7.930 3.079 ;
        RECT 7.930 1.465 7.940 3.079 ;
        RECT 7.940 1.475 7.950 3.079 ;
        RECT 7.735 1.270 7.745 1.520 ;
        RECT 7.745 1.280 7.755 1.530 ;
        RECT 7.755 1.290 7.765 1.540 ;
        RECT 7.765 1.300 7.775 1.550 ;
        RECT 7.775 1.305 7.781 1.559 ;
        RECT 7.605 1.220 7.615 1.390 ;
        RECT 7.615 1.220 7.625 1.400 ;
        RECT 7.625 1.220 7.635 1.410 ;
        RECT 7.635 1.220 7.645 1.420 ;
        RECT 7.645 1.220 7.655 1.430 ;
        RECT 7.655 1.220 7.665 1.440 ;
        RECT 7.665 1.220 7.675 1.450 ;
        RECT 7.675 1.220 7.685 1.460 ;
        RECT 7.685 1.220 7.695 1.470 ;
        RECT 7.695 1.220 7.705 1.480 ;
        RECT 7.705 1.220 7.715 1.490 ;
        RECT 7.715 1.220 7.725 1.500 ;
        RECT 7.725 1.220 7.735 1.510 ;
        RECT 6.705 2.740 6.715 2.974 ;
        RECT 6.715 2.750 6.725 2.974 ;
        RECT 6.725 2.760 6.735 2.974 ;
        RECT 6.735 2.770 6.745 2.974 ;
        RECT 6.745 2.780 6.755 2.974 ;
        RECT 6.755 2.790 6.765 2.974 ;
        RECT 6.765 2.800 6.775 2.974 ;
        RECT 6.775 2.805 6.781 2.975 ;
        RECT 6.620 2.655 6.630 2.889 ;
        RECT 6.630 2.665 6.640 2.899 ;
        RECT 6.640 2.675 6.650 2.909 ;
        RECT 6.650 2.685 6.660 2.919 ;
        RECT 6.660 2.695 6.670 2.929 ;
        RECT 6.670 2.705 6.680 2.939 ;
        RECT 6.680 2.715 6.690 2.949 ;
        RECT 6.690 2.725 6.700 2.959 ;
        RECT 6.700 2.730 6.706 2.970 ;
        RECT 6.545 2.645 6.555 2.815 ;
        RECT 6.555 2.645 6.565 2.825 ;
        RECT 6.565 2.645 6.575 2.835 ;
        RECT 6.575 2.645 6.585 2.845 ;
        RECT 6.585 2.645 6.595 2.855 ;
        RECT 6.595 2.645 6.605 2.865 ;
        RECT 6.605 2.645 6.615 2.875 ;
        RECT 6.615 2.645 6.621 2.885 ;
        RECT 6.010 2.645 6.020 2.879 ;
        RECT 6.020 2.645 6.030 2.869 ;
        RECT 6.030 2.645 6.040 2.859 ;
        RECT 6.040 2.645 6.050 2.849 ;
        RECT 6.050 2.645 6.060 2.839 ;
        RECT 6.060 2.645 6.070 2.829 ;
        RECT 6.070 2.645 6.080 2.819 ;
        RECT 6.080 2.645 6.086 2.815 ;
        RECT 5.985 2.670 5.995 2.904 ;
        RECT 5.995 2.660 6.005 2.894 ;
        RECT 6.005 2.650 6.011 2.890 ;
        RECT 5.910 2.745 5.920 2.915 ;
        RECT 5.920 2.735 5.930 2.915 ;
        RECT 5.930 2.725 5.940 2.915 ;
        RECT 5.940 2.715 5.950 2.915 ;
        RECT 5.950 2.705 5.960 2.915 ;
        RECT 5.960 2.695 5.970 2.915 ;
        RECT 5.970 2.685 5.980 2.915 ;
        RECT 5.980 2.675 5.986 2.915 ;
        RECT 8.485 1.460 8.655 1.760 ;
        RECT 8.485 1.460 9.520 1.630 ;
        RECT 9.140 1.110 9.440 1.630 ;
        RECT 9.350 1.460 9.520 2.305 ;
        RECT 9.350 2.135 9.800 2.305 ;
        RECT 8.690 0.760 8.860 1.280 ;
        RECT 8.560 1.110 8.860 1.280 ;
        RECT 9.600 0.640 9.900 0.930 ;
        RECT 8.690 0.760 9.900 0.930 ;
        RECT 7.010 0.850 7.180 2.245 ;
        RECT 7.010 2.075 7.355 2.245 ;
        RECT 7.010 0.850 7.795 1.020 ;
        RECT 8.400 1.995 9.135 2.165 ;
        RECT 8.965 1.995 9.135 2.655 ;
        RECT 9.320 2.485 9.620 2.735 ;
        RECT 10.380 1.550 10.550 2.655 ;
        RECT 8.965 2.485 10.550 2.655 ;
        RECT 8.315 1.920 8.325 2.164 ;
        RECT 8.325 1.930 8.335 2.164 ;
        RECT 8.335 1.940 8.345 2.164 ;
        RECT 8.345 1.950 8.355 2.164 ;
        RECT 8.355 1.960 8.365 2.164 ;
        RECT 8.365 1.970 8.375 2.164 ;
        RECT 8.375 1.980 8.385 2.164 ;
        RECT 8.385 1.990 8.395 2.164 ;
        RECT 8.395 1.995 8.401 2.165 ;
        RECT 8.305 1.910 8.315 2.154 ;
        RECT 8.135 1.125 8.145 1.985 ;
        RECT 8.145 1.135 8.155 1.995 ;
        RECT 8.155 1.145 8.165 2.005 ;
        RECT 8.165 1.155 8.175 2.015 ;
        RECT 8.175 1.165 8.185 2.025 ;
        RECT 8.185 1.175 8.195 2.035 ;
        RECT 8.195 1.185 8.205 2.045 ;
        RECT 8.205 1.195 8.215 2.055 ;
        RECT 8.215 1.205 8.225 2.065 ;
        RECT 8.225 1.215 8.235 2.075 ;
        RECT 8.235 1.225 8.245 2.085 ;
        RECT 8.245 1.235 8.255 2.095 ;
        RECT 8.255 1.245 8.265 2.105 ;
        RECT 8.265 1.255 8.275 2.115 ;
        RECT 8.275 1.265 8.285 2.125 ;
        RECT 8.285 1.275 8.295 2.135 ;
        RECT 8.295 1.285 8.305 2.145 ;
        RECT 7.870 0.860 7.880 1.094 ;
        RECT 7.880 0.870 7.890 1.104 ;
        RECT 7.890 0.880 7.900 1.114 ;
        RECT 7.900 0.890 7.910 1.124 ;
        RECT 7.910 0.900 7.920 1.134 ;
        RECT 7.920 0.910 7.930 1.144 ;
        RECT 7.930 0.920 7.940 1.154 ;
        RECT 7.940 0.930 7.950 1.164 ;
        RECT 7.950 0.940 7.960 1.174 ;
        RECT 7.960 0.950 7.970 1.184 ;
        RECT 7.970 0.960 7.980 1.194 ;
        RECT 7.980 0.970 7.990 1.204 ;
        RECT 7.990 0.980 8.000 1.214 ;
        RECT 8.000 0.990 8.010 1.224 ;
        RECT 8.010 1.000 8.020 1.234 ;
        RECT 8.020 1.010 8.030 1.244 ;
        RECT 8.030 1.020 8.040 1.254 ;
        RECT 8.040 1.030 8.050 1.264 ;
        RECT 8.050 1.040 8.060 1.274 ;
        RECT 8.060 1.050 8.070 1.284 ;
        RECT 8.070 1.060 8.080 1.294 ;
        RECT 8.080 1.070 8.090 1.304 ;
        RECT 8.090 1.080 8.100 1.314 ;
        RECT 8.100 1.090 8.110 1.324 ;
        RECT 8.110 1.100 8.120 1.334 ;
        RECT 8.120 1.110 8.130 1.344 ;
        RECT 8.130 1.115 8.136 1.355 ;
        RECT 7.795 0.850 7.805 1.020 ;
        RECT 7.805 0.850 7.815 1.030 ;
        RECT 7.815 0.850 7.825 1.040 ;
        RECT 7.825 0.850 7.835 1.050 ;
        RECT 7.835 0.850 7.845 1.060 ;
        RECT 7.845 0.850 7.855 1.070 ;
        RECT 7.855 0.850 7.865 1.080 ;
        RECT 7.865 0.850 7.871 1.090 ;
  END 
END FFDQSRHDLXHT

MACRO FFDQSRHD2XHT
  CLASS  CORE ;
  FOREIGN FFDQSRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.890 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.030 0.720 11.200 1.375 ;
        RECT 11.030 1.205 11.380 1.375 ;
        RECT 11.170 0.720 11.200 2.960 ;
        RECT 11.030 1.945 11.200 2.960 ;
        RECT 11.170 1.205 11.380 2.115 ;
        RECT 11.030 1.945 11.380 2.115 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.675 1.520 2.070 2.365 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.380 1.260 3.860 1.685 ;
        RECT 3.380 1.315 3.910 1.685 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.675 -0.300 0.975 0.715 ;
        RECT 1.625 -0.300 1.925 0.805 ;
        RECT 3.465 -0.300 3.765 1.020 ;
        RECT 6.395 -0.300 6.565 1.120 ;
        RECT 8.300 -0.300 8.600 0.815 ;
        RECT 10.385 -0.300 10.685 1.055 ;
        RECT 11.485 -0.300 11.785 1.055 ;
        RECT 0.000 -0.300 11.890 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.240 1.585 0.725 2.015 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 9.940 1.555 10.250 2.210 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.735 0.925 3.990 ;
        RECT 1.625 2.925 1.925 3.990 ;
        RECT 3.675 3.025 4.655 3.990 ;
        RECT 6.315 2.995 6.615 3.990 ;
        RECT 8.500 2.330 8.670 3.990 ;
        RECT 10.050 2.975 10.690 3.990 ;
        RECT 11.485 2.295 11.785 3.990 ;
        RECT 0.000 3.390 11.890 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 1.075 1.295 ;
        RECT 0.905 1.125 1.075 2.365 ;
        RECT 0.105 2.195 1.075 2.365 ;
        RECT 2.365 0.550 3.175 0.720 ;
        RECT 3.005 0.550 3.175 2.115 ;
        RECT 2.875 1.945 3.175 2.115 ;
        RECT 4.020 0.990 4.325 1.160 ;
        RECT 4.155 0.990 4.325 2.080 ;
        RECT 4.015 1.910 4.325 2.080 ;
        RECT 4.155 1.610 4.935 1.780 ;
        RECT 2.455 0.925 2.625 2.495 ;
        RECT 2.455 0.925 2.780 1.225 ;
        RECT 5.115 1.610 5.285 2.495 ;
        RECT 2.455 2.325 5.285 2.495 ;
        RECT 5.115 1.610 5.590 1.780 ;
        RECT 4.530 0.990 4.830 1.295 ;
        RECT 4.530 1.125 5.865 1.295 ;
        RECT 5.695 1.060 5.865 1.360 ;
        RECT 4.160 0.480 4.460 0.670 ;
        RECT 4.160 0.500 5.260 0.670 ;
        RECT 5.080 0.500 5.260 0.880 ;
        RECT 5.480 2.045 5.710 2.215 ;
        RECT 5.080 0.710 6.215 0.880 ;
        RECT 6.045 0.710 6.215 1.710 ;
        RECT 5.990 1.540 6.825 1.710 ;
        RECT 5.820 1.540 5.830 2.170 ;
        RECT 5.830 1.540 5.840 2.160 ;
        RECT 5.840 1.540 5.850 2.150 ;
        RECT 5.850 1.540 5.860 2.140 ;
        RECT 5.860 1.540 5.870 2.130 ;
        RECT 5.870 1.540 5.880 2.120 ;
        RECT 5.880 1.540 5.890 2.110 ;
        RECT 5.890 1.540 5.900 2.100 ;
        RECT 5.900 1.540 5.910 2.090 ;
        RECT 5.910 1.540 5.920 2.080 ;
        RECT 5.920 1.540 5.930 2.070 ;
        RECT 5.930 1.540 5.940 2.060 ;
        RECT 5.940 1.540 5.950 2.050 ;
        RECT 5.950 1.540 5.960 2.040 ;
        RECT 5.960 1.540 5.970 2.030 ;
        RECT 5.970 1.540 5.980 2.020 ;
        RECT 5.980 1.540 5.990 2.010 ;
        RECT 5.785 1.970 5.795 2.204 ;
        RECT 5.795 1.960 5.805 2.194 ;
        RECT 5.805 1.950 5.815 2.184 ;
        RECT 5.815 1.940 5.821 2.180 ;
        RECT 5.710 2.045 5.720 2.215 ;
        RECT 5.720 2.035 5.730 2.215 ;
        RECT 5.730 2.025 5.740 2.215 ;
        RECT 5.740 2.015 5.750 2.215 ;
        RECT 5.750 2.005 5.760 2.215 ;
        RECT 5.760 1.995 5.770 2.215 ;
        RECT 5.770 1.985 5.780 2.215 ;
        RECT 5.780 1.975 5.786 2.215 ;
        RECT 1.255 1.060 1.425 2.715 ;
        RECT 2.105 2.545 2.275 2.845 ;
        RECT 1.255 2.545 2.275 2.715 ;
        RECT 2.365 2.675 2.665 3.085 ;
        RECT 5.465 2.395 5.635 2.845 ;
        RECT 2.105 2.675 5.635 2.845 ;
        RECT 5.465 2.395 5.865 2.565 ;
        RECT 6.040 2.295 6.965 2.465 ;
        RECT 7.340 2.595 7.855 2.765 ;
        RECT 7.265 2.530 7.275 2.764 ;
        RECT 7.275 2.540 7.285 2.764 ;
        RECT 7.285 2.550 7.295 2.764 ;
        RECT 7.295 2.560 7.305 2.764 ;
        RECT 7.305 2.570 7.315 2.764 ;
        RECT 7.315 2.580 7.325 2.764 ;
        RECT 7.325 2.590 7.335 2.764 ;
        RECT 7.335 2.595 7.341 2.765 ;
        RECT 7.040 2.305 7.050 2.539 ;
        RECT 7.050 2.315 7.060 2.549 ;
        RECT 7.060 2.325 7.070 2.559 ;
        RECT 7.070 2.335 7.080 2.569 ;
        RECT 7.080 2.345 7.090 2.579 ;
        RECT 7.090 2.355 7.100 2.589 ;
        RECT 7.100 2.365 7.110 2.599 ;
        RECT 7.110 2.375 7.120 2.609 ;
        RECT 7.120 2.385 7.130 2.619 ;
        RECT 7.130 2.395 7.140 2.629 ;
        RECT 7.140 2.405 7.150 2.639 ;
        RECT 7.150 2.415 7.160 2.649 ;
        RECT 7.160 2.425 7.170 2.659 ;
        RECT 7.170 2.435 7.180 2.669 ;
        RECT 7.180 2.445 7.190 2.679 ;
        RECT 7.190 2.455 7.200 2.689 ;
        RECT 7.200 2.465 7.210 2.699 ;
        RECT 7.210 2.475 7.220 2.709 ;
        RECT 7.220 2.485 7.230 2.719 ;
        RECT 7.230 2.495 7.240 2.729 ;
        RECT 7.240 2.505 7.250 2.739 ;
        RECT 7.250 2.515 7.260 2.749 ;
        RECT 7.260 2.520 7.266 2.760 ;
        RECT 6.965 2.295 6.975 2.465 ;
        RECT 6.975 2.295 6.985 2.475 ;
        RECT 6.985 2.295 6.995 2.485 ;
        RECT 6.995 2.295 7.005 2.495 ;
        RECT 7.005 2.295 7.015 2.505 ;
        RECT 7.015 2.295 7.025 2.515 ;
        RECT 7.025 2.295 7.035 2.525 ;
        RECT 7.035 2.295 7.041 2.535 ;
        RECT 5.965 2.295 5.975 2.529 ;
        RECT 5.975 2.295 5.985 2.519 ;
        RECT 5.985 2.295 5.995 2.509 ;
        RECT 5.995 2.295 6.005 2.499 ;
        RECT 6.005 2.295 6.015 2.489 ;
        RECT 6.015 2.295 6.025 2.479 ;
        RECT 6.025 2.295 6.035 2.469 ;
        RECT 6.035 2.295 6.041 2.465 ;
        RECT 5.940 2.320 5.950 2.554 ;
        RECT 5.950 2.310 5.960 2.544 ;
        RECT 5.960 2.300 5.966 2.540 ;
        RECT 5.865 2.395 5.875 2.565 ;
        RECT 5.875 2.385 5.885 2.565 ;
        RECT 5.885 2.375 5.895 2.565 ;
        RECT 5.895 2.365 5.905 2.565 ;
        RECT 5.905 2.355 5.915 2.565 ;
        RECT 5.915 2.345 5.925 2.565 ;
        RECT 5.925 2.335 5.935 2.565 ;
        RECT 5.935 2.325 5.941 2.565 ;
        RECT 5.625 3.040 5.960 3.210 ;
        RECT 6.215 2.645 6.705 2.815 ;
        RECT 7.560 1.155 7.690 1.325 ;
        RECT 7.115 2.980 8.100 3.150 ;
        RECT 8.100 2.205 8.110 3.149 ;
        RECT 8.110 2.215 8.120 3.149 ;
        RECT 8.120 2.225 8.130 3.149 ;
        RECT 8.130 2.235 8.140 3.149 ;
        RECT 8.140 2.245 8.150 3.149 ;
        RECT 8.150 2.255 8.160 3.149 ;
        RECT 8.160 2.265 8.170 3.149 ;
        RECT 8.170 2.275 8.180 3.149 ;
        RECT 8.180 2.285 8.190 3.149 ;
        RECT 8.190 2.295 8.200 3.149 ;
        RECT 8.200 2.305 8.210 3.149 ;
        RECT 8.210 2.315 8.220 3.149 ;
        RECT 8.220 2.325 8.230 3.149 ;
        RECT 8.230 2.335 8.240 3.149 ;
        RECT 8.240 2.345 8.250 3.149 ;
        RECT 8.250 2.355 8.260 3.149 ;
        RECT 8.260 2.365 8.270 3.149 ;
        RECT 7.860 1.965 7.870 2.239 ;
        RECT 7.870 1.975 7.880 2.249 ;
        RECT 7.880 1.985 7.890 2.259 ;
        RECT 7.890 1.995 7.900 2.269 ;
        RECT 7.900 2.005 7.910 2.279 ;
        RECT 7.910 2.015 7.920 2.289 ;
        RECT 7.920 2.025 7.930 2.299 ;
        RECT 7.930 2.035 7.940 2.309 ;
        RECT 7.940 2.045 7.950 2.319 ;
        RECT 7.950 2.055 7.960 2.329 ;
        RECT 7.960 2.065 7.970 2.339 ;
        RECT 7.970 2.075 7.980 2.349 ;
        RECT 7.980 2.085 7.990 2.359 ;
        RECT 7.990 2.095 8.000 2.369 ;
        RECT 8.000 2.105 8.010 2.379 ;
        RECT 8.010 2.115 8.020 2.389 ;
        RECT 8.020 2.125 8.030 2.399 ;
        RECT 8.030 2.135 8.040 2.409 ;
        RECT 8.040 2.145 8.050 2.419 ;
        RECT 8.050 2.155 8.060 2.429 ;
        RECT 8.060 2.165 8.070 2.439 ;
        RECT 8.070 2.175 8.080 2.449 ;
        RECT 8.080 2.185 8.090 2.459 ;
        RECT 8.090 2.195 8.100 2.469 ;
        RECT 7.690 1.155 7.700 2.069 ;
        RECT 7.700 1.155 7.710 2.079 ;
        RECT 7.710 1.155 7.720 2.089 ;
        RECT 7.720 1.155 7.730 2.099 ;
        RECT 7.730 1.155 7.740 2.109 ;
        RECT 7.740 1.155 7.750 2.119 ;
        RECT 7.750 1.155 7.760 2.129 ;
        RECT 7.760 1.155 7.770 2.139 ;
        RECT 7.770 1.155 7.780 2.149 ;
        RECT 7.780 1.155 7.790 2.159 ;
        RECT 7.790 1.155 7.800 2.169 ;
        RECT 7.800 1.155 7.810 2.179 ;
        RECT 7.810 1.155 7.820 2.189 ;
        RECT 7.820 1.155 7.830 2.199 ;
        RECT 7.830 1.155 7.840 2.209 ;
        RECT 7.840 1.155 7.850 2.219 ;
        RECT 7.850 1.155 7.860 2.229 ;
        RECT 7.040 2.915 7.050 3.149 ;
        RECT 7.050 2.925 7.060 3.149 ;
        RECT 7.060 2.935 7.070 3.149 ;
        RECT 7.070 2.945 7.080 3.149 ;
        RECT 7.080 2.955 7.090 3.149 ;
        RECT 7.090 2.965 7.100 3.149 ;
        RECT 7.100 2.975 7.110 3.149 ;
        RECT 7.110 2.980 7.116 3.150 ;
        RECT 6.780 2.655 6.790 2.889 ;
        RECT 6.790 2.665 6.800 2.899 ;
        RECT 6.800 2.675 6.810 2.909 ;
        RECT 6.810 2.685 6.820 2.919 ;
        RECT 6.820 2.695 6.830 2.929 ;
        RECT 6.830 2.705 6.840 2.939 ;
        RECT 6.840 2.715 6.850 2.949 ;
        RECT 6.850 2.725 6.860 2.959 ;
        RECT 6.860 2.735 6.870 2.969 ;
        RECT 6.870 2.745 6.880 2.979 ;
        RECT 6.880 2.755 6.890 2.989 ;
        RECT 6.890 2.765 6.900 2.999 ;
        RECT 6.900 2.775 6.910 3.009 ;
        RECT 6.910 2.785 6.920 3.019 ;
        RECT 6.920 2.795 6.930 3.029 ;
        RECT 6.930 2.805 6.940 3.039 ;
        RECT 6.940 2.815 6.950 3.049 ;
        RECT 6.950 2.825 6.960 3.059 ;
        RECT 6.960 2.835 6.970 3.069 ;
        RECT 6.970 2.845 6.980 3.079 ;
        RECT 6.980 2.855 6.990 3.089 ;
        RECT 6.990 2.865 7.000 3.099 ;
        RECT 7.000 2.875 7.010 3.109 ;
        RECT 7.010 2.885 7.020 3.119 ;
        RECT 7.020 2.895 7.030 3.129 ;
        RECT 7.030 2.905 7.040 3.139 ;
        RECT 6.705 2.645 6.715 2.815 ;
        RECT 6.715 2.645 6.725 2.825 ;
        RECT 6.725 2.645 6.735 2.835 ;
        RECT 6.735 2.645 6.745 2.845 ;
        RECT 6.745 2.645 6.755 2.855 ;
        RECT 6.755 2.645 6.765 2.865 ;
        RECT 6.765 2.645 6.775 2.875 ;
        RECT 6.775 2.645 6.781 2.885 ;
        RECT 6.140 2.645 6.150 2.879 ;
        RECT 6.150 2.645 6.160 2.869 ;
        RECT 6.160 2.645 6.170 2.859 ;
        RECT 6.170 2.645 6.180 2.849 ;
        RECT 6.180 2.645 6.190 2.839 ;
        RECT 6.190 2.645 6.200 2.829 ;
        RECT 6.200 2.645 6.210 2.819 ;
        RECT 6.210 2.645 6.216 2.815 ;
        RECT 6.130 2.655 6.140 2.889 ;
        RECT 5.960 2.825 5.970 3.209 ;
        RECT 5.970 2.815 5.980 3.209 ;
        RECT 5.980 2.805 5.990 3.209 ;
        RECT 5.990 2.795 6.000 3.209 ;
        RECT 6.000 2.785 6.010 3.209 ;
        RECT 6.010 2.775 6.020 3.209 ;
        RECT 6.020 2.765 6.030 3.209 ;
        RECT 6.030 2.755 6.040 3.209 ;
        RECT 6.040 2.745 6.050 3.209 ;
        RECT 6.050 2.735 6.060 3.209 ;
        RECT 6.060 2.725 6.070 3.209 ;
        RECT 6.070 2.715 6.080 3.209 ;
        RECT 6.080 2.705 6.090 3.209 ;
        RECT 6.090 2.695 6.100 3.209 ;
        RECT 6.100 2.685 6.110 3.209 ;
        RECT 6.110 2.675 6.120 3.209 ;
        RECT 6.120 2.665 6.130 3.209 ;
        RECT 8.535 1.190 8.560 1.710 ;
        RECT 8.610 1.540 9.550 1.710 ;
        RECT 9.380 1.060 9.550 2.295 ;
        RECT 9.380 2.125 9.760 2.295 ;
        RECT 8.560 1.500 8.570 1.710 ;
        RECT 8.570 1.510 8.580 1.710 ;
        RECT 8.580 1.520 8.590 1.710 ;
        RECT 8.590 1.530 8.600 1.710 ;
        RECT 8.600 1.540 8.610 1.710 ;
        RECT 8.390 1.190 8.400 1.564 ;
        RECT 8.400 1.190 8.410 1.574 ;
        RECT 8.410 1.190 8.420 1.584 ;
        RECT 8.420 1.190 8.430 1.594 ;
        RECT 8.430 1.190 8.440 1.604 ;
        RECT 8.440 1.190 8.450 1.614 ;
        RECT 8.450 1.190 8.460 1.624 ;
        RECT 8.460 1.190 8.470 1.634 ;
        RECT 8.470 1.190 8.480 1.644 ;
        RECT 8.480 1.190 8.490 1.654 ;
        RECT 8.490 1.190 8.500 1.664 ;
        RECT 8.500 1.190 8.510 1.674 ;
        RECT 8.510 1.190 8.520 1.684 ;
        RECT 8.520 1.190 8.530 1.694 ;
        RECT 8.530 1.190 8.536 1.704 ;
        RECT 8.860 0.710 9.030 1.360 ;
        RECT 8.860 0.710 10.070 0.880 ;
        RECT 9.900 0.710 10.070 1.360 ;
        RECT 7.155 1.635 7.470 1.805 ;
        RECT 7.155 0.785 7.325 1.805 ;
        RECT 7.300 1.635 7.470 2.280 ;
        RECT 7.155 0.785 7.920 0.955 ;
        RECT 8.450 1.890 9.160 2.070 ;
        RECT 8.980 1.890 9.160 2.645 ;
        RECT 9.280 2.475 9.580 2.945 ;
        RECT 10.605 1.595 10.775 2.645 ;
        RECT 8.980 2.475 10.775 2.645 ;
        RECT 10.605 1.595 10.985 1.765 ;
        RECT 8.375 1.825 8.385 2.069 ;
        RECT 8.385 1.835 8.395 2.069 ;
        RECT 8.395 1.845 8.405 2.069 ;
        RECT 8.405 1.855 8.415 2.069 ;
        RECT 8.415 1.865 8.425 2.069 ;
        RECT 8.425 1.875 8.435 2.069 ;
        RECT 8.435 1.885 8.445 2.069 ;
        RECT 8.445 1.890 8.451 2.070 ;
        RECT 8.210 1.660 8.220 1.904 ;
        RECT 8.220 1.670 8.230 1.914 ;
        RECT 8.230 1.680 8.240 1.924 ;
        RECT 8.240 1.690 8.250 1.934 ;
        RECT 8.250 1.700 8.260 1.944 ;
        RECT 8.260 1.710 8.270 1.954 ;
        RECT 8.270 1.720 8.280 1.964 ;
        RECT 8.280 1.730 8.290 1.974 ;
        RECT 8.290 1.740 8.300 1.984 ;
        RECT 8.300 1.750 8.310 1.994 ;
        RECT 8.310 1.760 8.320 2.004 ;
        RECT 8.320 1.770 8.330 2.014 ;
        RECT 8.330 1.780 8.340 2.024 ;
        RECT 8.340 1.790 8.350 2.034 ;
        RECT 8.350 1.800 8.360 2.044 ;
        RECT 8.360 1.810 8.370 2.054 ;
        RECT 8.370 1.815 8.376 2.065 ;
        RECT 8.040 0.840 8.050 1.734 ;
        RECT 8.050 0.850 8.060 1.744 ;
        RECT 8.060 0.860 8.070 1.754 ;
        RECT 8.070 0.870 8.080 1.764 ;
        RECT 8.080 0.880 8.090 1.774 ;
        RECT 8.090 0.890 8.100 1.784 ;
        RECT 8.100 0.900 8.110 1.794 ;
        RECT 8.110 0.910 8.120 1.804 ;
        RECT 8.120 0.920 8.130 1.814 ;
        RECT 8.130 0.930 8.140 1.824 ;
        RECT 8.140 0.940 8.150 1.834 ;
        RECT 8.150 0.950 8.160 1.844 ;
        RECT 8.160 0.960 8.170 1.854 ;
        RECT 8.170 0.970 8.180 1.864 ;
        RECT 8.180 0.980 8.190 1.874 ;
        RECT 8.190 0.990 8.200 1.884 ;
        RECT 8.200 1.000 8.210 1.894 ;
        RECT 7.995 0.795 8.005 1.029 ;
        RECT 8.005 0.805 8.015 1.039 ;
        RECT 8.015 0.815 8.025 1.049 ;
        RECT 8.025 0.825 8.035 1.059 ;
        RECT 8.035 0.830 8.041 1.070 ;
        RECT 7.920 0.785 7.930 0.955 ;
        RECT 7.930 0.785 7.940 0.965 ;
        RECT 7.940 0.785 7.950 0.975 ;
        RECT 7.950 0.785 7.960 0.985 ;
        RECT 7.960 0.785 7.970 0.995 ;
        RECT 7.970 0.785 7.980 1.005 ;
        RECT 7.980 0.785 7.990 1.015 ;
        RECT 7.990 0.785 7.996 1.025 ;
  END 
END FFDQSRHD2XHT

MACRO FFDQSRHD1XHT
  CLASS  CORE ;
  FOREIGN FFDQSRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.070 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.700 0.720 10.970 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.265 2.070 1.845 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.380 1.410 3.850 2.030 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.505 -0.300 0.675 0.810 ;
        RECT 1.720 -0.300 2.020 0.565 ;
        RECT 3.500 -0.300 3.670 1.225 ;
        RECT 6.230 -0.300 6.400 1.220 ;
        RECT 8.125 -0.300 8.425 0.815 ;
        RECT 10.140 -0.300 10.440 0.715 ;
        RECT 0.000 -0.300 11.070 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.185 1.670 0.725 2.015 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 9.780 1.480 10.150 1.935 ;
        RECT 9.940 1.480 10.150 2.020 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.575 2.755 0.875 3.990 ;
        RECT 1.615 2.520 1.915 3.990 ;
        RECT 3.505 3.025 4.145 3.990 ;
        RECT 6.165 2.995 6.465 3.990 ;
        RECT 8.130 2.345 8.770 3.990 ;
        RECT 10.115 2.975 10.415 3.990 ;
        RECT 0.000 3.390 11.070 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 1.030 1.295 ;
        RECT 0.860 0.710 1.030 1.514 ;
        RECT 0.870 1.485 1.076 1.524 ;
        RECT 0.880 1.485 1.076 1.534 ;
        RECT 0.890 1.485 1.076 1.544 ;
        RECT 0.900 1.485 1.076 1.554 ;
        RECT 0.105 2.195 1.030 2.365 ;
        RECT 0.860 1.450 1.040 1.514 ;
        RECT 0.860 1.460 1.050 1.514 ;
        RECT 0.860 1.470 1.060 1.514 ;
        RECT 0.905 1.480 1.070 2.364 ;
        RECT 1.070 1.485 1.076 2.365 ;
        RECT 0.860 0.710 1.590 0.880 ;
        RECT 1.525 0.745 2.370 0.890 ;
        RECT 1.535 0.745 2.370 0.900 ;
        RECT 1.545 0.745 2.370 0.910 ;
        RECT 1.550 0.710 1.590 0.915 ;
        RECT 0.860 0.720 1.600 0.880 ;
        RECT 0.860 0.730 1.610 0.880 ;
        RECT 1.550 0.745 2.370 0.914 ;
        RECT 0.860 0.740 1.620 0.880 ;
        RECT 2.200 0.575 2.370 0.915 ;
        RECT 1.620 0.745 2.370 0.915 ;
        RECT 2.200 0.575 3.130 0.745 ;
        RECT 2.880 1.840 3.050 2.140 ;
        RECT 2.960 0.575 3.130 2.010 ;
        RECT 2.880 1.840 3.130 2.010 ;
        RECT 4.020 0.925 4.200 1.225 ;
        RECT 4.030 0.925 4.200 1.730 ;
        RECT 4.050 1.430 4.220 2.145 ;
        RECT 4.030 1.430 4.825 1.730 ;
        RECT 2.445 1.410 2.615 2.495 ;
        RECT 2.550 0.925 2.720 1.590 ;
        RECT 2.445 1.410 2.720 1.590 ;
        RECT 4.400 1.910 4.570 2.495 ;
        RECT 2.445 2.325 4.570 2.495 ;
        RECT 5.005 1.680 5.175 2.080 ;
        RECT 4.400 1.910 5.175 2.080 ;
        RECT 5.240 1.550 5.410 1.850 ;
        RECT 5.005 1.680 5.410 1.850 ;
        RECT 4.465 0.990 5.700 1.160 ;
        RECT 5.530 0.990 5.700 1.325 ;
        RECT 4.095 0.490 4.395 0.695 ;
        RECT 5.580 2.035 5.761 2.110 ;
        RECT 5.355 2.045 5.655 2.215 ;
        RECT 5.355 2.045 5.665 2.204 ;
        RECT 5.355 2.045 5.675 2.194 ;
        RECT 5.355 2.045 5.685 2.184 ;
        RECT 5.355 2.045 5.695 2.174 ;
        RECT 5.355 2.045 5.705 2.164 ;
        RECT 5.355 2.045 5.715 2.154 ;
        RECT 5.355 2.045 5.725 2.144 ;
        RECT 5.355 2.045 5.735 2.134 ;
        RECT 5.355 2.045 5.745 2.124 ;
        RECT 5.355 2.045 5.755 2.114 ;
        RECT 5.590 1.600 5.761 2.110 ;
        RECT 4.095 0.525 6.050 0.695 ;
        RECT 5.880 0.525 6.050 1.770 ;
        RECT 5.590 1.600 6.675 1.770 ;
        RECT 1.210 1.060 1.425 1.360 ;
        RECT 1.255 1.060 1.425 2.340 ;
        RECT 1.255 2.170 2.265 2.340 ;
        RECT 2.095 2.170 2.265 2.845 ;
        RECT 2.355 2.675 2.655 2.935 ;
        RECT 4.750 2.395 4.920 2.845 ;
        RECT 2.095 2.675 4.920 2.845 ;
        RECT 4.750 2.395 5.735 2.565 ;
        RECT 5.910 2.295 6.700 2.465 ;
        RECT 6.905 2.425 7.600 2.595 ;
        RECT 7.430 2.425 7.600 2.725 ;
        RECT 6.830 2.360 6.840 2.594 ;
        RECT 6.840 2.370 6.850 2.594 ;
        RECT 6.850 2.380 6.860 2.594 ;
        RECT 6.860 2.390 6.870 2.594 ;
        RECT 6.870 2.400 6.880 2.594 ;
        RECT 6.880 2.410 6.890 2.594 ;
        RECT 6.890 2.420 6.900 2.594 ;
        RECT 6.900 2.425 6.906 2.595 ;
        RECT 6.775 2.305 6.785 2.539 ;
        RECT 6.785 2.315 6.795 2.549 ;
        RECT 6.795 2.325 6.805 2.559 ;
        RECT 6.805 2.335 6.815 2.569 ;
        RECT 6.815 2.345 6.825 2.579 ;
        RECT 6.825 2.350 6.831 2.590 ;
        RECT 6.700 2.295 6.710 2.465 ;
        RECT 6.710 2.295 6.720 2.475 ;
        RECT 6.720 2.295 6.730 2.485 ;
        RECT 6.730 2.295 6.740 2.495 ;
        RECT 6.740 2.295 6.750 2.505 ;
        RECT 6.750 2.295 6.760 2.515 ;
        RECT 6.760 2.295 6.770 2.525 ;
        RECT 6.770 2.295 6.776 2.535 ;
        RECT 5.835 2.295 5.845 2.529 ;
        RECT 5.845 2.295 5.855 2.519 ;
        RECT 5.855 2.295 5.865 2.509 ;
        RECT 5.865 2.295 5.875 2.499 ;
        RECT 5.875 2.295 5.885 2.489 ;
        RECT 5.885 2.295 5.895 2.479 ;
        RECT 5.895 2.295 5.905 2.469 ;
        RECT 5.905 2.295 5.911 2.465 ;
        RECT 5.810 2.320 5.820 2.554 ;
        RECT 5.820 2.310 5.830 2.544 ;
        RECT 5.830 2.300 5.836 2.540 ;
        RECT 5.735 2.395 5.745 2.565 ;
        RECT 5.745 2.385 5.755 2.565 ;
        RECT 5.755 2.375 5.765 2.565 ;
        RECT 5.765 2.365 5.775 2.565 ;
        RECT 5.775 2.355 5.785 2.565 ;
        RECT 5.785 2.345 5.795 2.565 ;
        RECT 5.795 2.335 5.805 2.565 ;
        RECT 5.805 2.325 5.811 2.565 ;
        RECT 5.100 2.745 5.270 3.210 ;
        RECT 4.325 3.040 5.270 3.210 ;
        RECT 5.100 2.745 5.910 2.915 ;
        RECT 6.085 2.645 6.545 2.815 ;
        RECT 7.005 2.805 7.175 3.075 ;
        RECT 6.780 2.805 7.175 2.975 ;
        RECT 7.435 1.220 7.565 1.390 ;
        RECT 7.005 2.905 7.780 3.075 ;
        RECT 7.780 1.910 7.790 3.074 ;
        RECT 7.790 1.920 7.800 3.074 ;
        RECT 7.800 1.930 7.810 3.074 ;
        RECT 7.810 1.940 7.820 3.074 ;
        RECT 7.820 1.950 7.830 3.074 ;
        RECT 7.830 1.960 7.840 3.074 ;
        RECT 7.840 1.970 7.850 3.074 ;
        RECT 7.850 1.980 7.860 3.074 ;
        RECT 7.860 1.990 7.870 3.074 ;
        RECT 7.870 2.000 7.880 3.074 ;
        RECT 7.880 2.010 7.890 3.074 ;
        RECT 7.890 2.020 7.900 3.074 ;
        RECT 7.900 2.030 7.910 3.074 ;
        RECT 7.910 2.040 7.920 3.074 ;
        RECT 7.920 2.050 7.930 3.074 ;
        RECT 7.930 2.060 7.940 3.074 ;
        RECT 7.940 2.070 7.950 3.074 ;
        RECT 7.735 1.865 7.745 2.115 ;
        RECT 7.745 1.875 7.755 2.125 ;
        RECT 7.755 1.885 7.765 2.135 ;
        RECT 7.765 1.895 7.775 2.145 ;
        RECT 7.775 1.900 7.781 2.154 ;
        RECT 7.565 1.220 7.575 1.944 ;
        RECT 7.575 1.220 7.585 1.954 ;
        RECT 7.585 1.220 7.595 1.964 ;
        RECT 7.595 1.220 7.605 1.974 ;
        RECT 7.605 1.220 7.615 1.984 ;
        RECT 7.615 1.220 7.625 1.994 ;
        RECT 7.625 1.220 7.635 2.004 ;
        RECT 7.635 1.220 7.645 2.014 ;
        RECT 7.645 1.220 7.655 2.024 ;
        RECT 7.655 1.220 7.665 2.034 ;
        RECT 7.665 1.220 7.675 2.044 ;
        RECT 7.675 1.220 7.685 2.054 ;
        RECT 7.685 1.220 7.695 2.064 ;
        RECT 7.695 1.220 7.705 2.074 ;
        RECT 7.705 1.220 7.715 2.084 ;
        RECT 7.715 1.220 7.725 2.094 ;
        RECT 7.725 1.220 7.735 2.104 ;
        RECT 6.705 2.740 6.715 2.974 ;
        RECT 6.715 2.750 6.725 2.974 ;
        RECT 6.725 2.760 6.735 2.974 ;
        RECT 6.735 2.770 6.745 2.974 ;
        RECT 6.745 2.780 6.755 2.974 ;
        RECT 6.755 2.790 6.765 2.974 ;
        RECT 6.765 2.800 6.775 2.974 ;
        RECT 6.775 2.805 6.781 2.975 ;
        RECT 6.620 2.655 6.630 2.889 ;
        RECT 6.630 2.665 6.640 2.899 ;
        RECT 6.640 2.675 6.650 2.909 ;
        RECT 6.650 2.685 6.660 2.919 ;
        RECT 6.660 2.695 6.670 2.929 ;
        RECT 6.670 2.705 6.680 2.939 ;
        RECT 6.680 2.715 6.690 2.949 ;
        RECT 6.690 2.725 6.700 2.959 ;
        RECT 6.700 2.730 6.706 2.970 ;
        RECT 6.545 2.645 6.555 2.815 ;
        RECT 6.555 2.645 6.565 2.825 ;
        RECT 6.565 2.645 6.575 2.835 ;
        RECT 6.575 2.645 6.585 2.845 ;
        RECT 6.585 2.645 6.595 2.855 ;
        RECT 6.595 2.645 6.605 2.865 ;
        RECT 6.605 2.645 6.615 2.875 ;
        RECT 6.615 2.645 6.621 2.885 ;
        RECT 6.010 2.645 6.020 2.879 ;
        RECT 6.020 2.645 6.030 2.869 ;
        RECT 6.030 2.645 6.040 2.859 ;
        RECT 6.040 2.645 6.050 2.849 ;
        RECT 6.050 2.645 6.060 2.839 ;
        RECT 6.060 2.645 6.070 2.829 ;
        RECT 6.070 2.645 6.080 2.819 ;
        RECT 6.080 2.645 6.086 2.815 ;
        RECT 5.985 2.670 5.995 2.904 ;
        RECT 5.995 2.660 6.005 2.894 ;
        RECT 6.005 2.650 6.011 2.890 ;
        RECT 5.910 2.745 5.920 2.915 ;
        RECT 5.920 2.735 5.930 2.915 ;
        RECT 5.930 2.725 5.940 2.915 ;
        RECT 5.940 2.715 5.950 2.915 ;
        RECT 5.950 2.705 5.960 2.915 ;
        RECT 5.960 2.695 5.970 2.915 ;
        RECT 5.970 2.685 5.980 2.915 ;
        RECT 5.980 2.675 5.986 2.915 ;
        RECT 8.420 1.460 8.590 1.760 ;
        RECT 8.420 1.460 9.520 1.630 ;
        RECT 9.080 1.110 9.380 1.630 ;
        RECT 9.350 1.460 9.520 2.305 ;
        RECT 9.350 2.135 9.800 2.305 ;
        RECT 8.690 0.760 8.860 1.280 ;
        RECT 8.560 1.110 8.860 1.280 ;
        RECT 8.690 0.760 9.770 0.930 ;
        RECT 9.600 0.760 9.770 1.280 ;
        RECT 9.600 1.110 9.900 1.280 ;
        RECT 7.010 0.850 7.180 2.245 ;
        RECT 7.010 2.075 7.385 2.245 ;
        RECT 7.010 0.850 7.825 1.020 ;
        RECT 8.400 1.995 9.135 2.165 ;
        RECT 8.965 1.995 9.135 2.655 ;
        RECT 9.320 2.485 9.620 2.900 ;
        RECT 10.350 1.550 10.520 2.655 ;
        RECT 8.965 2.485 10.520 2.655 ;
        RECT 8.315 1.920 8.325 2.164 ;
        RECT 8.325 1.930 8.335 2.164 ;
        RECT 8.335 1.940 8.345 2.164 ;
        RECT 8.345 1.950 8.355 2.164 ;
        RECT 8.355 1.960 8.365 2.164 ;
        RECT 8.365 1.970 8.375 2.164 ;
        RECT 8.375 1.980 8.385 2.164 ;
        RECT 8.385 1.990 8.395 2.164 ;
        RECT 8.395 1.995 8.401 2.165 ;
        RECT 8.150 1.755 8.160 1.999 ;
        RECT 8.160 1.765 8.170 2.009 ;
        RECT 8.170 1.775 8.180 2.019 ;
        RECT 8.180 1.785 8.190 2.029 ;
        RECT 8.190 1.795 8.200 2.039 ;
        RECT 8.200 1.805 8.210 2.049 ;
        RECT 8.210 1.815 8.220 2.059 ;
        RECT 8.220 1.825 8.230 2.069 ;
        RECT 8.230 1.835 8.240 2.079 ;
        RECT 8.240 1.845 8.250 2.089 ;
        RECT 8.250 1.855 8.260 2.099 ;
        RECT 8.260 1.865 8.270 2.109 ;
        RECT 8.270 1.875 8.280 2.119 ;
        RECT 8.280 1.885 8.290 2.129 ;
        RECT 8.290 1.895 8.300 2.139 ;
        RECT 8.300 1.905 8.310 2.149 ;
        RECT 8.310 1.910 8.316 2.160 ;
        RECT 7.980 0.940 7.990 1.830 ;
        RECT 7.990 0.950 8.000 1.840 ;
        RECT 8.000 0.960 8.010 1.850 ;
        RECT 8.010 0.970 8.020 1.860 ;
        RECT 8.020 0.980 8.030 1.870 ;
        RECT 8.030 0.990 8.040 1.880 ;
        RECT 8.040 1.000 8.050 1.890 ;
        RECT 8.050 1.010 8.060 1.900 ;
        RECT 8.060 1.020 8.070 1.910 ;
        RECT 8.070 1.030 8.080 1.920 ;
        RECT 8.080 1.040 8.090 1.930 ;
        RECT 8.090 1.050 8.100 1.940 ;
        RECT 8.100 1.060 8.110 1.950 ;
        RECT 8.110 1.070 8.120 1.960 ;
        RECT 8.120 1.080 8.130 1.970 ;
        RECT 8.130 1.090 8.140 1.980 ;
        RECT 8.140 1.100 8.150 1.990 ;
        RECT 7.900 0.860 7.910 1.094 ;
        RECT 7.910 0.870 7.920 1.104 ;
        RECT 7.920 0.880 7.930 1.114 ;
        RECT 7.930 0.890 7.940 1.124 ;
        RECT 7.940 0.900 7.950 1.134 ;
        RECT 7.950 0.910 7.960 1.144 ;
        RECT 7.960 0.920 7.970 1.154 ;
        RECT 7.970 0.930 7.980 1.164 ;
        RECT 7.825 0.850 7.835 1.020 ;
        RECT 7.835 0.850 7.845 1.030 ;
        RECT 7.845 0.850 7.855 1.040 ;
        RECT 7.855 0.850 7.865 1.050 ;
        RECT 7.865 0.850 7.875 1.060 ;
        RECT 7.875 0.850 7.885 1.070 ;
        RECT 7.885 0.850 7.895 1.080 ;
        RECT 7.895 0.850 7.901 1.090 ;
  END 
END FFDQSRHD1XHT

MACRO FFDQSHDMXHT
  CLASS  CORE ;
  FOREIGN FFDQSHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.610 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.105 1.060 8.510 1.360 ;
        RECT 8.340 1.060 8.510 2.460 ;
        RECT 8.270 1.980 8.510 2.460 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.560 1.265 1.950 1.915 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.615 -0.300 0.915 0.825 ;
        RECT 1.495 -0.300 1.795 0.735 ;
        RECT 3.395 -0.300 3.695 1.020 ;
        RECT 4.475 -0.300 4.775 0.595 ;
        RECT 6.455 -0.300 6.625 0.720 ;
        RECT 8.040 -0.300 8.340 0.775 ;
        RECT 0.000 -0.300 8.610 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.085 0.755 4.385 0.945 ;
        RECT 5.035 0.605 5.205 0.945 ;
        RECT 4.085 0.775 5.205 0.945 ;
        RECT 5.035 0.605 6.225 0.775 ;
        RECT 6.055 0.605 6.225 1.130 ;
        RECT 7.025 0.540 7.195 1.130 ;
        RECT 6.055 0.920 7.195 1.130 ;
        RECT 7.025 0.540 7.430 0.710 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.810 0.955 3.990 ;
        RECT 1.460 2.810 1.630 3.990 ;
        RECT 3.395 3.160 3.695 3.990 ;
        RECT 4.475 3.160 4.775 3.990 ;
        RECT 6.445 2.745 6.745 3.990 ;
        RECT 7.585 2.745 7.885 3.990 ;
        RECT 0.000 3.390 8.610 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.510 0.830 2.680 1.485 ;
        RECT 2.510 1.305 2.865 1.485 ;
        RECT 2.695 1.305 2.865 2.280 ;
        RECT 2.535 2.110 2.865 2.280 ;
        RECT 2.695 1.675 3.905 1.845 ;
        RECT 3.135 1.245 4.370 1.415 ;
        RECT 4.200 1.125 4.370 2.215 ;
        RECT 3.945 2.045 4.370 2.215 ;
        RECT 4.200 1.125 4.985 1.295 ;
        RECT 0.170 0.590 0.340 1.295 ;
        RECT 0.170 2.460 0.340 2.900 ;
        RECT 0.170 1.125 0.965 1.295 ;
        RECT 0.795 1.125 0.965 2.630 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.170 2.460 1.980 2.630 ;
        RECT 1.810 2.460 1.980 2.980 ;
        RECT 1.810 2.810 5.545 2.980 ;
        RECT 1.170 0.915 1.380 1.360 ;
        RECT 1.210 0.915 1.380 2.280 ;
        RECT 1.170 1.980 1.380 2.280 ;
        RECT 1.170 0.915 2.330 1.085 ;
        RECT 2.160 0.480 2.330 2.630 ;
        RECT 2.160 1.740 2.485 1.910 ;
        RECT 2.160 0.480 2.985 0.650 ;
        RECT 5.070 1.565 5.240 2.630 ;
        RECT 5.230 1.265 5.400 1.735 ;
        RECT 5.070 1.565 5.400 1.735 ;
        RECT 5.825 2.425 6.125 2.630 ;
        RECT 2.160 2.460 6.125 2.630 ;
        RECT 6.280 1.325 7.545 1.495 ;
        RECT 7.375 0.890 7.545 2.215 ;
        RECT 6.995 2.045 7.545 2.215 ;
        RECT 5.535 0.955 5.835 1.125 ;
        RECT 5.665 0.955 5.835 2.215 ;
        RECT 5.560 2.045 5.860 2.215 ;
        RECT 6.330 1.675 6.500 2.565 ;
        RECT 5.665 1.675 7.075 1.845 ;
        RECT 7.920 1.610 8.090 2.565 ;
        RECT 6.330 2.395 8.090 2.565 ;
        RECT 7.920 1.610 8.100 1.910 ;
  END 
END FFDQSHDMXHT

MACRO FFDQSHDLXHT
  CLASS  CORE ;
  FOREIGN FFDQSHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.610 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.005 1.125 8.510 1.295 ;
        RECT 8.270 1.125 8.510 2.445 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.600 1.265 1.985 1.865 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.615 -0.300 0.915 0.865 ;
        RECT 1.535 -0.300 1.835 0.735 ;
        RECT 3.435 -0.300 3.735 1.045 ;
        RECT 4.550 -0.300 4.850 0.595 ;
        RECT 6.570 -0.300 6.740 0.760 ;
        RECT 8.005 -0.300 8.305 0.775 ;
        RECT 0.000 -0.300 8.610 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.155 0.755 4.455 0.945 ;
        RECT 5.165 0.605 5.335 0.945 ;
        RECT 4.155 0.775 5.335 0.945 ;
        RECT 5.165 0.605 6.355 0.775 ;
        RECT 6.185 0.605 6.355 1.145 ;
        RECT 7.005 0.920 7.340 1.145 ;
        RECT 7.170 0.540 7.340 1.145 ;
        RECT 6.185 0.975 7.340 1.145 ;
        RECT 7.170 0.540 7.545 0.710 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.685 2.810 0.985 3.990 ;
        RECT 1.500 2.810 1.670 3.990 ;
        RECT 3.435 3.235 3.735 3.990 ;
        RECT 4.550 3.235 4.850 3.990 ;
        RECT 6.575 2.745 6.875 3.990 ;
        RECT 7.655 2.745 7.955 3.990 ;
        RECT 0.000 3.390 8.610 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.550 1.190 2.815 1.390 ;
        RECT 2.550 0.830 2.720 1.390 ;
        RECT 2.645 1.190 2.815 2.355 ;
        RECT 2.570 2.055 2.815 2.355 ;
        RECT 2.645 1.675 3.945 1.845 ;
        RECT 3.175 1.245 4.470 1.415 ;
        RECT 4.270 1.125 4.470 2.215 ;
        RECT 3.985 2.045 4.470 2.215 ;
        RECT 4.270 1.125 5.115 1.295 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.195 0.965 2.365 ;
        RECT 0.795 1.125 0.965 2.630 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 2.460 2.020 2.630 ;
        RECT 1.850 2.460 2.020 3.055 ;
        RECT 1.850 2.885 5.515 3.055 ;
        RECT 1.210 0.915 1.400 1.360 ;
        RECT 1.230 0.915 1.400 2.280 ;
        RECT 1.210 1.980 1.400 2.280 ;
        RECT 1.210 0.915 2.370 1.085 ;
        RECT 2.200 0.480 2.370 2.705 ;
        RECT 2.200 1.610 2.460 1.910 ;
        RECT 2.200 0.480 2.995 0.650 ;
        RECT 5.360 1.265 5.530 2.705 ;
        RECT 5.955 2.460 6.255 2.705 ;
        RECT 2.200 2.535 6.255 2.705 ;
        RECT 6.395 1.325 7.690 1.495 ;
        RECT 7.520 0.890 7.690 2.215 ;
        RECT 7.155 2.045 7.690 2.215 ;
        RECT 5.755 0.955 5.925 2.280 ;
        RECT 5.665 0.955 5.965 1.125 ;
        RECT 6.460 1.675 6.630 2.565 ;
        RECT 5.755 1.675 7.205 1.845 ;
        RECT 7.920 1.540 8.090 2.565 ;
        RECT 6.460 2.395 8.090 2.565 ;
  END 
END FFDQSHDLXHT

MACRO FFDQSHD2XHT
  CLASS  CORE ;
  FOREIGN FFDQSHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.840 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.980 0.720 9.150 2.960 ;
        RECT 8.980 1.660 9.330 2.010 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.690 1.265 1.950 2.015 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.745 ;
        RECT 1.495 -0.300 1.795 0.735 ;
        RECT 3.395 -0.300 3.695 0.875 ;
        RECT 4.860 -0.300 5.030 0.780 ;
        RECT 6.890 -0.300 7.190 0.795 ;
        RECT 8.395 -0.300 8.695 1.055 ;
        RECT 9.435 -0.300 9.735 1.055 ;
        RECT 0.000 -0.300 9.840 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.545 0.555 2.015 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.925 0.960 5.095 1.495 ;
        RECT 4.405 1.325 5.095 1.495 ;
        RECT 5.210 0.605 5.380 1.130 ;
        RECT 4.925 0.960 5.380 1.130 ;
        RECT 5.210 0.605 6.570 0.775 ;
        RECT 6.400 0.605 6.570 1.145 ;
        RECT 7.415 0.920 7.770 1.145 ;
        RECT 7.600 0.560 7.770 1.145 ;
        RECT 6.400 0.975 7.770 1.145 ;
        RECT 7.600 0.560 7.930 0.730 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.545 2.810 0.845 3.990 ;
        RECT 1.495 3.095 1.795 3.990 ;
        RECT 3.510 3.095 3.810 3.990 ;
        RECT 4.650 3.095 4.950 3.990 ;
        RECT 6.890 2.790 7.190 3.990 ;
        RECT 8.000 2.975 8.640 3.990 ;
        RECT 9.435 2.295 9.735 3.990 ;
        RECT 0.000 3.390 9.840 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.510 0.830 2.845 1.130 ;
        RECT 2.675 0.830 2.845 2.215 ;
        RECT 2.590 2.045 2.890 2.215 ;
        RECT 2.675 1.675 3.855 1.845 ;
        RECT 3.685 1.610 3.855 1.910 ;
        RECT 3.135 1.245 3.435 1.465 ;
        RECT 3.135 1.245 4.225 1.415 ;
        RECT 4.055 0.945 4.225 2.215 ;
        RECT 4.055 2.045 4.370 2.215 ;
        RECT 4.055 0.945 4.585 1.115 ;
        RECT 4.055 1.675 5.275 1.845 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.195 0.965 2.365 ;
        RECT 0.795 1.125 0.965 2.630 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 2.460 2.035 2.630 ;
        RECT 1.865 2.460 2.035 2.915 ;
        RECT 2.930 2.745 3.230 2.995 ;
        RECT 1.865 2.745 5.855 2.915 ;
        RECT 5.675 2.745 5.855 3.185 ;
        RECT 5.675 3.015 6.295 3.185 ;
        RECT 1.160 0.915 1.380 1.360 ;
        RECT 1.210 0.915 1.380 2.280 ;
        RECT 1.160 1.980 1.380 2.280 ;
        RECT 1.160 0.915 2.330 1.085 ;
        RECT 2.160 0.480 2.330 1.985 ;
        RECT 2.215 1.685 2.385 2.565 ;
        RECT 2.160 1.685 2.420 1.985 ;
        RECT 2.160 0.480 2.995 0.650 ;
        RECT 5.520 1.290 5.690 2.565 ;
        RECT 2.215 2.395 6.385 2.565 ;
        RECT 6.215 2.395 6.385 2.770 ;
        RECT 6.620 1.325 8.120 1.495 ;
        RECT 7.950 0.910 8.120 2.215 ;
        RECT 7.450 2.045 8.120 2.215 ;
        RECT 5.880 0.955 6.180 1.125 ;
        RECT 6.010 0.955 6.180 2.215 ;
        RECT 5.925 2.045 6.245 2.215 ;
        RECT 7.020 1.675 7.190 2.610 ;
        RECT 6.010 1.675 7.435 1.845 ;
        RECT 8.630 1.540 8.800 2.610 ;
        RECT 7.020 2.440 8.800 2.610 ;
  END 
END FFDQSHD2XHT

MACRO FFDQSHD1XHT
  CLASS  CORE ;
  FOREIGN FFDQSHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.020 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.680 0.720 8.920 1.360 ;
        RECT 8.710 0.720 8.920 2.960 ;
        RECT 8.680 1.980 8.920 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.670 1.495 2.060 2.050 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.745 ;
        RECT 1.585 -0.300 1.885 0.880 ;
        RECT 3.475 -0.300 3.775 1.020 ;
        RECT 4.680 -0.300 4.980 0.595 ;
        RECT 6.665 -0.300 6.965 0.575 ;
        RECT 8.095 -0.300 8.395 1.055 ;
        RECT 0.000 -0.300 9.020 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.215 0.705 4.515 0.945 ;
        RECT 5.295 0.605 5.465 0.945 ;
        RECT 4.215 0.775 5.465 0.945 ;
        RECT 5.295 0.605 6.485 0.775 ;
        RECT 6.315 0.605 6.485 1.130 ;
        RECT 7.300 0.540 7.470 1.130 ;
        RECT 6.315 0.920 7.470 1.130 ;
        RECT 7.300 0.540 7.705 0.710 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 2.810 0.835 3.990 ;
        RECT 1.550 2.810 1.720 3.990 ;
        RECT 3.505 3.160 3.805 3.990 ;
        RECT 4.680 3.160 4.980 3.990 ;
        RECT 6.685 2.770 6.985 3.990 ;
        RECT 7.325 2.945 7.625 3.990 ;
        RECT 8.095 2.975 8.395 3.990 ;
        RECT 0.000 3.390 9.020 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.600 0.915 2.935 1.130 ;
        RECT 2.600 0.830 2.770 1.130 ;
        RECT 2.720 1.980 2.890 2.280 ;
        RECT 2.765 0.915 2.935 2.215 ;
        RECT 2.720 1.980 2.935 2.215 ;
        RECT 2.765 1.675 4.005 1.845 ;
        RECT 3.225 1.245 4.355 1.415 ;
        RECT 4.185 1.125 4.355 2.215 ;
        RECT 4.055 2.045 4.355 2.215 ;
        RECT 4.185 1.125 5.245 1.295 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.195 0.965 2.365 ;
        RECT 0.795 1.125 0.965 2.630 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 2.460 2.070 2.630 ;
        RECT 1.900 2.460 2.070 2.980 ;
        RECT 1.900 2.810 5.755 2.980 ;
        RECT 1.150 1.060 1.380 1.360 ;
        RECT 1.210 1.060 1.380 2.280 ;
        RECT 1.150 1.980 1.380 2.280 ;
        RECT 1.150 1.060 2.420 1.230 ;
        RECT 2.250 0.480 2.420 2.630 ;
        RECT 2.250 1.685 2.510 1.985 ;
        RECT 2.250 0.480 3.075 0.650 ;
        RECT 5.445 1.645 5.615 2.630 ;
        RECT 5.490 1.245 5.660 1.815 ;
        RECT 5.445 1.645 5.660 1.815 ;
        RECT 2.250 2.460 6.300 2.630 ;
        RECT 6.130 2.460 6.300 2.795 ;
        RECT 6.535 1.325 7.820 1.495 ;
        RECT 7.650 0.890 7.820 2.215 ;
        RECT 7.235 2.045 7.820 2.215 ;
        RECT 5.795 0.955 6.095 1.125 ;
        RECT 5.925 0.955 6.095 2.215 ;
        RECT 5.795 2.045 6.095 2.215 ;
        RECT 6.590 1.675 6.760 2.590 ;
        RECT 5.925 1.675 7.335 1.845 ;
        RECT 8.330 1.530 8.500 2.590 ;
        RECT 6.590 2.420 8.500 2.590 ;
        RECT 8.330 1.530 8.510 1.830 ;
  END 
END FFDQSHD1XHT

MACRO FFDQRHDMXHT
  CLASS  CORE ;
  FOREIGN FFDQRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.840 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.500 1.040 9.740 1.340 ;
        RECT 9.570 1.040 9.740 2.450 ;
        RECT 9.500 1.980 9.740 2.450 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.695 1.270 1.985 1.945 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.430 1.505 5.885 2.010 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.825 ;
        RECT 1.535 -0.300 1.835 0.740 ;
        RECT 3.465 -0.300 3.765 1.020 ;
        RECT 4.455 -0.300 4.755 0.595 ;
        RECT 5.525 -0.300 5.695 0.810 ;
        RECT 7.465 -0.300 7.765 0.575 ;
        RECT 8.915 -0.300 9.215 1.125 ;
        RECT 0.000 -0.300 9.840 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.010 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 2.810 0.865 3.990 ;
        RECT 1.495 2.810 1.665 3.990 ;
        RECT 3.435 3.195 3.735 3.990 ;
        RECT 5.535 3.195 5.835 3.990 ;
        RECT 7.565 2.745 7.865 3.990 ;
        RECT 8.885 2.825 9.185 3.990 ;
        RECT 0.000 3.390 9.840 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.550 1.190 2.875 1.390 ;
        RECT 2.550 0.830 2.720 1.390 ;
        RECT 2.705 1.190 2.875 2.315 ;
        RECT 2.545 2.080 2.875 2.315 ;
        RECT 2.705 1.675 3.935 1.845 ;
        RECT 3.205 1.245 4.285 1.415 ;
        RECT 4.080 0.775 4.250 1.415 ;
        RECT 4.115 1.245 4.285 2.215 ;
        RECT 4.115 2.045 4.655 2.215 ;
        RECT 4.940 0.480 5.110 0.945 ;
        RECT 4.080 0.775 5.110 0.945 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.190 0.965 2.360 ;
        RECT 0.795 1.125 0.965 2.630 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 2.460 2.015 2.630 ;
        RECT 1.845 2.460 2.015 3.015 ;
        RECT 5.860 2.745 6.030 3.015 ;
        RECT 1.845 2.845 6.030 3.015 ;
        RECT 5.860 2.745 6.605 2.915 ;
        RECT 1.210 0.920 1.400 1.360 ;
        RECT 1.230 0.920 1.400 2.280 ;
        RECT 1.210 1.980 1.400 2.280 ;
        RECT 1.210 0.920 2.365 1.090 ;
        RECT 2.195 0.480 2.365 2.665 ;
        RECT 2.195 1.720 2.525 1.890 ;
        RECT 2.195 0.480 3.025 0.650 ;
        RECT 5.505 2.395 5.675 2.665 ;
        RECT 2.195 2.495 5.675 2.665 ;
        RECT 6.245 1.330 6.415 2.565 ;
        RECT 6.225 1.330 6.525 1.500 ;
        RECT 5.505 2.395 7.185 2.565 ;
        RECT 6.885 2.395 7.185 2.595 ;
        RECT 4.465 1.595 5.210 1.765 ;
        RECT 5.040 1.125 5.210 2.280 ;
        RECT 5.875 0.605 6.045 1.295 ;
        RECT 5.015 1.125 6.045 1.295 ;
        RECT 7.090 0.605 7.260 0.945 ;
        RECT 5.875 0.605 7.260 0.775 ;
        RECT 7.090 0.775 8.735 0.945 ;
        RECT 8.565 0.775 8.735 1.730 ;
        RECT 8.015 1.125 8.385 1.495 ;
        RECT 7.255 1.325 8.385 1.495 ;
        RECT 8.215 1.125 8.385 2.215 ;
        RECT 8.215 2.045 8.785 2.215 ;
        RECT 6.515 0.955 6.875 1.125 ;
        RECT 6.705 0.955 6.875 2.215 ;
        RECT 6.620 2.045 6.920 2.215 ;
        RECT 6.705 1.675 8.035 1.845 ;
        RECT 7.865 1.675 8.035 2.565 ;
        RECT 9.150 1.545 9.320 2.565 ;
        RECT 7.865 2.395 9.320 2.565 ;
  END 
END FFDQRHDMXHT

MACRO FFDQRHDLXHT
  CLASS  CORE ;
  FOREIGN FFDQRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.840 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.500 1.060 9.740 1.360 ;
        RECT 9.530 1.060 9.740 2.280 ;
        RECT 9.500 1.980 9.740 2.280 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.600 1.270 1.990 1.800 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.430 1.515 5.885 2.010 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.855 ;
        RECT 1.535 -0.300 1.835 0.740 ;
        RECT 3.465 -0.300 3.765 1.020 ;
        RECT 4.455 -0.300 4.755 0.595 ;
        RECT 5.525 -0.300 5.695 0.810 ;
        RECT 7.465 -0.300 7.765 0.575 ;
        RECT 8.950 -0.300 9.120 1.190 ;
        RECT 0.000 -0.300 9.840 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.010 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 2.810 0.865 3.990 ;
        RECT 1.495 2.810 1.665 3.990 ;
        RECT 3.435 3.195 3.735 3.990 ;
        RECT 5.535 3.195 5.835 3.990 ;
        RECT 7.565 2.745 7.865 3.990 ;
        RECT 8.885 2.800 9.185 3.990 ;
        RECT 0.000 3.390 9.840 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.550 1.190 2.875 1.390 ;
        RECT 2.550 0.830 2.720 1.390 ;
        RECT 2.705 1.190 2.875 2.260 ;
        RECT 2.545 2.090 2.875 2.260 ;
        RECT 2.705 1.675 3.935 1.845 ;
        RECT 3.205 1.245 4.285 1.415 ;
        RECT 4.110 0.775 4.280 1.415 ;
        RECT 4.115 1.245 4.285 2.215 ;
        RECT 4.115 2.045 4.655 2.215 ;
        RECT 4.940 0.480 5.110 0.945 ;
        RECT 4.110 0.775 5.110 0.945 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.190 0.965 2.360 ;
        RECT 0.795 1.125 0.965 2.630 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 2.460 2.015 2.630 ;
        RECT 1.845 2.460 2.015 3.015 ;
        RECT 5.860 2.745 6.030 3.015 ;
        RECT 1.845 2.845 6.030 3.015 ;
        RECT 5.860 2.745 6.480 2.915 ;
        RECT 1.210 0.920 1.400 1.360 ;
        RECT 1.230 0.920 1.400 2.280 ;
        RECT 1.210 1.980 1.400 2.280 ;
        RECT 1.210 0.920 2.365 1.090 ;
        RECT 2.195 0.480 2.365 2.665 ;
        RECT 2.195 1.720 2.525 1.890 ;
        RECT 2.195 0.480 3.025 0.650 ;
        RECT 5.505 2.395 5.675 2.665 ;
        RECT 2.195 2.495 5.675 2.665 ;
        RECT 6.245 1.330 6.415 2.565 ;
        RECT 6.225 1.330 6.525 1.500 ;
        RECT 5.505 2.395 7.185 2.565 ;
        RECT 6.885 2.395 7.185 2.585 ;
        RECT 4.465 1.585 5.210 1.755 ;
        RECT 5.040 1.125 5.210 2.280 ;
        RECT 5.875 0.605 6.045 1.295 ;
        RECT 5.015 1.125 6.045 1.295 ;
        RECT 7.090 0.605 7.260 0.945 ;
        RECT 5.875 0.605 7.260 0.775 ;
        RECT 7.090 0.775 8.735 0.945 ;
        RECT 8.565 0.775 8.735 1.765 ;
        RECT 7.255 1.325 8.385 1.495 ;
        RECT 8.015 1.125 8.315 1.495 ;
        RECT 8.215 1.325 8.385 2.215 ;
        RECT 8.215 2.045 8.785 2.215 ;
        RECT 6.515 0.955 6.875 1.125 ;
        RECT 6.705 0.955 6.875 2.215 ;
        RECT 6.620 2.045 6.920 2.215 ;
        RECT 6.705 1.675 8.035 1.845 ;
        RECT 7.865 1.675 8.035 2.565 ;
        RECT 9.150 1.525 9.320 2.565 ;
        RECT 7.865 2.395 9.320 2.565 ;
  END 
END FFDQRHDLXHT

MACRO FFDQRHD2XHT
  CLASS  CORE ;
  FOREIGN FFDQRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.800 0.720 9.970 2.960 ;
        RECT 9.800 1.630 10.150 2.015 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.270 2.140 1.840 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.655 1.555 6.050 1.855 ;
        RECT 5.695 1.555 6.050 2.170 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.745 ;
        RECT 1.690 -0.300 1.990 1.020 ;
        RECT 3.610 -0.300 3.910 1.020 ;
        RECT 4.680 -0.300 4.980 0.595 ;
        RECT 5.850 -0.300 6.020 0.780 ;
        RECT 7.685 -0.300 7.985 0.595 ;
        RECT 9.215 -0.300 9.515 1.055 ;
        RECT 10.255 -0.300 10.555 1.055 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.600 2.810 0.900 3.990 ;
        RECT 1.690 3.140 1.990 3.990 ;
        RECT 3.545 3.140 3.845 3.990 ;
        RECT 5.755 3.095 6.055 3.990 ;
        RECT 7.785 2.810 8.085 3.990 ;
        RECT 9.215 2.975 9.515 3.990 ;
        RECT 10.255 2.295 10.555 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.705 1.190 3.030 1.370 ;
        RECT 2.705 0.885 2.875 1.370 ;
        RECT 2.860 1.190 3.030 2.260 ;
        RECT 2.705 2.090 3.030 2.260 ;
        RECT 2.860 1.675 4.090 1.845 ;
        RECT 3.360 1.245 4.440 1.415 ;
        RECT 4.195 0.735 4.365 1.415 ;
        RECT 4.270 1.245 4.440 2.215 ;
        RECT 4.270 2.045 4.810 2.215 ;
        RECT 5.160 0.480 5.330 0.945 ;
        RECT 4.195 0.775 5.330 0.945 ;
        RECT 0.105 1.125 1.020 1.295 ;
        RECT 0.105 2.220 1.020 2.390 ;
        RECT 0.850 1.125 1.020 2.630 ;
        RECT 0.850 1.525 1.085 1.825 ;
        RECT 0.850 2.460 2.175 2.630 ;
        RECT 2.005 2.460 2.175 2.960 ;
        RECT 3.010 2.790 3.310 2.975 ;
        RECT 5.325 2.745 5.495 2.960 ;
        RECT 2.005 2.790 5.495 2.960 ;
        RECT 5.325 2.745 6.655 2.915 ;
        RECT 6.485 2.745 6.655 3.210 ;
        RECT 6.485 3.040 7.315 3.210 ;
        RECT 1.245 1.060 1.435 1.360 ;
        RECT 1.265 1.060 1.435 2.280 ;
        RECT 1.245 1.980 1.435 2.280 ;
        RECT 1.245 2.090 2.525 2.280 ;
        RECT 2.355 0.480 2.525 2.610 ;
        RECT 2.355 1.720 2.680 1.890 ;
        RECT 2.355 0.480 3.180 0.650 ;
        RECT 4.970 2.395 5.140 2.610 ;
        RECT 2.355 2.440 5.140 2.610 ;
        RECT 6.445 1.355 6.615 2.565 ;
        RECT 6.445 1.355 6.745 1.525 ;
        RECT 4.970 2.395 7.340 2.565 ;
        RECT 7.170 2.395 7.340 2.795 ;
        RECT 4.620 1.575 5.405 1.745 ;
        RECT 5.235 1.125 5.405 2.215 ;
        RECT 5.195 2.045 5.495 2.215 ;
        RECT 5.735 0.960 5.905 1.295 ;
        RECT 5.235 1.125 5.905 1.295 ;
        RECT 5.735 0.960 6.370 1.130 ;
        RECT 6.200 0.635 6.370 1.130 ;
        RECT 7.320 0.635 7.490 0.945 ;
        RECT 6.200 0.635 7.490 0.805 ;
        RECT 7.320 0.775 8.985 0.945 ;
        RECT 8.815 0.775 8.985 1.775 ;
        RECT 8.265 1.125 8.605 1.495 ;
        RECT 7.425 1.325 8.605 1.495 ;
        RECT 8.435 1.125 8.605 2.215 ;
        RECT 8.435 2.045 9.005 2.215 ;
        RECT 6.735 0.985 7.140 1.155 ;
        RECT 6.970 0.985 7.140 2.215 ;
        RECT 6.840 2.045 7.140 2.215 ;
        RECT 6.970 1.675 8.255 1.845 ;
        RECT 8.085 1.675 8.255 2.565 ;
        RECT 9.450 1.525 9.620 2.565 ;
        RECT 8.085 2.395 9.620 2.565 ;
  END 
END FFDQRHD2XHT

MACRO FFDQHDMXHT
  CLASS  CORE ;
  FOREIGN FFDQHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.200 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.860 1.060 8.100 1.360 ;
        RECT 7.890 1.060 8.100 2.460 ;
        RECT 7.860 1.980 8.100 2.460 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.600 1.265 1.985 1.760 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.825 ;
        RECT 1.535 -0.300 1.835 0.720 ;
        RECT 3.335 -0.300 3.635 0.605 ;
        RECT 4.395 -0.300 4.695 1.110 ;
        RECT 6.295 -0.300 6.595 0.470 ;
        RECT 7.340 -0.300 7.510 1.210 ;
        RECT 0.000 -0.300 8.200 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 2.745 0.865 3.990 ;
        RECT 1.500 2.760 1.670 3.990 ;
        RECT 3.435 3.160 3.735 3.990 ;
        RECT 4.405 3.160 4.705 3.990 ;
        RECT 6.305 2.745 6.605 3.990 ;
        RECT 7.245 2.745 7.545 3.990 ;
        RECT 0.000 3.390 8.200 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.550 0.865 2.720 2.280 ;
        RECT 2.550 1.675 3.955 1.845 ;
        RECT 3.950 0.840 4.120 1.445 ;
        RECT 3.175 1.275 4.305 1.445 ;
        RECT 4.135 1.275 4.305 2.215 ;
        RECT 3.895 2.045 4.305 2.215 ;
        RECT 4.135 1.410 4.815 1.580 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.195 0.965 2.365 ;
        RECT 0.795 1.125 0.965 2.565 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 2.395 2.020 2.565 ;
        RECT 1.850 2.395 2.020 3.010 ;
        RECT 2.855 2.810 3.155 3.010 ;
        RECT 1.850 2.840 3.155 3.010 ;
        RECT 2.855 2.810 5.395 2.980 ;
        RECT 1.210 0.995 1.400 1.295 ;
        RECT 1.230 0.995 1.400 2.215 ;
        RECT 1.145 2.045 2.370 2.215 ;
        RECT 2.200 0.515 2.370 2.660 ;
        RECT 2.200 2.460 2.575 2.660 ;
        RECT 2.200 0.515 2.995 0.685 ;
        RECT 4.995 0.500 5.165 2.630 ;
        RECT 4.995 0.500 5.395 0.670 ;
        RECT 4.995 2.440 5.905 2.630 ;
        RECT 2.200 2.460 5.905 2.630 ;
        RECT 6.055 1.220 7.160 1.390 ;
        RECT 6.830 0.785 7.000 1.390 ;
        RECT 6.990 1.220 7.160 2.215 ;
        RECT 6.735 2.045 7.160 2.215 ;
        RECT 5.410 0.875 5.580 2.215 ;
        RECT 5.345 2.045 5.645 2.215 ;
        RECT 6.385 1.675 6.555 2.565 ;
        RECT 5.410 1.675 6.810 1.845 ;
        RECT 7.510 1.520 7.680 2.565 ;
        RECT 6.385 2.395 7.680 2.565 ;
        RECT 7.510 1.520 7.700 1.820 ;
  END 
END FFDQHDMXHT

MACRO LATHDLXHT
  CLASS  CORE ;
  FOREIGN LATHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.150 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.805 1.060 5.975 2.425 ;
        RECT 5.805 2.085 6.050 2.425 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.545 0.510 4.935 0.720 ;
        RECT 4.765 0.510 4.935 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.670 1.585 2.245 1.950 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.495 0.510 2.930 ;
    END
  END G
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.785 ;
        RECT 1.655 -0.300 1.955 1.035 ;
        RECT 3.555 -0.300 3.855 1.295 ;
        RECT 5.220 -0.300 5.520 1.295 ;
        RECT 0.000 -0.300 6.150 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.120 0.860 3.990 ;
        RECT 1.715 2.530 2.015 3.990 ;
        RECT 3.495 2.925 3.795 3.990 ;
        RECT 5.190 2.925 5.490 3.990 ;
        RECT 0.000 3.390 6.150 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.020 0.340 2.280 ;
        RECT 0.170 1.520 1.030 1.820 ;
        RECT 1.210 1.020 1.380 2.300 ;
        RECT 1.210 2.130 2.465 2.300 ;
        RECT 2.265 0.705 2.435 1.385 ;
        RECT 1.210 1.215 2.435 1.385 ;
        RECT 2.295 2.130 2.465 3.095 ;
        RECT 2.265 0.705 2.695 0.875 ;
        RECT 2.295 2.925 3.115 3.095 ;
        RECT 3.345 1.850 3.645 2.020 ;
        RECT 3.475 1.850 3.645 2.395 ;
        RECT 4.105 1.125 4.475 1.295 ;
        RECT 4.305 1.125 4.475 2.395 ;
        RECT 3.475 2.225 4.475 2.395 ;
        RECT 4.305 1.520 4.585 1.820 ;
        RECT 2.670 1.060 2.870 1.360 ;
        RECT 2.700 1.060 2.870 2.745 ;
        RECT 2.700 1.500 4.125 1.670 ;
        RECT 5.455 1.520 5.625 2.745 ;
        RECT 2.700 2.575 5.625 2.745 ;
  END 
END LATHDLXHT

MACRO FFDQHDLXHT
  CLASS  CORE ;
  FOREIGN FFDQHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.200 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.860 1.060 8.100 1.360 ;
        RECT 7.890 1.060 8.100 2.280 ;
        RECT 7.860 1.980 8.100 2.280 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.600 1.265 1.985 1.670 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.855 ;
        RECT 1.535 -0.300 1.835 0.785 ;
        RECT 3.335 -0.300 3.635 0.565 ;
        RECT 4.405 -0.300 4.705 0.680 ;
        RECT 6.295 -0.300 6.595 0.550 ;
        RECT 7.340 -0.300 7.510 1.330 ;
        RECT 0.000 -0.300 8.200 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 2.745 0.865 3.990 ;
        RECT 1.500 2.745 1.670 3.990 ;
        RECT 3.435 3.160 3.735 3.990 ;
        RECT 4.405 3.160 4.705 3.990 ;
        RECT 6.305 2.745 6.605 3.990 ;
        RECT 7.245 2.745 7.545 3.990 ;
        RECT 0.000 3.390 8.200 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.550 0.865 2.720 2.280 ;
        RECT 2.550 1.675 3.955 1.845 ;
        RECT 3.960 0.840 4.130 1.445 ;
        RECT 3.175 1.275 4.815 1.445 ;
        RECT 4.645 1.275 4.815 2.215 ;
        RECT 3.895 2.045 4.815 2.215 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.195 0.965 2.365 ;
        RECT 0.795 1.125 0.965 2.565 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 2.395 2.020 2.565 ;
        RECT 1.850 2.395 2.020 2.995 ;
        RECT 2.855 2.810 3.025 2.995 ;
        RECT 1.850 2.825 3.025 2.995 ;
        RECT 2.855 2.810 5.285 2.980 ;
        RECT 1.210 1.060 1.400 1.360 ;
        RECT 1.230 1.060 1.400 2.215 ;
        RECT 1.145 2.045 2.370 2.215 ;
        RECT 2.200 0.515 2.370 2.645 ;
        RECT 2.200 2.460 2.575 2.645 ;
        RECT 2.200 0.515 2.995 0.685 ;
        RECT 4.995 0.525 5.165 2.630 ;
        RECT 4.995 0.525 5.385 0.695 ;
        RECT 2.200 2.460 5.865 2.630 ;
        RECT 6.055 1.220 7.160 1.390 ;
        RECT 6.830 0.785 7.000 1.390 ;
        RECT 6.990 1.220 7.160 2.215 ;
        RECT 6.735 2.045 7.160 2.215 ;
        RECT 5.410 0.875 5.580 2.215 ;
        RECT 5.345 2.045 5.645 2.215 ;
        RECT 6.385 1.675 6.555 2.565 ;
        RECT 5.410 1.675 6.810 1.845 ;
        RECT 7.510 1.520 7.680 2.565 ;
        RECT 6.385 2.395 7.680 2.565 ;
        RECT 7.510 1.520 7.700 1.820 ;
  END 
END FFDQHDLXHT

MACRO FFDQHD2XHT
  CLASS  CORE ;
  FOREIGN FFDQHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.020 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.160 0.720 8.330 2.960 ;
        RECT 8.160 1.640 8.510 2.015 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.585 1.265 2.080 1.670 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.745 ;
        RECT 1.630 -0.300 1.930 0.875 ;
        RECT 3.650 -0.300 3.950 1.020 ;
        RECT 4.700 -0.300 5.000 1.055 ;
        RECT 6.475 -0.300 6.645 0.780 ;
        RECT 7.640 -0.300 7.810 0.780 ;
        RECT 8.615 -0.300 8.915 1.055 ;
        RECT 0.000 -0.300 9.020 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.520 2.015 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.515 2.745 0.815 3.990 ;
        RECT 1.620 2.745 1.790 3.990 ;
        RECT 3.620 3.095 3.920 3.990 ;
        RECT 4.575 3.095 4.875 3.990 ;
        RECT 6.595 2.805 6.765 3.990 ;
        RECT 7.575 2.975 7.875 3.990 ;
        RECT 8.615 2.295 8.915 3.990 ;
        RECT 0.000 3.390 9.020 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.670 0.850 2.970 1.020 ;
        RECT 2.800 0.850 2.970 2.215 ;
        RECT 2.670 2.045 2.970 2.215 ;
        RECT 2.800 1.675 4.190 1.845 ;
        RECT 4.255 0.985 4.425 1.445 ;
        RECT 3.390 1.275 5.120 1.445 ;
        RECT 4.950 1.275 5.120 2.215 ;
        RECT 4.170 2.045 5.120 2.215 ;
        RECT 0.105 1.125 0.880 1.295 ;
        RECT 0.105 2.195 0.880 2.365 ;
        RECT 0.710 1.125 0.880 2.565 ;
        RECT 0.710 1.525 1.035 1.825 ;
        RECT 0.710 2.395 2.140 2.565 ;
        RECT 1.970 2.395 2.140 2.915 ;
        RECT 5.015 2.745 5.185 2.975 ;
        RECT 1.970 2.745 5.185 2.915 ;
        RECT 5.015 2.805 5.685 2.975 ;
        RECT 5.515 2.805 5.685 3.210 ;
        RECT 5.515 3.040 6.200 3.210 ;
        RECT 6.390 1.590 7.345 1.760 ;
        RECT 7.175 1.060 7.345 2.280 ;
        RECT 1.215 1.060 1.385 2.215 ;
        RECT 1.085 2.045 2.490 2.215 ;
        RECT 2.320 0.480 2.490 2.565 ;
        RECT 2.320 1.605 2.555 1.905 ;
        RECT 2.320 0.480 3.240 0.650 ;
        RECT 5.300 0.710 5.470 2.565 ;
        RECT 5.365 2.395 5.535 2.610 ;
        RECT 2.320 2.395 5.535 2.565 ;
        RECT 5.365 2.440 6.135 2.610 ;
        RECT 5.300 0.710 6.240 0.880 ;
        RECT 5.965 2.440 6.135 2.795 ;
        RECT 6.070 0.710 6.240 1.140 ;
        RECT 6.825 0.480 6.995 1.140 ;
        RECT 6.070 0.970 6.995 1.140 ;
        RECT 6.825 0.480 7.460 0.650 ;
        RECT 5.715 1.060 5.885 2.215 ;
        RECT 5.650 2.045 6.995 2.215 ;
        RECT 6.825 2.045 6.995 2.630 ;
        RECT 6.965 2.460 7.135 2.770 ;
        RECT 7.810 1.530 7.980 2.630 ;
        RECT 6.825 2.460 7.980 2.630 ;
  END 
END FFDQHD2XHT

MACRO FFDQHD1XHT
  CLASS  CORE ;
  FOREIGN FFDQHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.200 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.860 0.720 8.100 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.600 1.265 1.985 1.670 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.745 ;
        RECT 1.535 -0.300 1.835 0.720 ;
        RECT 3.345 -0.300 3.645 0.525 ;
        RECT 4.405 -0.300 4.705 1.040 ;
        RECT 6.295 -0.300 6.595 0.490 ;
        RECT 7.275 -0.300 7.575 1.055 ;
        RECT 0.000 -0.300 8.200 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 2.745 0.865 3.990 ;
        RECT 1.500 2.770 1.670 3.990 ;
        RECT 3.435 3.160 3.735 3.990 ;
        RECT 4.405 3.160 4.705 3.990 ;
        RECT 6.305 2.745 6.605 3.990 ;
        RECT 7.275 2.975 7.575 3.990 ;
        RECT 0.000 3.390 8.200 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.550 0.865 2.720 2.280 ;
        RECT 2.550 1.675 3.955 1.845 ;
        RECT 3.960 0.840 4.130 1.445 ;
        RECT 3.175 1.275 4.815 1.445 ;
        RECT 4.645 1.275 4.815 2.215 ;
        RECT 3.895 2.045 4.815 2.215 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.195 0.965 2.365 ;
        RECT 0.795 1.125 0.965 2.565 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 2.395 2.020 2.565 ;
        RECT 1.850 2.395 2.020 3.170 ;
        RECT 2.855 2.810 3.155 3.170 ;
        RECT 1.850 3.000 3.155 3.170 ;
        RECT 2.855 2.810 5.395 2.980 ;
        RECT 1.210 0.995 1.400 1.295 ;
        RECT 1.230 0.995 1.400 2.215 ;
        RECT 1.145 2.045 2.370 2.215 ;
        RECT 2.200 0.515 2.370 2.820 ;
        RECT 2.200 2.460 2.575 2.820 ;
        RECT 2.200 0.515 2.995 0.685 ;
        RECT 4.995 0.500 5.165 2.630 ;
        RECT 4.995 0.500 5.395 0.670 ;
        RECT 4.995 2.440 5.905 2.630 ;
        RECT 2.200 2.460 5.905 2.630 ;
        RECT 5.605 2.440 5.905 2.705 ;
        RECT 6.035 1.240 7.160 1.410 ;
        RECT 6.830 0.805 7.000 1.410 ;
        RECT 6.990 1.240 7.160 2.215 ;
        RECT 6.735 2.045 7.160 2.215 ;
        RECT 5.410 0.945 5.580 2.215 ;
        RECT 5.345 2.045 5.645 2.215 ;
        RECT 6.385 1.675 6.555 2.565 ;
        RECT 5.410 1.675 6.810 1.845 ;
        RECT 7.510 1.520 7.680 2.565 ;
        RECT 6.385 2.395 7.680 2.565 ;
  END 
END FFDQHD1XHT

MACRO FFDNSRHDMXHT
  CLASS  CORE ;
  FOREIGN FFDNSRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.890 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.605 0.550 2.060 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.540 1.060 11.715 2.430 ;
        RECT 11.540 2.070 11.790 2.430 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.440 1.125 10.970 1.295 ;
        RECT 10.760 1.125 10.970 2.280 ;
        RECT 10.440 1.980 10.970 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.655 1.330 2.050 1.785 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.380 1.580 3.850 2.035 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.825 ;
        RECT 1.655 -0.300 1.955 0.690 ;
        RECT 3.435 -0.300 3.735 1.160 ;
        RECT 6.140 -0.300 6.440 0.730 ;
        RECT 8.005 -0.300 8.305 0.730 ;
        RECT 9.930 -0.300 10.230 0.735 ;
        RECT 10.920 -0.300 11.220 0.595 ;
        RECT 0.000 -0.300 11.890 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 9.530 1.635 9.910 2.020 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.785 2.810 1.765 3.990 ;
        RECT 3.600 3.025 4.580 3.990 ;
        RECT 6.160 3.025 6.460 3.990 ;
        RECT 8.130 2.515 8.430 3.990 ;
        RECT 9.845 2.945 10.145 3.990 ;
        RECT 10.925 2.945 11.225 3.990 ;
        RECT 0.000 3.390 11.890 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.210 0.870 1.380 2.280 ;
        RECT 2.135 0.620 2.305 1.040 ;
        RECT 1.210 0.870 2.305 1.040 ;
        RECT 2.135 0.620 3.135 0.790 ;
        RECT 2.965 0.620 3.135 2.085 ;
        RECT 2.775 1.915 3.135 2.085 ;
        RECT 4.020 0.925 4.220 1.225 ;
        RECT 4.050 0.925 4.220 2.145 ;
        RECT 4.050 1.470 4.845 1.770 ;
        RECT 2.425 1.425 2.595 2.465 ;
        RECT 2.485 0.990 2.655 1.595 ;
        RECT 2.425 1.425 2.655 1.595 ;
        RECT 2.485 0.990 2.785 1.160 ;
        RECT 2.545 2.295 2.845 2.495 ;
        RECT 2.425 2.295 2.845 2.465 ;
        RECT 2.545 2.325 4.885 2.495 ;
        RECT 5.195 1.550 5.360 1.850 ;
        RECT 5.025 1.550 5.035 2.424 ;
        RECT 5.035 1.550 5.045 2.414 ;
        RECT 5.045 1.550 5.055 2.404 ;
        RECT 5.055 1.550 5.065 2.394 ;
        RECT 5.065 1.550 5.075 2.384 ;
        RECT 5.075 1.550 5.085 2.374 ;
        RECT 5.085 1.550 5.095 2.364 ;
        RECT 5.095 1.550 5.105 2.354 ;
        RECT 5.105 1.550 5.115 2.344 ;
        RECT 5.115 1.550 5.125 2.334 ;
        RECT 5.125 1.550 5.135 2.324 ;
        RECT 5.135 1.550 5.145 2.314 ;
        RECT 5.145 1.550 5.155 2.304 ;
        RECT 5.155 1.550 5.165 2.294 ;
        RECT 5.165 1.550 5.175 2.284 ;
        RECT 5.175 1.550 5.185 2.274 ;
        RECT 5.185 1.550 5.195 2.264 ;
        RECT 4.965 2.245 4.975 2.485 ;
        RECT 4.975 2.235 4.985 2.475 ;
        RECT 4.985 2.225 4.995 2.465 ;
        RECT 4.995 2.215 5.005 2.455 ;
        RECT 5.005 2.205 5.015 2.445 ;
        RECT 5.015 2.195 5.025 2.435 ;
        RECT 4.885 2.325 4.895 2.495 ;
        RECT 4.895 2.315 4.905 2.495 ;
        RECT 4.905 2.305 4.915 2.495 ;
        RECT 4.915 2.295 4.925 2.495 ;
        RECT 4.925 2.285 4.935 2.495 ;
        RECT 4.935 2.275 4.945 2.495 ;
        RECT 4.945 2.265 4.955 2.495 ;
        RECT 4.955 2.255 4.965 2.495 ;
        RECT 4.465 0.990 4.765 1.230 ;
        RECT 4.465 1.060 5.700 1.230 ;
        RECT 5.530 1.060 5.700 1.360 ;
        RECT 4.095 0.560 5.625 0.730 ;
        RECT 5.540 1.590 5.710 2.215 ;
        RECT 5.410 2.045 5.710 2.215 ;
        RECT 5.540 1.590 5.880 1.760 ;
        RECT 6.050 1.590 6.465 1.760 ;
        RECT 5.880 0.740 5.890 1.760 ;
        RECT 5.890 0.750 5.900 1.760 ;
        RECT 5.900 0.760 5.910 1.760 ;
        RECT 5.910 0.770 5.920 1.760 ;
        RECT 5.920 0.780 5.930 1.760 ;
        RECT 5.930 0.790 5.940 1.760 ;
        RECT 5.940 0.800 5.950 1.760 ;
        RECT 5.950 0.810 5.960 1.760 ;
        RECT 5.960 0.820 5.970 1.760 ;
        RECT 5.970 0.830 5.980 1.760 ;
        RECT 5.980 0.840 5.990 1.760 ;
        RECT 5.990 0.850 6.000 1.760 ;
        RECT 6.000 0.860 6.010 1.760 ;
        RECT 6.010 0.870 6.020 1.760 ;
        RECT 6.020 0.880 6.030 1.760 ;
        RECT 6.030 0.890 6.040 1.760 ;
        RECT 6.040 0.900 6.050 1.760 ;
        RECT 5.710 0.570 5.720 0.814 ;
        RECT 5.720 0.580 5.730 0.824 ;
        RECT 5.730 0.590 5.740 0.834 ;
        RECT 5.740 0.600 5.750 0.844 ;
        RECT 5.750 0.610 5.760 0.854 ;
        RECT 5.760 0.620 5.770 0.864 ;
        RECT 5.770 0.630 5.780 0.874 ;
        RECT 5.780 0.640 5.790 0.884 ;
        RECT 5.790 0.650 5.800 0.894 ;
        RECT 5.800 0.660 5.810 0.904 ;
        RECT 5.810 0.670 5.820 0.914 ;
        RECT 5.820 0.680 5.830 0.924 ;
        RECT 5.830 0.690 5.840 0.934 ;
        RECT 5.840 0.700 5.850 0.944 ;
        RECT 5.850 0.710 5.860 0.954 ;
        RECT 5.860 0.720 5.870 0.964 ;
        RECT 5.870 0.730 5.880 0.974 ;
        RECT 5.625 0.560 5.635 0.730 ;
        RECT 5.635 0.560 5.645 0.740 ;
        RECT 5.645 0.560 5.655 0.750 ;
        RECT 5.655 0.560 5.665 0.760 ;
        RECT 5.665 0.560 5.675 0.770 ;
        RECT 5.675 0.560 5.685 0.780 ;
        RECT 5.685 0.560 5.695 0.790 ;
        RECT 5.695 0.560 5.705 0.800 ;
        RECT 5.705 0.560 5.711 0.810 ;
        RECT 0.105 1.125 1.030 1.295 ;
        RECT 0.105 2.245 1.030 2.415 ;
        RECT 0.860 1.125 1.030 2.630 ;
        RECT 0.860 2.460 2.170 2.630 ;
        RECT 2.000 2.460 2.170 2.845 ;
        RECT 2.000 2.675 5.140 2.845 ;
        RECT 5.495 2.395 5.785 2.565 ;
        RECT 5.960 2.295 6.700 2.465 ;
        RECT 6.875 2.395 7.385 2.565 ;
        RECT 7.215 2.395 7.385 2.770 ;
        RECT 6.800 2.330 6.810 2.564 ;
        RECT 6.810 2.340 6.820 2.564 ;
        RECT 6.820 2.350 6.830 2.564 ;
        RECT 6.830 2.360 6.840 2.564 ;
        RECT 6.840 2.370 6.850 2.564 ;
        RECT 6.850 2.380 6.860 2.564 ;
        RECT 6.860 2.390 6.870 2.564 ;
        RECT 6.870 2.395 6.876 2.565 ;
        RECT 6.775 2.305 6.785 2.539 ;
        RECT 6.785 2.315 6.795 2.549 ;
        RECT 6.795 2.320 6.801 2.560 ;
        RECT 6.700 2.295 6.710 2.465 ;
        RECT 6.710 2.295 6.720 2.475 ;
        RECT 6.720 2.295 6.730 2.485 ;
        RECT 6.730 2.295 6.740 2.495 ;
        RECT 6.740 2.295 6.750 2.505 ;
        RECT 6.750 2.295 6.760 2.515 ;
        RECT 6.760 2.295 6.770 2.525 ;
        RECT 6.770 2.295 6.776 2.535 ;
        RECT 5.885 2.295 5.895 2.529 ;
        RECT 5.895 2.295 5.905 2.519 ;
        RECT 5.905 2.295 5.915 2.509 ;
        RECT 5.915 2.295 5.925 2.499 ;
        RECT 5.925 2.295 5.935 2.489 ;
        RECT 5.935 2.295 5.945 2.479 ;
        RECT 5.945 2.295 5.955 2.469 ;
        RECT 5.955 2.295 5.961 2.465 ;
        RECT 5.860 2.320 5.870 2.554 ;
        RECT 5.870 2.310 5.880 2.544 ;
        RECT 5.880 2.300 5.886 2.540 ;
        RECT 5.785 2.395 5.795 2.565 ;
        RECT 5.795 2.385 5.805 2.565 ;
        RECT 5.805 2.375 5.815 2.565 ;
        RECT 5.815 2.365 5.825 2.565 ;
        RECT 5.825 2.355 5.835 2.565 ;
        RECT 5.835 2.345 5.845 2.565 ;
        RECT 5.845 2.335 5.855 2.565 ;
        RECT 5.855 2.325 5.861 2.565 ;
        RECT 5.380 2.395 5.390 2.669 ;
        RECT 5.390 2.395 5.400 2.659 ;
        RECT 5.400 2.395 5.410 2.649 ;
        RECT 5.410 2.395 5.420 2.639 ;
        RECT 5.420 2.395 5.430 2.629 ;
        RECT 5.430 2.395 5.440 2.619 ;
        RECT 5.440 2.395 5.450 2.609 ;
        RECT 5.450 2.395 5.460 2.599 ;
        RECT 5.460 2.395 5.470 2.589 ;
        RECT 5.470 2.395 5.480 2.579 ;
        RECT 5.480 2.395 5.490 2.569 ;
        RECT 5.490 2.395 5.496 2.565 ;
        RECT 5.215 2.600 5.225 2.834 ;
        RECT 5.225 2.590 5.235 2.824 ;
        RECT 5.235 2.580 5.245 2.814 ;
        RECT 5.245 2.570 5.255 2.804 ;
        RECT 5.255 2.560 5.265 2.794 ;
        RECT 5.265 2.550 5.275 2.784 ;
        RECT 5.275 2.540 5.285 2.774 ;
        RECT 5.285 2.530 5.295 2.764 ;
        RECT 5.295 2.520 5.305 2.754 ;
        RECT 5.305 2.510 5.315 2.744 ;
        RECT 5.315 2.500 5.325 2.734 ;
        RECT 5.325 2.490 5.335 2.724 ;
        RECT 5.335 2.480 5.345 2.714 ;
        RECT 5.345 2.470 5.355 2.704 ;
        RECT 5.355 2.460 5.365 2.694 ;
        RECT 5.365 2.450 5.375 2.684 ;
        RECT 5.375 2.440 5.381 2.680 ;
        RECT 5.140 2.675 5.150 2.845 ;
        RECT 5.150 2.665 5.160 2.845 ;
        RECT 5.160 2.655 5.170 2.845 ;
        RECT 5.170 2.645 5.180 2.845 ;
        RECT 5.180 2.635 5.190 2.845 ;
        RECT 5.190 2.625 5.200 2.845 ;
        RECT 5.200 2.615 5.210 2.845 ;
        RECT 5.210 2.605 5.216 2.845 ;
        RECT 5.585 2.745 5.755 3.210 ;
        RECT 4.765 3.040 5.755 3.210 ;
        RECT 5.585 2.745 5.940 2.915 ;
        RECT 6.115 2.645 6.510 2.815 ;
        RECT 6.610 2.645 6.625 2.915 ;
        RECT 6.725 2.745 6.950 2.915 ;
        RECT 6.780 2.745 6.950 3.120 ;
        RECT 7.380 1.230 7.735 1.530 ;
        RECT 7.565 1.230 7.735 3.120 ;
        RECT 6.780 2.950 7.735 3.120 ;
        RECT 6.625 2.655 6.635 2.915 ;
        RECT 6.635 2.665 6.645 2.915 ;
        RECT 6.645 2.675 6.655 2.915 ;
        RECT 6.655 2.685 6.665 2.915 ;
        RECT 6.665 2.695 6.675 2.915 ;
        RECT 6.675 2.705 6.685 2.915 ;
        RECT 6.685 2.715 6.695 2.915 ;
        RECT 6.695 2.725 6.705 2.915 ;
        RECT 6.705 2.735 6.715 2.915 ;
        RECT 6.715 2.745 6.725 2.915 ;
        RECT 6.510 2.645 6.520 2.815 ;
        RECT 6.520 2.645 6.530 2.825 ;
        RECT 6.530 2.645 6.540 2.835 ;
        RECT 6.540 2.645 6.550 2.845 ;
        RECT 6.550 2.645 6.560 2.855 ;
        RECT 6.560 2.645 6.570 2.865 ;
        RECT 6.570 2.645 6.580 2.875 ;
        RECT 6.580 2.645 6.590 2.885 ;
        RECT 6.590 2.645 6.600 2.895 ;
        RECT 6.600 2.645 6.610 2.905 ;
        RECT 6.040 2.645 6.050 2.879 ;
        RECT 6.050 2.645 6.060 2.869 ;
        RECT 6.060 2.645 6.070 2.859 ;
        RECT 6.070 2.645 6.080 2.849 ;
        RECT 6.080 2.645 6.090 2.839 ;
        RECT 6.090 2.645 6.100 2.829 ;
        RECT 6.100 2.645 6.110 2.819 ;
        RECT 6.110 2.645 6.116 2.815 ;
        RECT 6.015 2.670 6.025 2.904 ;
        RECT 6.025 2.660 6.035 2.894 ;
        RECT 6.035 2.650 6.041 2.890 ;
        RECT 5.940 2.745 5.950 2.915 ;
        RECT 5.950 2.735 5.960 2.915 ;
        RECT 5.960 2.725 5.970 2.915 ;
        RECT 5.970 2.715 5.980 2.915 ;
        RECT 5.980 2.705 5.990 2.915 ;
        RECT 5.990 2.695 6.000 2.915 ;
        RECT 6.000 2.685 6.010 2.915 ;
        RECT 6.010 2.675 6.016 2.915 ;
        RECT 8.570 0.775 8.740 1.295 ;
        RECT 8.440 1.125 8.740 1.295 ;
        RECT 8.570 0.775 9.650 0.945 ;
        RECT 9.480 0.775 9.650 1.295 ;
        RECT 9.480 1.125 9.780 1.295 ;
        RECT 8.265 1.495 8.435 1.795 ;
        RECT 8.960 1.125 9.300 1.295 ;
        RECT 8.265 1.625 9.300 1.795 ;
        RECT 9.125 1.125 9.300 2.415 ;
        RECT 10.090 1.480 10.260 2.415 ;
        RECT 9.125 2.245 10.260 2.415 ;
        RECT 10.090 1.480 10.580 1.780 ;
        RECT 6.970 0.880 7.140 2.215 ;
        RECT 6.955 2.045 7.255 2.215 ;
        RECT 6.970 0.880 7.810 1.050 ;
        RECT 8.085 1.975 8.945 2.145 ;
        RECT 8.775 1.975 8.945 2.765 ;
        RECT 9.085 2.595 9.385 3.055 ;
        RECT 11.190 1.530 11.360 2.765 ;
        RECT 8.775 2.595 11.360 2.765 ;
        RECT 7.915 0.910 7.925 2.144 ;
        RECT 7.925 0.920 7.935 2.144 ;
        RECT 7.935 0.930 7.945 2.144 ;
        RECT 7.945 0.940 7.955 2.144 ;
        RECT 7.955 0.950 7.965 2.144 ;
        RECT 7.965 0.960 7.975 2.144 ;
        RECT 7.975 0.970 7.985 2.144 ;
        RECT 7.985 0.980 7.995 2.144 ;
        RECT 7.995 0.990 8.005 2.144 ;
        RECT 8.005 1.000 8.015 2.144 ;
        RECT 8.015 1.010 8.025 2.144 ;
        RECT 8.025 1.020 8.035 2.144 ;
        RECT 8.035 1.030 8.045 2.144 ;
        RECT 8.045 1.040 8.055 2.144 ;
        RECT 8.055 1.050 8.065 2.144 ;
        RECT 8.065 1.060 8.075 2.144 ;
        RECT 8.075 1.070 8.085 2.144 ;
        RECT 7.895 0.890 7.905 1.134 ;
        RECT 7.905 0.900 7.915 1.144 ;
        RECT 7.810 0.880 7.820 1.050 ;
        RECT 7.820 0.880 7.830 1.060 ;
        RECT 7.830 0.880 7.840 1.070 ;
        RECT 7.840 0.880 7.850 1.080 ;
        RECT 7.850 0.880 7.860 1.090 ;
        RECT 7.860 0.880 7.870 1.100 ;
        RECT 7.870 0.880 7.880 1.110 ;
        RECT 7.880 0.880 7.890 1.120 ;
        RECT 7.890 0.880 7.896 1.130 ;
  END 
END FFDNSRHDMXHT

MACRO FFDNSRHD2XHT
  CLASS  CORE ;
  FOREIGN FFDNSRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.940 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.350 1.525 0.720 2.015 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 12.805 1.235 13.275 1.405 ;
        RECT 12.805 0.785 13.105 1.405 ;
        RECT 12.805 2.045 13.105 2.895 ;
        RECT 13.105 1.235 13.275 2.215 ;
        RECT 12.805 2.045 13.275 2.215 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.765 0.785 12.065 1.295 ;
        RECT 11.765 1.125 12.265 1.295 ;
        RECT 12.095 1.125 12.265 2.360 ;
        RECT 11.765 2.150 12.265 2.360 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.230 2.070 1.765 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.670 1.520 3.880 1.960 ;
        RECT 3.290 1.740 3.880 1.960 ;
        RECT 3.670 1.520 4.075 1.755 ;
        RECT 3.290 1.740 4.075 1.755 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.575 -0.300 0.875 0.715 ;
        RECT 1.625 -0.300 1.925 0.700 ;
        RECT 3.565 -0.300 3.865 1.155 ;
        RECT 6.505 -0.300 6.675 1.120 ;
        RECT 8.640 -0.300 8.810 0.730 ;
        RECT 10.825 -0.300 11.465 1.055 ;
        RECT 12.285 -0.300 12.585 0.715 ;
        RECT 13.325 -0.300 13.625 1.055 ;
        RECT 0.000 -0.300 13.940 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 10.830 1.325 11.000 1.840 ;
        RECT 10.830 1.325 11.445 1.545 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.645 0.925 3.990 ;
        RECT 1.625 2.780 1.925 3.990 ;
        RECT 3.725 3.025 4.710 3.990 ;
        RECT 6.425 2.995 6.725 3.990 ;
        RECT 8.530 2.575 8.700 3.990 ;
        RECT 10.275 2.920 10.575 3.990 ;
        RECT 11.245 2.975 11.545 3.990 ;
        RECT 12.285 2.975 12.585 3.990 ;
        RECT 13.325 2.635 13.625 3.990 ;
        RECT 0.000 3.390 13.940 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.255 0.880 1.440 1.275 ;
        RECT 1.270 0.880 1.440 2.230 ;
        RECT 2.105 0.520 2.275 1.050 ;
        RECT 1.255 0.880 2.275 1.050 ;
        RECT 2.105 0.520 3.195 0.690 ;
        RECT 2.940 1.335 3.110 2.080 ;
        RECT 3.025 0.520 3.195 1.515 ;
        RECT 2.940 1.335 3.195 1.515 ;
        RECT 4.115 1.020 4.450 1.190 ;
        RECT 4.280 1.020 4.450 2.145 ;
        RECT 4.150 1.975 4.450 2.145 ;
        RECT 4.280 1.600 5.030 1.770 ;
        RECT 2.525 0.985 2.695 2.495 ;
        RECT 2.525 0.985 2.845 1.155 ;
        RECT 5.245 1.680 5.415 2.495 ;
        RECT 2.525 2.325 5.415 2.495 ;
        RECT 5.405 1.550 5.575 1.850 ;
        RECT 5.245 1.680 5.575 1.850 ;
        RECT 4.705 0.965 4.875 1.370 ;
        RECT 5.805 0.965 5.975 1.370 ;
        RECT 4.705 1.200 5.975 1.370 ;
        RECT 4.270 0.480 4.570 0.765 ;
        RECT 5.160 0.595 5.460 1.000 ;
        RECT 5.755 1.550 5.925 2.215 ;
        RECT 5.625 2.045 5.925 2.215 ;
        RECT 4.270 0.595 6.325 0.765 ;
        RECT 6.155 0.595 6.325 1.720 ;
        RECT 5.755 1.550 6.935 1.720 ;
        RECT 0.170 2.240 0.340 2.880 ;
        RECT 0.105 1.125 0.945 1.295 ;
        RECT 0.905 1.125 0.945 2.410 ;
        RECT 0.170 2.240 0.945 2.410 ;
        RECT 1.210 2.430 2.315 2.600 ;
        RECT 2.145 2.430 2.315 2.845 ;
        RECT 5.605 2.405 5.775 2.845 ;
        RECT 2.145 2.675 5.775 2.845 ;
        RECT 5.605 2.405 6.005 2.575 ;
        RECT 6.190 2.295 6.965 2.465 ;
        RECT 7.760 1.590 7.930 2.630 ;
        RECT 7.205 2.460 7.930 2.630 ;
        RECT 7.130 2.395 7.140 2.629 ;
        RECT 7.140 2.405 7.150 2.629 ;
        RECT 7.150 2.415 7.160 2.629 ;
        RECT 7.160 2.425 7.170 2.629 ;
        RECT 7.170 2.435 7.180 2.629 ;
        RECT 7.180 2.445 7.190 2.629 ;
        RECT 7.190 2.455 7.200 2.629 ;
        RECT 7.200 2.460 7.206 2.630 ;
        RECT 7.040 2.305 7.050 2.539 ;
        RECT 7.050 2.315 7.060 2.549 ;
        RECT 7.060 2.325 7.070 2.559 ;
        RECT 7.070 2.335 7.080 2.569 ;
        RECT 7.080 2.345 7.090 2.579 ;
        RECT 7.090 2.355 7.100 2.589 ;
        RECT 7.100 2.365 7.110 2.599 ;
        RECT 7.110 2.375 7.120 2.609 ;
        RECT 7.120 2.385 7.130 2.619 ;
        RECT 6.965 2.295 6.975 2.465 ;
        RECT 6.975 2.295 6.985 2.475 ;
        RECT 6.985 2.295 6.995 2.485 ;
        RECT 6.995 2.295 7.005 2.495 ;
        RECT 7.005 2.295 7.015 2.505 ;
        RECT 7.015 2.295 7.025 2.515 ;
        RECT 7.025 2.295 7.035 2.525 ;
        RECT 7.035 2.295 7.041 2.535 ;
        RECT 6.115 2.295 6.125 2.529 ;
        RECT 6.125 2.295 6.135 2.519 ;
        RECT 6.135 2.295 6.145 2.509 ;
        RECT 6.145 2.295 6.155 2.499 ;
        RECT 6.155 2.295 6.165 2.489 ;
        RECT 6.165 2.295 6.175 2.479 ;
        RECT 6.175 2.295 6.185 2.469 ;
        RECT 6.185 2.295 6.191 2.465 ;
        RECT 6.080 2.330 6.090 2.564 ;
        RECT 6.090 2.320 6.100 2.554 ;
        RECT 6.100 2.310 6.110 2.544 ;
        RECT 6.110 2.300 6.116 2.540 ;
        RECT 6.005 2.405 6.015 2.575 ;
        RECT 6.015 2.395 6.025 2.575 ;
        RECT 6.025 2.385 6.035 2.575 ;
        RECT 6.035 2.375 6.045 2.575 ;
        RECT 6.045 2.365 6.055 2.575 ;
        RECT 6.055 2.355 6.065 2.575 ;
        RECT 6.065 2.345 6.075 2.575 ;
        RECT 6.075 2.335 6.081 2.575 ;
        RECT 1.135 2.365 1.145 2.599 ;
        RECT 1.145 2.375 1.155 2.599 ;
        RECT 1.155 2.385 1.165 2.599 ;
        RECT 1.165 2.395 1.175 2.599 ;
        RECT 1.175 2.405 1.185 2.599 ;
        RECT 1.185 2.415 1.195 2.599 ;
        RECT 1.195 2.425 1.205 2.599 ;
        RECT 1.205 2.430 1.211 2.600 ;
        RECT 1.075 2.305 1.085 2.539 ;
        RECT 1.085 2.315 1.095 2.549 ;
        RECT 1.095 2.325 1.105 2.559 ;
        RECT 1.105 2.335 1.115 2.569 ;
        RECT 1.115 2.345 1.125 2.579 ;
        RECT 1.125 2.355 1.135 2.589 ;
        RECT 0.945 1.125 0.955 2.409 ;
        RECT 0.955 1.125 0.965 2.419 ;
        RECT 0.965 1.125 0.975 2.429 ;
        RECT 0.975 1.125 0.985 2.439 ;
        RECT 0.985 1.125 0.995 2.449 ;
        RECT 0.995 1.125 1.005 2.459 ;
        RECT 1.005 1.125 1.015 2.469 ;
        RECT 1.015 1.125 1.025 2.479 ;
        RECT 1.025 1.125 1.035 2.489 ;
        RECT 1.035 1.125 1.045 2.499 ;
        RECT 1.045 1.125 1.055 2.509 ;
        RECT 1.055 1.125 1.065 2.519 ;
        RECT 1.065 1.125 1.075 2.529 ;
        RECT 5.735 3.040 6.075 3.210 ;
        RECT 6.350 2.645 6.810 2.815 ;
        RECT 7.845 1.155 8.145 1.410 ;
        RECT 7.845 1.240 8.340 1.410 ;
        RECT 8.170 1.240 8.340 3.085 ;
        RECT 7.155 2.915 8.340 3.085 ;
        RECT 7.080 2.850 7.090 3.084 ;
        RECT 7.090 2.860 7.100 3.084 ;
        RECT 7.100 2.870 7.110 3.084 ;
        RECT 7.110 2.880 7.120 3.084 ;
        RECT 7.120 2.890 7.130 3.084 ;
        RECT 7.130 2.900 7.140 3.084 ;
        RECT 7.140 2.910 7.150 3.084 ;
        RECT 7.150 2.915 7.156 3.085 ;
        RECT 6.885 2.655 6.895 2.889 ;
        RECT 6.895 2.665 6.905 2.899 ;
        RECT 6.905 2.675 6.915 2.909 ;
        RECT 6.915 2.685 6.925 2.919 ;
        RECT 6.925 2.695 6.935 2.929 ;
        RECT 6.935 2.705 6.945 2.939 ;
        RECT 6.945 2.715 6.955 2.949 ;
        RECT 6.955 2.725 6.965 2.959 ;
        RECT 6.965 2.735 6.975 2.969 ;
        RECT 6.975 2.745 6.985 2.979 ;
        RECT 6.985 2.755 6.995 2.989 ;
        RECT 6.995 2.765 7.005 2.999 ;
        RECT 7.005 2.775 7.015 3.009 ;
        RECT 7.015 2.785 7.025 3.019 ;
        RECT 7.025 2.795 7.035 3.029 ;
        RECT 7.035 2.805 7.045 3.039 ;
        RECT 7.045 2.815 7.055 3.049 ;
        RECT 7.055 2.825 7.065 3.059 ;
        RECT 7.065 2.835 7.075 3.069 ;
        RECT 7.075 2.840 7.081 3.080 ;
        RECT 6.810 2.645 6.820 2.815 ;
        RECT 6.820 2.645 6.830 2.825 ;
        RECT 6.830 2.645 6.840 2.835 ;
        RECT 6.840 2.645 6.850 2.845 ;
        RECT 6.850 2.645 6.860 2.855 ;
        RECT 6.860 2.645 6.870 2.865 ;
        RECT 6.870 2.645 6.880 2.875 ;
        RECT 6.880 2.645 6.886 2.885 ;
        RECT 6.265 2.645 6.275 2.889 ;
        RECT 6.275 2.645 6.285 2.879 ;
        RECT 6.285 2.645 6.295 2.869 ;
        RECT 6.295 2.645 6.305 2.859 ;
        RECT 6.305 2.645 6.315 2.849 ;
        RECT 6.315 2.645 6.325 2.839 ;
        RECT 6.325 2.645 6.335 2.829 ;
        RECT 6.335 2.645 6.345 2.819 ;
        RECT 6.345 2.645 6.351 2.815 ;
        RECT 6.245 2.665 6.255 2.909 ;
        RECT 6.255 2.655 6.265 2.899 ;
        RECT 6.075 2.835 6.085 3.209 ;
        RECT 6.085 2.825 6.095 3.209 ;
        RECT 6.095 2.815 6.105 3.209 ;
        RECT 6.105 2.805 6.115 3.209 ;
        RECT 6.115 2.795 6.125 3.209 ;
        RECT 6.125 2.785 6.135 3.209 ;
        RECT 6.135 2.775 6.145 3.209 ;
        RECT 6.145 2.765 6.155 3.209 ;
        RECT 6.155 2.755 6.165 3.209 ;
        RECT 6.165 2.745 6.175 3.209 ;
        RECT 6.175 2.735 6.185 3.209 ;
        RECT 6.185 2.725 6.195 3.209 ;
        RECT 6.195 2.715 6.205 3.209 ;
        RECT 6.205 2.705 6.215 3.209 ;
        RECT 6.215 2.695 6.225 3.209 ;
        RECT 6.225 2.685 6.235 3.209 ;
        RECT 6.235 2.675 6.245 3.209 ;
        RECT 8.905 1.650 10.300 1.820 ;
        RECT 10.130 1.650 10.300 1.975 ;
        RECT 9.085 0.645 9.385 0.905 ;
        RECT 9.085 0.645 10.470 0.815 ;
        RECT 10.170 0.645 10.470 0.920 ;
        RECT 8.870 1.105 9.040 1.405 ;
        RECT 9.355 2.370 9.795 2.540 ;
        RECT 9.610 1.035 9.910 1.405 ;
        RECT 8.870 1.235 10.650 1.405 ;
        RECT 10.480 1.235 10.650 2.390 ;
        RECT 11.405 1.780 11.575 2.390 ;
        RECT 10.020 2.220 11.575 2.390 ;
        RECT 11.735 1.540 11.905 1.950 ;
        RECT 11.405 1.780 11.905 1.950 ;
        RECT 9.945 2.220 9.955 2.454 ;
        RECT 9.955 2.220 9.965 2.444 ;
        RECT 9.965 2.220 9.975 2.434 ;
        RECT 9.975 2.220 9.985 2.424 ;
        RECT 9.985 2.220 9.995 2.414 ;
        RECT 9.995 2.220 10.005 2.404 ;
        RECT 10.005 2.220 10.015 2.394 ;
        RECT 10.015 2.220 10.021 2.390 ;
        RECT 9.870 2.295 9.880 2.529 ;
        RECT 9.880 2.285 9.890 2.519 ;
        RECT 9.890 2.275 9.900 2.509 ;
        RECT 9.900 2.265 9.910 2.499 ;
        RECT 9.910 2.255 9.920 2.489 ;
        RECT 9.920 2.245 9.930 2.479 ;
        RECT 9.930 2.235 9.940 2.469 ;
        RECT 9.940 2.225 9.946 2.465 ;
        RECT 9.795 2.370 9.805 2.540 ;
        RECT 9.805 2.360 9.815 2.540 ;
        RECT 9.815 2.350 9.825 2.540 ;
        RECT 9.825 2.340 9.835 2.540 ;
        RECT 9.835 2.330 9.845 2.540 ;
        RECT 9.845 2.320 9.855 2.540 ;
        RECT 9.855 2.310 9.865 2.540 ;
        RECT 9.865 2.300 9.871 2.540 ;
        RECT 7.410 0.785 7.580 2.280 ;
        RECT 7.410 0.785 8.355 0.955 ;
        RECT 8.980 2.000 9.150 2.935 ;
        RECT 8.690 2.000 9.730 2.170 ;
        RECT 8.980 2.765 9.910 2.935 ;
        RECT 12.445 1.585 12.615 2.740 ;
        RECT 10.180 2.570 12.615 2.740 ;
        RECT 12.445 1.585 12.925 1.755 ;
        RECT 10.105 2.570 10.115 2.804 ;
        RECT 10.115 2.570 10.125 2.794 ;
        RECT 10.125 2.570 10.135 2.784 ;
        RECT 10.135 2.570 10.145 2.774 ;
        RECT 10.145 2.570 10.155 2.764 ;
        RECT 10.155 2.570 10.165 2.754 ;
        RECT 10.165 2.570 10.175 2.744 ;
        RECT 10.175 2.570 10.181 2.740 ;
        RECT 9.985 2.690 9.995 2.924 ;
        RECT 9.995 2.680 10.005 2.914 ;
        RECT 10.005 2.670 10.015 2.904 ;
        RECT 10.015 2.660 10.025 2.894 ;
        RECT 10.025 2.650 10.035 2.884 ;
        RECT 10.035 2.640 10.045 2.874 ;
        RECT 10.045 2.630 10.055 2.864 ;
        RECT 10.055 2.620 10.065 2.854 ;
        RECT 10.065 2.610 10.075 2.844 ;
        RECT 10.075 2.600 10.085 2.834 ;
        RECT 10.085 2.590 10.095 2.824 ;
        RECT 10.095 2.580 10.105 2.814 ;
        RECT 9.910 2.765 9.920 2.935 ;
        RECT 9.920 2.755 9.930 2.935 ;
        RECT 9.930 2.745 9.940 2.935 ;
        RECT 9.940 2.735 9.950 2.935 ;
        RECT 9.950 2.725 9.960 2.935 ;
        RECT 9.960 2.715 9.970 2.935 ;
        RECT 9.970 2.705 9.980 2.935 ;
        RECT 9.980 2.695 9.986 2.935 ;
        RECT 8.520 0.885 8.530 2.169 ;
        RECT 8.530 0.895 8.540 2.169 ;
        RECT 8.540 0.905 8.550 2.169 ;
        RECT 8.550 0.915 8.560 2.169 ;
        RECT 8.560 0.925 8.570 2.169 ;
        RECT 8.570 0.935 8.580 2.169 ;
        RECT 8.580 0.945 8.590 2.169 ;
        RECT 8.590 0.955 8.600 2.169 ;
        RECT 8.600 0.965 8.610 2.169 ;
        RECT 8.610 0.975 8.620 2.169 ;
        RECT 8.620 0.985 8.630 2.169 ;
        RECT 8.630 0.995 8.640 2.169 ;
        RECT 8.640 1.005 8.650 2.169 ;
        RECT 8.650 1.015 8.660 2.169 ;
        RECT 8.660 1.025 8.670 2.169 ;
        RECT 8.670 1.035 8.680 2.169 ;
        RECT 8.680 1.045 8.690 2.169 ;
        RECT 8.430 0.795 8.440 1.029 ;
        RECT 8.440 0.805 8.450 1.039 ;
        RECT 8.450 0.815 8.460 1.049 ;
        RECT 8.460 0.825 8.470 1.059 ;
        RECT 8.470 0.835 8.480 1.069 ;
        RECT 8.480 0.845 8.490 1.079 ;
        RECT 8.490 0.855 8.500 1.089 ;
        RECT 8.500 0.865 8.510 1.099 ;
        RECT 8.510 0.875 8.520 1.109 ;
        RECT 8.355 0.785 8.365 0.955 ;
        RECT 8.365 0.785 8.375 0.965 ;
        RECT 8.375 0.785 8.385 0.975 ;
        RECT 8.385 0.785 8.395 0.985 ;
        RECT 8.395 0.785 8.405 0.995 ;
        RECT 8.405 0.785 8.415 1.005 ;
        RECT 8.415 0.785 8.425 1.015 ;
        RECT 8.425 0.785 8.431 1.025 ;
  END 
END FFDNSRHD2XHT

MACRO FFDNSRHD1XHT
  CLASS  CORE ;
  FOREIGN FFDNSRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.300 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.350 1.670 0.720 2.015 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.955 0.720 12.200 1.360 ;
        RECT 12.030 0.720 12.125 2.960 ;
        RECT 11.955 1.980 12.125 2.960 ;
        RECT 12.030 0.720 12.200 2.480 ;
        RECT 11.955 1.980 12.200 2.480 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.760 0.785 11.255 1.295 ;
        RECT 11.085 0.785 11.255 2.215 ;
        RECT 10.850 2.045 11.255 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.675 1.320 2.135 1.750 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.495 1.375 3.665 1.950 ;
        RECT 3.315 1.740 3.665 1.950 ;
        RECT 3.495 1.375 3.935 1.545 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.575 -0.300 0.875 0.745 ;
        RECT 1.625 -0.300 1.925 0.790 ;
        RECT 3.435 -0.300 3.735 1.130 ;
        RECT 6.340 -0.300 6.510 1.325 ;
        RECT 8.525 -0.300 8.695 0.835 ;
        RECT 10.280 -0.300 10.580 0.680 ;
        RECT 11.435 -0.300 11.605 1.120 ;
        RECT 0.000 -0.300 12.300 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 9.875 1.540 10.315 1.955 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.545 0.955 3.990 ;
        RECT 1.625 2.885 1.925 3.990 ;
        RECT 3.635 2.995 4.615 3.990 ;
        RECT 6.265 2.995 6.565 3.990 ;
        RECT 8.480 2.840 9.120 3.990 ;
        RECT 10.290 2.840 10.590 3.990 ;
        RECT 11.370 2.975 11.670 3.990 ;
        RECT 0.000 3.390 12.300 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 1.055 1.295 ;
        RECT 0.885 1.125 1.055 1.575 ;
        RECT 0.895 1.520 1.075 1.585 ;
        RECT 0.105 2.195 1.055 2.365 ;
        RECT 0.885 1.510 1.065 1.575 ;
        RECT 0.905 1.520 1.075 2.364 ;
        RECT 1.235 0.970 1.440 1.360 ;
        RECT 1.270 0.970 1.440 2.340 ;
        RECT 2.105 0.500 2.275 1.140 ;
        RECT 1.235 0.970 2.275 1.140 ;
        RECT 2.105 0.500 3.195 0.670 ;
        RECT 2.900 1.355 3.070 2.090 ;
        RECT 2.835 1.920 3.135 2.090 ;
        RECT 3.025 0.500 3.195 1.525 ;
        RECT 2.900 1.355 3.195 1.525 ;
        RECT 3.955 0.960 4.285 1.130 ;
        RECT 4.115 0.960 4.285 2.110 ;
        RECT 4.115 1.520 4.345 2.110 ;
        RECT 4.045 1.940 4.345 2.110 ;
        RECT 4.115 1.520 4.880 1.820 ;
        RECT 2.455 0.960 2.625 2.460 ;
        RECT 2.455 0.960 2.845 1.130 ;
        RECT 5.085 1.680 5.255 2.460 ;
        RECT 2.455 2.290 5.255 2.460 ;
        RECT 5.240 1.550 5.410 1.850 ;
        RECT 5.085 1.680 5.410 1.850 ;
        RECT 4.465 1.020 5.800 1.190 ;
        RECT 5.630 1.020 5.800 1.325 ;
        RECT 5.015 0.560 5.315 0.840 ;
        RECT 4.095 0.560 5.315 0.730 ;
        RECT 5.590 1.535 5.760 2.215 ;
        RECT 5.460 2.045 5.760 2.215 ;
        RECT 5.015 0.670 6.160 0.840 ;
        RECT 5.990 0.670 6.160 1.705 ;
        RECT 5.590 1.535 6.815 1.705 ;
        RECT 1.140 2.535 1.310 2.835 ;
        RECT 2.105 2.535 2.275 2.810 ;
        RECT 1.140 2.535 2.275 2.705 ;
        RECT 2.325 2.645 2.625 3.085 ;
        RECT 2.135 2.645 5.590 2.815 ;
        RECT 6.015 2.295 6.880 2.465 ;
        RECT 7.705 1.810 7.875 2.565 ;
        RECT 7.055 2.395 7.875 2.565 ;
        RECT 6.980 2.330 6.990 2.564 ;
        RECT 6.990 2.340 7.000 2.564 ;
        RECT 7.000 2.350 7.010 2.564 ;
        RECT 7.010 2.360 7.020 2.564 ;
        RECT 7.020 2.370 7.030 2.564 ;
        RECT 7.030 2.380 7.040 2.564 ;
        RECT 7.040 2.390 7.050 2.564 ;
        RECT 7.050 2.395 7.056 2.565 ;
        RECT 6.955 2.305 6.965 2.539 ;
        RECT 6.965 2.315 6.975 2.549 ;
        RECT 6.975 2.320 6.981 2.560 ;
        RECT 6.880 2.295 6.890 2.465 ;
        RECT 6.890 2.295 6.900 2.475 ;
        RECT 6.900 2.295 6.910 2.485 ;
        RECT 6.910 2.295 6.920 2.495 ;
        RECT 6.920 2.295 6.930 2.505 ;
        RECT 6.930 2.295 6.940 2.515 ;
        RECT 6.940 2.295 6.950 2.525 ;
        RECT 6.950 2.295 6.956 2.535 ;
        RECT 5.940 2.295 5.950 2.529 ;
        RECT 5.950 2.295 5.960 2.519 ;
        RECT 5.960 2.295 5.970 2.509 ;
        RECT 5.970 2.295 5.980 2.499 ;
        RECT 5.980 2.295 5.990 2.489 ;
        RECT 5.990 2.295 6.000 2.479 ;
        RECT 6.000 2.295 6.010 2.469 ;
        RECT 6.010 2.295 6.016 2.465 ;
        RECT 5.665 2.570 5.675 2.804 ;
        RECT 5.675 2.560 5.685 2.794 ;
        RECT 5.685 2.550 5.695 2.784 ;
        RECT 5.695 2.540 5.705 2.774 ;
        RECT 5.705 2.530 5.715 2.764 ;
        RECT 5.715 2.520 5.725 2.754 ;
        RECT 5.725 2.510 5.735 2.744 ;
        RECT 5.735 2.500 5.745 2.734 ;
        RECT 5.745 2.490 5.755 2.724 ;
        RECT 5.755 2.480 5.765 2.714 ;
        RECT 5.765 2.470 5.775 2.704 ;
        RECT 5.775 2.460 5.785 2.694 ;
        RECT 5.785 2.450 5.795 2.684 ;
        RECT 5.795 2.440 5.805 2.674 ;
        RECT 5.805 2.430 5.815 2.664 ;
        RECT 5.815 2.420 5.825 2.654 ;
        RECT 5.825 2.410 5.835 2.644 ;
        RECT 5.835 2.400 5.845 2.634 ;
        RECT 5.845 2.390 5.855 2.624 ;
        RECT 5.855 2.380 5.865 2.614 ;
        RECT 5.865 2.370 5.875 2.604 ;
        RECT 5.875 2.360 5.885 2.594 ;
        RECT 5.885 2.350 5.895 2.584 ;
        RECT 5.895 2.340 5.905 2.574 ;
        RECT 5.905 2.330 5.915 2.564 ;
        RECT 5.915 2.320 5.925 2.554 ;
        RECT 5.925 2.310 5.935 2.544 ;
        RECT 5.935 2.300 5.941 2.540 ;
        RECT 5.590 2.645 5.600 2.815 ;
        RECT 5.600 2.635 5.610 2.815 ;
        RECT 5.610 2.625 5.620 2.815 ;
        RECT 5.620 2.615 5.630 2.815 ;
        RECT 5.630 2.605 5.640 2.815 ;
        RECT 5.640 2.595 5.650 2.815 ;
        RECT 5.650 2.585 5.660 2.815 ;
        RECT 5.660 2.575 5.666 2.815 ;
        RECT 4.805 2.995 5.105 3.210 ;
        RECT 4.805 2.995 5.915 3.165 ;
        RECT 6.185 2.645 6.650 2.815 ;
        RECT 7.675 1.270 7.975 1.630 ;
        RECT 7.675 1.460 8.225 1.630 ;
        RECT 8.055 1.460 8.225 2.915 ;
        RECT 6.825 2.745 8.225 2.915 ;
        RECT 6.750 2.680 6.760 2.914 ;
        RECT 6.760 2.690 6.770 2.914 ;
        RECT 6.770 2.700 6.780 2.914 ;
        RECT 6.780 2.710 6.790 2.914 ;
        RECT 6.790 2.720 6.800 2.914 ;
        RECT 6.800 2.730 6.810 2.914 ;
        RECT 6.810 2.740 6.820 2.914 ;
        RECT 6.820 2.745 6.826 2.915 ;
        RECT 6.725 2.655 6.735 2.889 ;
        RECT 6.735 2.665 6.745 2.899 ;
        RECT 6.745 2.670 6.751 2.910 ;
        RECT 6.650 2.645 6.660 2.815 ;
        RECT 6.660 2.645 6.670 2.825 ;
        RECT 6.670 2.645 6.680 2.835 ;
        RECT 6.680 2.645 6.690 2.845 ;
        RECT 6.690 2.645 6.700 2.855 ;
        RECT 6.700 2.645 6.710 2.865 ;
        RECT 6.710 2.645 6.720 2.875 ;
        RECT 6.720 2.645 6.726 2.885 ;
        RECT 6.095 2.645 6.105 2.895 ;
        RECT 6.105 2.645 6.115 2.885 ;
        RECT 6.115 2.645 6.125 2.875 ;
        RECT 6.125 2.645 6.135 2.865 ;
        RECT 6.135 2.645 6.145 2.855 ;
        RECT 6.145 2.645 6.155 2.845 ;
        RECT 6.155 2.645 6.165 2.835 ;
        RECT 6.165 2.645 6.175 2.825 ;
        RECT 6.175 2.645 6.185 2.815 ;
        RECT 6.085 2.655 6.095 2.905 ;
        RECT 5.915 2.825 5.925 3.165 ;
        RECT 5.925 2.815 5.935 3.165 ;
        RECT 5.935 2.805 5.945 3.165 ;
        RECT 5.945 2.795 5.955 3.165 ;
        RECT 5.955 2.785 5.965 3.165 ;
        RECT 5.965 2.775 5.975 3.165 ;
        RECT 5.975 2.765 5.985 3.165 ;
        RECT 5.985 2.755 5.995 3.165 ;
        RECT 5.995 2.745 6.005 3.165 ;
        RECT 6.005 2.735 6.015 3.165 ;
        RECT 6.015 2.725 6.025 3.165 ;
        RECT 6.025 2.715 6.035 3.165 ;
        RECT 6.035 2.705 6.045 3.165 ;
        RECT 6.045 2.695 6.055 3.165 ;
        RECT 6.055 2.685 6.065 3.165 ;
        RECT 6.065 2.675 6.075 3.165 ;
        RECT 6.075 2.665 6.085 3.165 ;
        RECT 8.980 0.760 9.150 1.280 ;
        RECT 8.850 1.110 9.150 1.280 ;
        RECT 8.980 0.760 10.060 0.930 ;
        RECT 9.890 0.760 10.060 1.280 ;
        RECT 9.890 1.110 10.190 1.280 ;
        RECT 8.755 1.460 8.925 1.760 ;
        RECT 9.370 1.110 9.670 1.630 ;
        RECT 8.755 1.460 9.670 1.630 ;
        RECT 9.500 1.110 9.670 2.305 ;
        RECT 10.495 1.520 10.665 2.305 ;
        RECT 9.500 2.135 10.665 2.305 ;
        RECT 10.495 1.520 10.905 1.820 ;
        RECT 7.225 0.900 7.395 2.215 ;
        RECT 7.225 2.045 7.525 2.215 ;
        RECT 7.225 0.900 8.325 1.070 ;
        RECT 8.155 0.900 8.325 1.280 ;
        RECT 8.155 1.110 8.575 1.280 ;
        RECT 8.405 1.110 8.575 2.660 ;
        RECT 9.560 2.490 9.860 2.985 ;
        RECT 11.485 1.585 11.655 2.660 ;
        RECT 8.405 2.490 11.655 2.660 ;
        RECT 11.485 1.585 11.850 1.755 ;
  END 
END FFDNSRHD1XHT

MACRO FFDNSHDMXHT
  CLASS  CORE ;
  FOREIGN FFDNSHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.430 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.090 1.060 9.330 1.360 ;
        RECT 9.120 1.060 9.330 2.435 ;
        RECT 9.090 1.980 9.330 2.435 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.050 1.060 8.220 1.360 ;
        RECT 8.050 1.190 8.510 1.360 ;
        RECT 8.300 1.190 8.510 2.240 ;
        RECT 7.985 2.070 8.510 2.240 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.560 1.495 1.950 2.050 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 0.530 ;
        RECT 1.475 -0.300 1.775 0.530 ;
        RECT 3.375 -0.300 3.675 1.020 ;
        RECT 4.570 -0.300 4.870 0.595 ;
        RECT 6.620 -0.300 6.790 0.720 ;
        RECT 8.535 -0.300 8.835 0.595 ;
        RECT 0.000 -0.300 9.430 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.115 0.755 4.415 0.945 ;
        RECT 5.185 0.605 5.355 0.945 ;
        RECT 4.115 0.775 5.355 0.945 ;
        RECT 5.185 0.605 6.375 0.775 ;
        RECT 6.205 0.605 6.375 1.145 ;
        RECT 7.005 0.920 7.360 1.145 ;
        RECT 7.190 0.540 7.360 1.145 ;
        RECT 6.205 0.975 7.360 1.145 ;
        RECT 7.190 0.540 7.595 0.710 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.610 0.955 3.990 ;
        RECT 1.440 2.580 1.610 3.990 ;
        RECT 3.395 3.160 3.695 3.990 ;
        RECT 4.570 3.160 4.870 3.990 ;
        RECT 6.575 2.770 6.875 3.990 ;
        RECT 7.215 2.945 7.515 3.990 ;
        RECT 8.535 2.975 8.835 3.990 ;
        RECT 0.000 3.390 9.430 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.490 0.830 2.660 1.130 ;
        RECT 2.490 0.960 2.895 1.130 ;
        RECT 2.610 1.980 2.780 2.280 ;
        RECT 2.725 0.960 2.895 2.150 ;
        RECT 2.610 1.980 2.895 2.150 ;
        RECT 2.725 1.675 3.895 1.845 ;
        RECT 3.115 1.245 4.245 1.415 ;
        RECT 4.075 1.125 4.245 2.215 ;
        RECT 3.945 2.045 4.245 2.215 ;
        RECT 4.075 1.125 5.135 1.295 ;
        RECT 1.150 1.060 1.380 1.360 ;
        RECT 1.210 1.060 1.380 2.400 ;
        RECT 1.150 1.980 1.380 2.400 ;
        RECT 1.150 2.230 1.960 2.400 ;
        RECT 1.790 2.230 1.960 2.980 ;
        RECT 1.790 2.810 5.515 2.980 ;
        RECT 0.105 0.655 0.405 0.880 ;
        RECT 0.225 2.195 0.405 2.935 ;
        RECT 0.105 2.765 0.405 2.935 ;
        RECT 0.795 0.710 0.965 2.365 ;
        RECT 0.225 2.195 0.965 2.365 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.105 0.710 2.310 0.880 ;
        RECT 2.140 0.480 2.310 2.630 ;
        RECT 2.140 1.685 2.400 1.985 ;
        RECT 2.140 0.480 2.935 0.650 ;
        RECT 5.340 1.645 5.510 2.630 ;
        RECT 5.380 1.245 5.550 1.815 ;
        RECT 5.340 1.645 5.550 1.815 ;
        RECT 2.140 2.460 6.255 2.630 ;
        RECT 6.445 1.325 7.710 1.495 ;
        RECT 7.540 0.890 7.710 2.215 ;
        RECT 7.125 2.045 7.710 2.215 ;
        RECT 7.540 1.540 8.120 1.840 ;
        RECT 5.775 0.955 5.945 2.215 ;
        RECT 5.685 0.955 5.985 1.125 ;
        RECT 5.690 2.045 5.990 2.215 ;
        RECT 6.480 1.675 6.650 2.590 ;
        RECT 5.775 1.675 7.225 1.845 ;
        RECT 8.740 1.530 8.910 2.590 ;
        RECT 6.480 2.420 8.910 2.590 ;
        RECT 8.740 1.530 8.920 1.830 ;
  END 
END FFDNSHDMXHT

MACRO FFDNSHDLXHT
  CLASS  CORE ;
  FOREIGN FFDNSHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.430 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.090 1.060 9.330 1.360 ;
        RECT 9.120 1.060 9.330 2.435 ;
        RECT 9.090 1.980 9.330 2.435 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.050 1.060 8.220 1.360 ;
        RECT 8.050 1.190 8.510 1.360 ;
        RECT 8.300 1.190 8.510 2.240 ;
        RECT 7.985 2.070 8.510 2.240 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.620 1.495 2.010 2.050 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.530 ;
        RECT 1.535 -0.300 1.835 0.530 ;
        RECT 3.435 -0.300 3.735 1.020 ;
        RECT 4.570 -0.300 4.870 0.595 ;
        RECT 6.590 -0.300 6.760 0.760 ;
        RECT 8.535 -0.300 8.835 0.745 ;
        RECT 0.000 -0.300 9.430 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.175 0.775 5.355 0.925 ;
        RECT 4.180 0.755 4.475 0.945 ;
        RECT 4.175 0.755 4.475 0.925 ;
        RECT 5.185 0.605 5.355 0.945 ;
        RECT 4.180 0.775 5.355 0.945 ;
        RECT 5.185 0.605 6.375 0.775 ;
        RECT 6.205 0.605 6.375 1.145 ;
        RECT 7.005 0.920 7.360 1.145 ;
        RECT 7.190 0.540 7.360 1.145 ;
        RECT 6.205 0.975 7.360 1.145 ;
        RECT 7.190 0.540 7.565 0.710 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.685 2.580 0.985 3.990 ;
        RECT 1.495 2.580 1.665 3.990 ;
        RECT 3.485 3.160 3.785 3.990 ;
        RECT 4.600 3.160 4.900 3.990 ;
        RECT 6.575 2.770 6.875 3.990 ;
        RECT 7.155 2.875 7.455 3.990 ;
        RECT 8.535 2.770 8.835 3.990 ;
        RECT 0.000 3.390 9.430 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.550 0.915 2.885 1.130 ;
        RECT 2.550 0.830 2.720 1.130 ;
        RECT 2.715 0.915 2.885 2.280 ;
        RECT 2.660 1.980 2.885 2.280 ;
        RECT 2.715 1.675 3.965 1.845 ;
        RECT 3.175 1.245 4.335 1.415 ;
        RECT 4.165 1.245 4.335 2.215 ;
        RECT 4.035 2.045 4.335 2.215 ;
        RECT 4.170 1.125 5.135 1.295 ;
        RECT 1.210 1.060 1.420 1.360 ;
        RECT 1.250 1.060 1.420 2.400 ;
        RECT 1.210 1.990 1.420 2.400 ;
        RECT 1.210 2.230 2.020 2.400 ;
        RECT 1.850 2.230 2.020 2.980 ;
        RECT 1.850 2.810 5.675 2.980 ;
        RECT 0.105 1.125 1.010 1.295 ;
        RECT 0.840 0.710 1.010 2.365 ;
        RECT 0.105 2.195 1.010 2.365 ;
        RECT 0.840 1.525 1.070 1.825 ;
        RECT 0.840 0.710 2.370 0.880 ;
        RECT 2.200 0.480 2.370 2.630 ;
        RECT 2.200 1.685 2.460 1.985 ;
        RECT 2.200 0.480 3.025 0.650 ;
        RECT 5.380 1.245 5.550 2.630 ;
        RECT 2.200 2.460 6.255 2.630 ;
        RECT 6.415 1.325 7.710 1.495 ;
        RECT 7.540 0.890 7.710 2.215 ;
        RECT 7.155 2.045 7.710 2.215 ;
        RECT 7.540 1.540 8.120 1.840 ;
        RECT 5.755 0.955 5.925 2.280 ;
        RECT 5.685 0.955 5.990 1.125 ;
        RECT 6.805 1.675 6.975 2.590 ;
        RECT 5.755 1.675 7.225 1.845 ;
        RECT 8.740 1.525 8.910 2.590 ;
        RECT 6.805 2.420 8.910 2.590 ;
        RECT 8.740 1.525 8.920 1.825 ;
  END 
END FFDNSHDLXHT

MACRO FFDNSHD2XHT
  CLASS  CORE ;
  FOREIGN FFDNSHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.070 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.210 0.720 10.380 2.960 ;
        RECT 10.210 1.665 10.560 2.015 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.120 0.720 9.340 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.560 1.265 1.950 1.900 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.545 -0.300 0.845 0.530 ;
        RECT 1.495 -0.300 1.795 0.530 ;
        RECT 3.395 -0.300 3.695 1.020 ;
        RECT 4.915 -0.300 5.215 0.715 ;
        RECT 7.080 -0.300 7.380 0.740 ;
        RECT 8.585 -0.300 8.885 1.055 ;
        RECT 9.625 -0.300 9.925 1.055 ;
        RECT 10.665 -0.300 10.965 1.055 ;
        RECT 0.000 -0.300 11.070 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.700 1.240 4.870 1.565 ;
        RECT 4.985 0.960 5.165 1.410 ;
        RECT 4.700 1.240 5.165 1.410 ;
        RECT 5.395 0.605 5.565 1.130 ;
        RECT 4.985 0.960 5.565 1.130 ;
        RECT 5.395 0.605 6.725 0.775 ;
        RECT 6.555 0.605 6.725 1.145 ;
        RECT 7.770 0.920 7.940 1.845 ;
        RECT 7.415 0.920 7.960 1.145 ;
        RECT 6.555 0.975 7.960 1.145 ;
        RECT 7.770 1.675 8.120 1.845 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.645 0.925 3.990 ;
        RECT 1.535 2.555 1.705 3.990 ;
        RECT 3.395 3.095 3.695 3.990 ;
        RECT 4.550 3.095 5.190 3.990 ;
        RECT 6.965 2.790 7.265 3.990 ;
        RECT 8.075 2.790 8.375 3.990 ;
        RECT 8.585 2.975 8.885 3.990 ;
        RECT 9.625 2.975 9.925 3.990 ;
        RECT 10.665 2.295 10.965 3.990 ;
        RECT 0.000 3.390 11.070 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.510 0.960 2.845 1.130 ;
        RECT 2.510 0.830 2.680 1.130 ;
        RECT 2.675 0.960 2.845 2.215 ;
        RECT 2.595 2.045 2.895 2.215 ;
        RECT 2.675 1.675 3.925 1.845 ;
        RECT 3.135 1.245 4.485 1.415 ;
        RECT 4.315 0.850 4.485 2.215 ;
        RECT 3.945 2.045 4.485 2.215 ;
        RECT 4.315 0.850 4.645 1.020 ;
        RECT 5.195 1.610 5.365 1.915 ;
        RECT 4.315 1.745 5.365 1.915 ;
        RECT 1.160 1.060 1.380 1.360 ;
        RECT 1.210 1.060 1.380 2.335 ;
        RECT 1.160 1.980 1.380 2.335 ;
        RECT 1.160 2.165 2.055 2.335 ;
        RECT 1.885 2.165 2.055 2.915 ;
        RECT 2.905 2.745 3.205 2.970 ;
        RECT 1.885 2.745 6.010 2.915 ;
        RECT 5.830 2.745 6.010 3.185 ;
        RECT 5.830 3.015 6.450 3.185 ;
        RECT 0.170 2.195 0.340 2.880 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.795 0.710 0.965 2.365 ;
        RECT 0.170 2.195 0.965 2.365 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 0.710 2.330 0.880 ;
        RECT 2.160 0.480 2.330 1.985 ;
        RECT 2.235 1.685 2.405 2.565 ;
        RECT 2.160 1.685 2.420 1.985 ;
        RECT 2.160 0.480 2.955 0.650 ;
        RECT 5.675 1.290 5.845 2.565 ;
        RECT 2.235 2.395 6.540 2.565 ;
        RECT 6.370 2.395 6.540 2.770 ;
        RECT 8.140 1.060 8.310 1.495 ;
        RECT 8.140 1.325 8.940 1.495 ;
        RECT 8.770 1.325 8.940 2.215 ;
        RECT 7.525 2.045 8.940 2.215 ;
        RECT 6.165 0.955 6.335 2.215 ;
        RECT 6.075 0.955 6.375 1.125 ;
        RECT 6.100 2.045 6.400 2.215 ;
        RECT 7.175 1.610 7.345 2.610 ;
        RECT 6.165 1.610 7.590 1.780 ;
        RECT 8.570 2.440 8.815 2.630 ;
        RECT 7.175 2.440 8.815 2.610 ;
        RECT 9.860 1.530 10.030 2.630 ;
        RECT 8.570 2.460 10.030 2.630 ;
  END 
END FFDNSHD2XHT

MACRO FFDNSHD1XHT
  CLASS  CORE ;
  FOREIGN FFDNSHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.430 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.090 0.720 9.330 1.360 ;
        RECT 9.120 0.720 9.330 2.960 ;
        RECT 9.090 1.980 9.330 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.050 0.720 8.220 1.360 ;
        RECT 8.050 1.190 8.510 1.360 ;
        RECT 8.300 1.190 8.510 2.240 ;
        RECT 7.985 2.070 8.510 2.240 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.560 1.495 1.950 2.050 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.530 ;
        RECT 1.475 -0.300 1.775 0.530 ;
        RECT 3.365 -0.300 3.665 1.020 ;
        RECT 4.570 -0.300 4.870 0.595 ;
        RECT 6.620 -0.300 6.790 0.640 ;
        RECT 8.505 -0.300 8.805 0.715 ;
        RECT 0.000 -0.300 9.430 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.105 0.705 4.405 0.945 ;
        RECT 5.185 0.605 5.355 0.945 ;
        RECT 4.105 0.775 5.355 0.945 ;
        RECT 5.185 0.605 6.375 0.775 ;
        RECT 6.205 0.605 6.375 1.130 ;
        RECT 7.190 0.535 7.360 1.130 ;
        RECT 6.205 0.920 7.360 1.130 ;
        RECT 7.190 0.535 7.595 0.705 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.645 0.955 3.990 ;
        RECT 1.440 2.580 1.610 3.990 ;
        RECT 3.395 3.160 3.695 3.990 ;
        RECT 4.570 3.160 4.870 3.990 ;
        RECT 6.575 2.770 6.875 3.990 ;
        RECT 7.215 3.005 7.515 3.990 ;
        RECT 8.505 2.975 8.805 3.990 ;
        RECT 0.000 3.390 9.430 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.490 0.960 2.825 1.130 ;
        RECT 2.490 0.830 2.660 1.130 ;
        RECT 2.610 1.980 2.780 2.280 ;
        RECT 2.655 0.960 2.825 2.215 ;
        RECT 2.610 1.980 2.825 2.215 ;
        RECT 2.655 1.675 3.895 1.845 ;
        RECT 3.115 1.245 4.245 1.415 ;
        RECT 4.075 1.125 4.245 2.215 ;
        RECT 3.945 2.045 4.245 2.215 ;
        RECT 4.075 1.125 5.135 1.295 ;
        RECT 1.150 1.060 1.380 1.360 ;
        RECT 1.210 1.060 1.380 2.400 ;
        RECT 1.150 1.980 1.380 2.400 ;
        RECT 1.150 2.230 1.960 2.400 ;
        RECT 1.790 2.230 1.960 2.980 ;
        RECT 1.790 2.810 5.675 2.980 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.795 0.710 0.965 2.465 ;
        RECT 0.105 2.295 0.965 2.465 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 0.710 2.310 0.880 ;
        RECT 2.140 0.480 2.310 2.630 ;
        RECT 2.140 1.685 2.400 1.985 ;
        RECT 2.140 0.480 2.935 0.650 ;
        RECT 5.255 1.645 5.425 2.630 ;
        RECT 5.380 1.245 5.550 1.815 ;
        RECT 5.255 1.645 5.550 1.815 ;
        RECT 2.140 2.460 6.255 2.630 ;
        RECT 5.955 2.460 6.255 2.705 ;
        RECT 6.445 1.325 7.710 1.495 ;
        RECT 7.540 0.890 7.710 2.215 ;
        RECT 7.125 2.045 7.710 2.215 ;
        RECT 7.540 1.540 8.120 1.840 ;
        RECT 5.685 0.955 5.990 1.125 ;
        RECT 5.820 0.955 5.990 2.215 ;
        RECT 5.690 2.045 5.990 2.215 ;
        RECT 6.480 1.675 6.650 2.590 ;
        RECT 5.820 1.675 7.225 1.845 ;
        RECT 8.740 1.555 8.910 2.590 ;
        RECT 6.480 2.420 8.910 2.590 ;
        RECT 8.740 1.555 8.920 1.855 ;
  END 
END FFDNSHD1XHT

MACRO FFDNRHDMXHT
  CLASS  CORE ;
  FOREIGN FFDNRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.590 2.010 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.220 1.060 10.560 1.360 ;
        RECT 10.350 1.060 10.560 2.440 ;
        RECT 10.220 1.980 10.560 2.440 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.120 0.855 9.370 1.470 ;
        RECT 9.120 1.300 9.690 1.470 ;
        RECT 9.520 1.300 9.690 2.215 ;
        RECT 9.115 2.045 9.690 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.640 1.270 2.030 1.775 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.430 1.610 5.925 2.010 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.530 ;
        RECT 1.575 -0.300 1.875 0.530 ;
        RECT 3.505 -0.300 3.805 1.020 ;
        RECT 4.495 -0.300 4.795 0.595 ;
        RECT 5.565 -0.300 5.735 0.810 ;
        RECT 7.475 -0.300 7.775 0.595 ;
        RECT 8.635 -0.300 8.935 0.595 ;
        RECT 9.665 -0.300 9.965 0.595 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.605 0.955 3.990 ;
        RECT 1.540 2.490 1.710 3.990 ;
        RECT 3.475 3.195 3.775 3.990 ;
        RECT 5.605 3.195 5.905 3.990 ;
        RECT 7.605 2.810 7.905 3.990 ;
        RECT 9.605 2.925 9.905 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.590 1.190 2.850 1.390 ;
        RECT 2.590 0.830 2.760 1.390 ;
        RECT 2.680 1.190 2.850 2.305 ;
        RECT 2.680 1.675 3.975 1.845 ;
        RECT 3.245 1.245 4.325 1.415 ;
        RECT 4.120 0.775 4.290 1.415 ;
        RECT 4.155 1.245 4.325 2.215 ;
        RECT 4.155 2.045 4.695 2.215 ;
        RECT 4.980 0.480 5.150 0.945 ;
        RECT 4.120 0.775 5.150 0.945 ;
        RECT 1.250 1.060 1.440 1.360 ;
        RECT 1.270 1.060 1.440 2.280 ;
        RECT 1.250 1.980 1.440 2.280 ;
        RECT 1.250 2.110 2.060 2.280 ;
        RECT 1.890 2.110 2.060 3.015 ;
        RECT 5.900 2.745 6.070 3.015 ;
        RECT 1.890 2.845 6.070 3.015 ;
        RECT 5.900 2.745 6.645 2.915 ;
        RECT 0.105 1.125 1.005 1.295 ;
        RECT 0.835 0.710 1.005 2.360 ;
        RECT 0.105 2.190 1.005 2.360 ;
        RECT 0.835 1.525 1.070 1.825 ;
        RECT 0.835 0.710 2.410 0.880 ;
        RECT 2.240 0.480 2.410 2.665 ;
        RECT 2.240 1.655 2.500 1.955 ;
        RECT 2.240 0.480 3.065 0.650 ;
        RECT 5.545 2.395 5.715 2.665 ;
        RECT 2.240 2.495 5.715 2.665 ;
        RECT 6.285 1.330 6.455 2.565 ;
        RECT 6.265 1.330 6.565 1.500 ;
        RECT 5.545 2.395 7.225 2.565 ;
        RECT 6.925 2.395 7.225 2.595 ;
        RECT 4.505 1.675 5.250 1.845 ;
        RECT 5.080 1.125 5.250 2.280 ;
        RECT 5.915 0.605 6.085 1.295 ;
        RECT 5.055 1.125 6.085 1.295 ;
        RECT 7.095 0.605 7.265 0.945 ;
        RECT 5.915 0.605 7.265 0.775 ;
        RECT 7.095 0.775 8.775 0.945 ;
        RECT 8.605 0.775 8.775 1.515 ;
        RECT 8.055 1.125 8.425 1.495 ;
        RECT 7.295 1.325 8.425 1.495 ;
        RECT 8.255 1.125 8.425 1.865 ;
        RECT 8.590 1.695 8.760 2.280 ;
        RECT 9.040 1.675 9.340 1.865 ;
        RECT 8.255 1.695 9.340 1.865 ;
        RECT 6.555 0.955 6.915 1.125 ;
        RECT 6.745 0.955 6.915 2.215 ;
        RECT 6.660 2.045 6.960 2.215 ;
        RECT 6.745 1.675 8.075 1.845 ;
        RECT 7.905 1.675 8.075 2.630 ;
        RECT 9.870 1.525 10.040 2.630 ;
        RECT 7.905 2.460 10.040 2.630 ;
  END 
END FFDNRHDMXHT

MACRO FFDNRHDLXHT
  CLASS  CORE ;
  FOREIGN FFDNRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.590 2.010 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.220 1.060 10.560 1.360 ;
        RECT 10.350 1.060 10.560 2.445 ;
        RECT 10.220 1.980 10.560 2.445 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.120 0.855 9.370 1.470 ;
        RECT 9.120 1.300 9.690 1.470 ;
        RECT 9.520 1.300 9.690 2.215 ;
        RECT 9.115 2.045 9.690 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.640 1.270 2.030 1.775 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.430 1.610 5.925 2.010 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.685 -0.300 0.985 0.530 ;
        RECT 1.575 -0.300 1.875 0.530 ;
        RECT 3.505 -0.300 3.805 1.020 ;
        RECT 4.495 -0.300 4.795 0.595 ;
        RECT 5.565 -0.300 5.735 0.810 ;
        RECT 7.505 -0.300 7.805 0.595 ;
        RECT 8.605 -0.300 8.905 0.595 ;
        RECT 9.665 -0.300 9.965 0.745 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.685 2.540 0.985 3.990 ;
        RECT 1.540 2.490 1.710 3.990 ;
        RECT 3.505 3.195 3.805 3.990 ;
        RECT 5.605 3.195 5.905 3.990 ;
        RECT 7.605 2.810 7.905 3.990 ;
        RECT 9.605 2.810 9.905 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.590 1.190 2.850 1.390 ;
        RECT 2.590 0.830 2.760 1.390 ;
        RECT 2.680 1.190 2.850 2.305 ;
        RECT 2.680 1.675 3.975 1.845 ;
        RECT 3.245 1.245 4.325 1.415 ;
        RECT 4.150 0.775 4.320 1.415 ;
        RECT 4.155 1.245 4.325 2.215 ;
        RECT 4.155 2.045 4.725 2.215 ;
        RECT 5.010 0.480 5.180 0.945 ;
        RECT 4.150 0.775 5.180 0.945 ;
        RECT 1.250 1.060 1.440 1.360 ;
        RECT 1.270 1.060 1.440 2.280 ;
        RECT 1.250 1.980 1.440 2.280 ;
        RECT 1.250 2.110 2.060 2.280 ;
        RECT 1.890 2.110 2.060 3.015 ;
        RECT 5.900 2.745 6.070 3.015 ;
        RECT 1.890 2.845 6.070 3.015 ;
        RECT 5.900 2.745 6.645 2.915 ;
        RECT 0.105 1.125 1.005 1.295 ;
        RECT 0.835 0.710 1.005 2.360 ;
        RECT 0.105 2.190 1.005 2.360 ;
        RECT 0.835 1.525 1.070 1.825 ;
        RECT 0.835 0.710 2.410 0.880 ;
        RECT 2.240 0.480 2.410 2.665 ;
        RECT 2.240 1.655 2.500 1.955 ;
        RECT 2.240 0.480 3.065 0.650 ;
        RECT 5.545 2.395 5.715 2.665 ;
        RECT 2.240 2.495 5.715 2.665 ;
        RECT 6.265 1.330 6.435 2.565 ;
        RECT 6.265 1.330 6.565 1.500 ;
        RECT 5.545 2.395 7.225 2.565 ;
        RECT 6.925 2.395 7.225 2.585 ;
        RECT 4.505 1.590 5.250 1.760 ;
        RECT 5.080 1.125 5.250 2.280 ;
        RECT 5.915 0.605 6.085 1.295 ;
        RECT 5.055 1.125 6.085 1.295 ;
        RECT 7.130 0.605 7.300 0.945 ;
        RECT 5.915 0.605 7.300 0.775 ;
        RECT 7.130 0.775 8.775 0.945 ;
        RECT 8.605 0.775 8.775 1.515 ;
        RECT 8.055 1.125 8.425 1.495 ;
        RECT 7.295 1.325 8.425 1.495 ;
        RECT 8.255 1.125 8.425 1.865 ;
        RECT 8.590 1.695 8.760 2.280 ;
        RECT 9.040 1.675 9.340 1.865 ;
        RECT 8.255 1.695 9.340 1.865 ;
        RECT 6.555 0.955 6.915 1.125 ;
        RECT 6.745 0.955 6.915 2.215 ;
        RECT 6.660 2.045 6.960 2.215 ;
        RECT 6.745 1.675 8.075 1.845 ;
        RECT 7.905 1.675 8.075 2.630 ;
        RECT 9.870 1.530 10.040 2.630 ;
        RECT 7.905 2.460 10.040 2.630 ;
  END 
END FFDNRHDLXHT

MACRO FFDNRHD2XHT
  CLASS  CORE ;
  FOREIGN FFDNRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.480 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.620 0.720 10.790 2.960 ;
        RECT 10.620 1.655 10.970 2.015 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.530 0.720 9.750 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.580 1.270 1.965 1.765 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.360 1.565 6.050 1.735 ;
        RECT 5.680 1.565 6.050 2.130 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.575 -0.300 0.875 0.500 ;
        RECT 1.515 -0.300 1.815 0.500 ;
        RECT 3.435 -0.300 3.735 1.020 ;
        RECT 4.505 -0.300 4.805 0.595 ;
        RECT 5.610 -0.300 5.910 0.715 ;
        RECT 7.510 -0.300 7.810 0.595 ;
        RECT 8.995 -0.300 9.295 1.055 ;
        RECT 10.035 -0.300 10.335 1.055 ;
        RECT 11.075 -0.300 11.375 1.055 ;
        RECT 0.000 -0.300 11.480 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.645 0.925 3.990 ;
        RECT 1.480 2.525 1.650 3.990 ;
        RECT 3.450 3.140 3.750 3.990 ;
        RECT 5.610 3.095 5.910 3.990 ;
        RECT 7.620 2.910 7.920 3.990 ;
        RECT 8.995 2.975 9.295 3.990 ;
        RECT 10.035 2.975 10.335 3.990 ;
        RECT 11.075 2.295 11.375 3.990 ;
        RECT 0.000 3.390 11.480 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.530 1.085 2.855 1.285 ;
        RECT 2.530 0.885 2.700 1.285 ;
        RECT 2.685 1.085 2.855 2.260 ;
        RECT 2.530 2.090 2.855 2.260 ;
        RECT 2.685 1.675 3.915 1.845 ;
        RECT 3.185 1.245 4.265 1.415 ;
        RECT 4.020 0.735 4.190 1.415 ;
        RECT 4.095 1.245 4.265 2.215 ;
        RECT 4.095 2.045 4.715 2.215 ;
        RECT 4.985 0.480 5.155 0.945 ;
        RECT 4.020 0.775 5.155 0.945 ;
        RECT 1.190 1.060 1.380 1.360 ;
        RECT 1.210 1.060 1.380 2.280 ;
        RECT 1.190 1.980 1.380 2.280 ;
        RECT 1.190 2.090 2.000 2.280 ;
        RECT 1.830 2.090 2.000 2.960 ;
        RECT 2.835 2.790 3.135 2.975 ;
        RECT 5.190 2.745 5.360 2.960 ;
        RECT 1.830 2.790 5.360 2.960 ;
        RECT 5.190 2.745 6.480 2.915 ;
        RECT 6.310 2.745 6.480 3.210 ;
        RECT 6.310 3.040 7.140 3.210 ;
        RECT 0.170 2.195 0.340 2.835 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.795 0.710 0.965 2.390 ;
        RECT 0.170 2.195 0.965 2.390 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 0.710 2.350 0.880 ;
        RECT 2.180 0.480 2.350 2.610 ;
        RECT 2.180 1.720 2.505 1.890 ;
        RECT 2.180 0.480 3.005 0.650 ;
        RECT 4.835 2.395 5.005 2.610 ;
        RECT 2.180 2.440 5.005 2.610 ;
        RECT 6.270 1.355 6.440 2.565 ;
        RECT 6.270 1.355 6.570 1.525 ;
        RECT 4.835 2.395 7.165 2.565 ;
        RECT 6.995 2.395 7.165 2.795 ;
        RECT 4.445 1.575 5.160 1.745 ;
        RECT 4.990 1.125 5.160 2.215 ;
        RECT 4.990 2.045 5.320 2.215 ;
        RECT 5.560 0.960 5.730 1.295 ;
        RECT 4.990 1.125 5.730 1.295 ;
        RECT 5.560 0.960 6.320 1.130 ;
        RECT 6.150 0.635 6.320 1.130 ;
        RECT 7.145 0.635 7.315 0.945 ;
        RECT 6.150 0.635 7.315 0.805 ;
        RECT 7.145 0.775 8.780 0.945 ;
        RECT 8.610 0.775 8.780 1.735 ;
        RECT 8.060 1.125 8.430 1.495 ;
        RECT 7.250 1.325 8.430 1.495 ;
        RECT 8.260 1.125 8.430 2.240 ;
        RECT 9.180 1.525 9.350 2.240 ;
        RECT 8.260 2.070 9.350 2.240 ;
        RECT 6.560 0.985 6.965 1.155 ;
        RECT 6.795 0.985 6.965 2.215 ;
        RECT 6.665 2.045 6.965 2.215 ;
        RECT 6.795 1.675 8.080 1.845 ;
        RECT 7.910 1.675 8.080 2.655 ;
        RECT 10.270 1.520 10.440 2.655 ;
        RECT 7.910 2.485 10.440 2.655 ;
  END 
END FFDNRHD2XHT

MACRO FFDNRHD1XHT
  CLASS  CORE ;
  FOREIGN FFDNRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.010 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.180 0.720 10.560 1.360 ;
        RECT 10.350 0.720 10.560 2.960 ;
        RECT 10.180 1.980 10.560 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.120 1.300 9.650 1.345 ;
        RECT 9.125 0.720 9.330 1.470 ;
        RECT 9.120 0.720 9.330 1.345 ;
        RECT 9.125 1.300 9.650 1.470 ;
        RECT 9.480 1.300 9.650 2.280 ;
        RECT 9.075 2.110 9.650 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.600 1.270 1.990 1.795 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.430 1.610 5.885 2.010 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.530 ;
        RECT 1.535 -0.300 1.835 0.530 ;
        RECT 3.435 -0.300 3.735 1.020 ;
        RECT 4.455 -0.300 4.755 0.595 ;
        RECT 5.525 -0.300 5.695 0.810 ;
        RECT 7.435 -0.300 7.735 0.495 ;
        RECT 8.565 -0.300 8.865 0.480 ;
        RECT 9.595 -0.300 9.895 1.055 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.605 0.955 3.990 ;
        RECT 1.500 2.525 1.670 3.990 ;
        RECT 3.435 3.195 3.735 3.990 ;
        RECT 5.565 3.195 5.865 3.990 ;
        RECT 7.565 2.810 7.865 3.990 ;
        RECT 9.595 2.975 9.895 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.550 1.190 2.810 1.390 ;
        RECT 2.550 0.830 2.720 1.390 ;
        RECT 2.640 1.190 2.810 2.305 ;
        RECT 2.640 1.675 3.935 1.845 ;
        RECT 3.205 1.245 4.285 1.415 ;
        RECT 4.050 0.775 4.220 1.415 ;
        RECT 4.115 1.245 4.285 2.240 ;
        RECT 4.115 2.070 4.655 2.240 ;
        RECT 4.940 0.480 5.110 0.945 ;
        RECT 4.050 0.775 5.110 0.945 ;
        RECT 1.210 1.060 1.400 1.360 ;
        RECT 1.230 1.060 1.400 2.280 ;
        RECT 1.210 1.980 1.400 2.280 ;
        RECT 1.210 2.110 2.020 2.280 ;
        RECT 1.850 2.110 2.020 3.015 ;
        RECT 5.860 2.745 6.030 3.015 ;
        RECT 1.850 2.845 6.030 3.015 ;
        RECT 5.860 2.745 6.605 2.915 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.795 0.710 0.965 2.425 ;
        RECT 0.105 2.255 0.965 2.425 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 0.710 2.370 0.880 ;
        RECT 2.200 0.480 2.370 2.665 ;
        RECT 2.200 1.655 2.460 1.955 ;
        RECT 2.200 0.480 3.025 0.650 ;
        RECT 5.505 2.395 5.675 2.665 ;
        RECT 2.200 2.495 5.675 2.665 ;
        RECT 6.225 1.330 6.395 2.565 ;
        RECT 6.225 1.330 6.525 1.500 ;
        RECT 5.505 2.395 7.120 2.565 ;
        RECT 6.950 2.395 7.120 2.795 ;
        RECT 4.465 1.600 5.210 1.770 ;
        RECT 5.040 1.125 5.210 2.280 ;
        RECT 5.875 0.605 6.045 1.295 ;
        RECT 5.015 1.125 6.045 1.295 ;
        RECT 7.090 0.605 7.260 0.945 ;
        RECT 5.875 0.605 7.260 0.775 ;
        RECT 8.265 0.705 8.565 0.945 ;
        RECT 7.090 0.775 8.565 0.945 ;
        RECT 8.015 1.125 8.315 1.495 ;
        RECT 7.255 1.325 8.655 1.495 ;
        RECT 8.485 1.325 8.655 2.280 ;
        RECT 8.485 1.675 8.785 2.280 ;
        RECT 8.485 1.675 9.300 1.845 ;
        RECT 6.515 0.955 6.875 1.125 ;
        RECT 6.705 0.955 6.875 2.215 ;
        RECT 6.620 2.045 6.920 2.215 ;
        RECT 6.705 1.675 8.035 1.845 ;
        RECT 7.865 1.675 8.035 2.630 ;
        RECT 9.830 1.530 10.000 2.630 ;
        RECT 7.865 2.460 10.000 2.630 ;
  END 
END FFDNRHD1XHT

MACRO FFDNHDMXHT
  CLASS  CORE ;
  FOREIGN FFDNHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.610 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.270 1.060 8.510 1.360 ;
        RECT 8.300 1.060 8.510 2.435 ;
        RECT 8.270 1.980 8.510 2.435 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.230 1.060 7.400 1.385 ;
        RECT 7.230 2.000 7.400 2.300 ;
        RECT 7.230 1.205 7.690 1.385 ;
        RECT 7.480 1.205 7.690 2.235 ;
        RECT 7.230 2.000 7.690 2.235 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.625 1.210 1.985 1.740 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.530 ;
        RECT 1.535 -0.300 1.835 0.530 ;
        RECT 3.315 -0.300 3.615 0.630 ;
        RECT 4.295 -0.300 4.595 0.630 ;
        RECT 6.185 -0.300 6.485 0.470 ;
        RECT 7.715 -0.300 8.015 0.595 ;
        RECT 0.000 -0.300 8.610 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.545 0.955 3.990 ;
        RECT 1.500 2.520 1.670 3.990 ;
        RECT 3.435 3.160 3.735 3.990 ;
        RECT 4.295 3.160 4.595 3.990 ;
        RECT 6.195 2.830 6.495 3.990 ;
        RECT 7.715 2.925 8.015 3.990 ;
        RECT 0.000 3.390 8.610 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.550 0.865 2.720 2.280 ;
        RECT 2.550 1.675 3.955 1.845 ;
        RECT 3.930 0.865 4.100 1.470 ;
        RECT 3.175 1.300 4.705 1.470 ;
        RECT 4.535 1.300 4.705 2.215 ;
        RECT 3.865 2.045 4.705 2.215 ;
        RECT 1.145 1.060 1.445 1.230 ;
        RECT 1.275 1.060 1.445 2.245 ;
        RECT 1.145 2.075 2.020 2.245 ;
        RECT 1.850 2.075 2.020 3.075 ;
        RECT 2.855 2.810 3.155 3.075 ;
        RECT 1.850 2.905 3.155 3.075 ;
        RECT 2.855 2.810 5.180 2.980 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.795 0.710 0.965 2.365 ;
        RECT 0.105 2.195 0.965 2.365 ;
        RECT 0.795 1.600 1.095 1.770 ;
        RECT 0.795 0.710 2.370 0.880 ;
        RECT 2.200 0.515 2.370 2.725 ;
        RECT 2.200 2.460 2.575 2.725 ;
        RECT 2.200 0.515 2.995 0.685 ;
        RECT 4.885 0.500 5.055 2.630 ;
        RECT 4.885 0.500 5.285 0.670 ;
        RECT 4.885 2.440 5.755 2.630 ;
        RECT 2.200 2.460 5.755 2.630 ;
        RECT 5.945 1.220 7.050 1.390 ;
        RECT 6.720 0.785 6.890 1.390 ;
        RECT 6.880 1.220 7.050 2.215 ;
        RECT 6.625 2.045 7.050 2.215 ;
        RECT 6.880 1.565 7.275 1.735 ;
        RECT 5.300 0.875 5.470 2.215 ;
        RECT 5.235 2.045 6.445 2.215 ;
        RECT 6.275 1.675 6.445 2.650 ;
        RECT 6.275 1.675 6.700 1.845 ;
        RECT 7.920 1.520 8.090 2.650 ;
        RECT 6.275 2.480 8.090 2.650 ;
        RECT 7.920 1.520 8.110 1.820 ;
  END 
END FFDNHDMXHT

MACRO FFDNHDLXHT
  CLASS  CORE ;
  FOREIGN FFDNHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.610 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.270 1.060 8.510 1.360 ;
        RECT 8.300 1.060 8.510 2.430 ;
        RECT 8.270 1.980 8.510 2.430 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.230 1.060 7.400 1.470 ;
        RECT 7.230 2.000 7.400 2.300 ;
        RECT 7.230 1.290 7.690 1.470 ;
        RECT 7.480 1.290 7.690 2.235 ;
        RECT 7.230 2.000 7.690 2.235 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.625 1.240 1.985 1.770 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.595 ;
        RECT 1.535 -0.300 1.835 0.595 ;
        RECT 3.315 -0.300 3.615 0.670 ;
        RECT 4.320 -0.300 4.620 0.625 ;
        RECT 6.185 -0.300 6.485 0.550 ;
        RECT 7.715 -0.300 8.015 0.745 ;
        RECT 0.000 -0.300 8.610 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.545 0.955 3.990 ;
        RECT 1.500 2.500 1.670 3.990 ;
        RECT 3.435 3.160 3.735 3.990 ;
        RECT 4.295 3.160 4.595 3.990 ;
        RECT 6.195 2.830 6.495 3.990 ;
        RECT 7.715 2.830 8.015 3.990 ;
        RECT 0.000 3.390 8.610 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.550 0.865 2.720 2.280 ;
        RECT 2.550 1.675 3.955 1.845 ;
        RECT 3.960 0.865 4.130 1.470 ;
        RECT 3.175 1.300 4.705 1.470 ;
        RECT 4.535 1.300 4.705 2.215 ;
        RECT 3.865 2.045 4.705 2.215 ;
        RECT 1.145 1.125 1.445 1.295 ;
        RECT 1.275 1.125 1.445 2.225 ;
        RECT 1.145 2.055 2.020 2.225 ;
        RECT 1.850 2.055 2.020 2.995 ;
        RECT 2.625 2.810 2.855 2.995 ;
        RECT 1.850 2.825 2.855 2.995 ;
        RECT 2.625 2.810 5.175 2.980 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.795 0.775 0.965 2.365 ;
        RECT 0.105 2.195 0.965 2.365 ;
        RECT 0.795 1.590 1.095 1.760 ;
        RECT 0.795 0.775 2.370 0.945 ;
        RECT 2.200 0.515 2.370 2.645 ;
        RECT 2.200 2.460 2.525 2.645 ;
        RECT 2.200 0.515 2.995 0.685 ;
        RECT 4.885 0.500 5.055 2.630 ;
        RECT 4.885 0.500 5.285 0.670 ;
        RECT 2.200 2.460 5.755 2.630 ;
        RECT 5.945 1.220 7.050 1.390 ;
        RECT 6.720 0.785 6.890 1.390 ;
        RECT 6.880 1.220 7.050 2.215 ;
        RECT 6.625 2.045 7.050 2.215 ;
        RECT 6.880 1.650 7.275 1.820 ;
        RECT 5.300 0.875 5.470 2.215 ;
        RECT 5.245 2.045 6.445 2.215 ;
        RECT 6.275 1.675 6.445 2.650 ;
        RECT 6.275 1.675 6.700 1.845 ;
        RECT 7.920 1.520 8.090 2.650 ;
        RECT 6.275 2.480 8.090 2.650 ;
        RECT 7.920 1.520 8.110 1.820 ;
  END 
END FFDNHDLXHT

MACRO FFDNHD2XHT
  CLASS  CORE ;
  FOREIGN FFDNHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.250 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.520 2.015 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.390 0.720 9.560 2.960 ;
        RECT 9.390 1.645 9.740 2.015 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.300 0.720 8.520 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.640 1.265 2.080 1.760 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.600 -0.300 0.900 0.595 ;
        RECT 1.630 -0.300 1.930 0.595 ;
        RECT 3.650 -0.300 3.950 1.020 ;
        RECT 4.700 -0.300 5.000 1.055 ;
        RECT 6.475 -0.300 6.645 0.810 ;
        RECT 7.830 -0.300 8.000 1.120 ;
        RECT 8.805 -0.300 9.105 1.055 ;
        RECT 9.845 -0.300 10.145 1.055 ;
        RECT 0.000 -0.300 10.250 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.645 0.925 3.990 ;
        RECT 1.620 2.480 1.790 3.990 ;
        RECT 3.620 3.095 3.920 3.990 ;
        RECT 4.575 3.095 4.875 3.990 ;
        RECT 6.620 2.785 6.790 3.990 ;
        RECT 7.765 2.975 8.065 3.990 ;
        RECT 8.805 2.975 9.105 3.990 ;
        RECT 9.845 2.295 10.145 3.990 ;
        RECT 0.000 3.390 10.250 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.670 0.850 2.970 1.020 ;
        RECT 2.800 0.850 2.970 2.215 ;
        RECT 2.670 2.045 2.970 2.215 ;
        RECT 2.800 1.675 4.190 1.845 ;
        RECT 4.255 0.985 4.425 1.445 ;
        RECT 3.390 1.275 5.120 1.445 ;
        RECT 4.950 1.275 5.120 2.215 ;
        RECT 4.170 2.045 5.120 2.215 ;
        RECT 1.150 1.125 1.460 1.295 ;
        RECT 1.290 1.125 1.460 2.215 ;
        RECT 1.085 2.045 2.140 2.215 ;
        RECT 1.970 2.045 2.140 2.915 ;
        RECT 1.970 2.745 5.685 2.915 ;
        RECT 5.515 2.745 5.685 3.210 ;
        RECT 5.515 3.040 6.200 3.210 ;
        RECT 0.170 2.195 0.340 2.835 ;
        RECT 0.105 1.125 0.880 1.295 ;
        RECT 0.710 0.775 0.880 2.365 ;
        RECT 0.170 2.195 0.880 2.365 ;
        RECT 0.710 1.590 1.110 1.760 ;
        RECT 0.710 0.775 2.490 0.945 ;
        RECT 2.320 0.480 2.490 2.565 ;
        RECT 2.320 1.605 2.555 1.905 ;
        RECT 2.320 0.480 3.240 0.650 ;
        RECT 5.300 0.710 5.470 2.565 ;
        RECT 2.320 2.395 6.135 2.565 ;
        RECT 5.300 0.710 6.240 0.880 ;
        RECT 5.965 2.395 6.135 2.795 ;
        RECT 6.070 0.710 6.240 1.160 ;
        RECT 6.825 0.480 6.995 1.160 ;
        RECT 6.070 0.990 6.995 1.160 ;
        RECT 6.825 0.480 7.650 0.650 ;
        RECT 6.390 1.675 7.415 1.845 ;
        RECT 7.175 1.060 7.345 1.845 ;
        RECT 7.245 1.600 7.415 2.280 ;
        RECT 7.175 1.600 8.120 1.770 ;
        RECT 5.715 1.060 5.885 2.215 ;
        RECT 5.650 2.045 7.065 2.215 ;
        RECT 6.895 2.045 7.065 2.630 ;
        RECT 6.970 2.460 7.270 3.125 ;
        RECT 9.040 1.535 9.210 2.630 ;
        RECT 6.895 2.460 9.210 2.630 ;
  END 
END FFDNHD2XHT

MACRO FFDNHD1XHT
  CLASS  CORE ;
  FOREIGN FFDNHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.610 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.270 0.720 8.510 1.360 ;
        RECT 8.300 0.720 8.510 2.960 ;
        RECT 8.270 1.980 8.510 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.230 0.720 7.400 1.470 ;
        RECT 7.230 2.000 7.400 2.300 ;
        RECT 7.230 1.290 7.690 1.470 ;
        RECT 7.480 1.290 7.690 2.170 ;
        RECT 7.230 2.000 7.690 2.170 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.625 1.140 1.985 1.605 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.595 ;
        RECT 1.535 -0.300 1.835 0.595 ;
        RECT 3.435 -0.300 3.735 0.525 ;
        RECT 4.295 -0.300 4.595 0.565 ;
        RECT 6.185 -0.300 6.485 0.530 ;
        RECT 7.685 -0.300 7.985 1.055 ;
        RECT 0.000 -0.300 8.610 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.685 2.610 0.985 3.990 ;
        RECT 1.435 2.555 1.605 3.990 ;
        RECT 3.435 3.170 3.735 3.990 ;
        RECT 4.295 3.170 4.595 3.990 ;
        RECT 6.195 2.830 6.495 3.990 ;
        RECT 7.685 2.975 7.985 3.990 ;
        RECT 0.000 3.390 8.610 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.550 1.275 2.875 1.445 ;
        RECT 2.550 0.935 2.720 1.445 ;
        RECT 2.705 1.275 2.875 2.290 ;
        RECT 2.485 2.120 2.875 2.290 ;
        RECT 2.705 1.675 3.955 1.845 ;
        RECT 3.930 0.840 4.100 1.445 ;
        RECT 3.175 1.275 4.705 1.445 ;
        RECT 4.535 1.275 4.705 2.215 ;
        RECT 3.865 2.045 4.705 2.215 ;
        RECT 1.230 1.125 1.400 2.215 ;
        RECT 1.145 1.125 1.445 1.295 ;
        RECT 1.145 2.045 1.955 2.215 ;
        RECT 1.785 2.045 1.955 2.990 ;
        RECT 1.785 2.820 5.285 2.990 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.795 0.775 0.965 2.365 ;
        RECT 0.105 2.195 0.965 2.365 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 0.775 2.370 0.945 ;
        RECT 2.135 1.785 2.305 2.640 ;
        RECT 2.200 0.480 2.370 1.940 ;
        RECT 2.200 1.750 2.525 1.940 ;
        RECT 2.200 0.480 2.995 0.650 ;
        RECT 4.885 0.495 5.055 2.640 ;
        RECT 4.885 0.495 5.285 0.665 ;
        RECT 4.885 2.440 5.795 2.640 ;
        RECT 2.135 2.470 5.795 2.640 ;
        RECT 5.495 2.440 5.795 2.705 ;
        RECT 5.945 1.280 7.050 1.450 ;
        RECT 6.720 0.845 6.890 1.450 ;
        RECT 6.880 1.280 7.050 2.215 ;
        RECT 6.625 2.045 7.050 2.215 ;
        RECT 6.880 1.650 7.300 1.820 ;
        RECT 5.300 0.845 5.470 2.215 ;
        RECT 5.235 2.045 5.535 2.215 ;
        RECT 6.275 1.675 6.445 2.650 ;
        RECT 5.300 1.675 6.700 1.845 ;
        RECT 7.920 1.520 8.090 2.650 ;
        RECT 6.275 2.480 8.090 2.650 ;
        RECT 7.920 1.520 8.110 1.820 ;
  END 
END FFDNHD1XHT

MACRO FFDHQHDMXHT
  CLASS  CORE ;
  FOREIGN FFDHQHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.020 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.680 1.060 8.920 2.460 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.420 1.265 2.805 1.800 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 -0.300 0.860 1.060 ;
        RECT 2.380 -0.300 2.550 1.000 ;
        RECT 4.165 -0.300 4.465 0.525 ;
        RECT 5.225 -0.300 5.525 1.095 ;
        RECT 6.950 -0.300 7.120 0.780 ;
        RECT 8.160 -0.300 8.330 1.210 ;
        RECT 0.000 -0.300 9.020 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.850 1.525 1.340 1.950 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.385 2.895 1.685 3.990 ;
        RECT 2.320 2.760 2.490 3.990 ;
        RECT 4.255 3.160 4.555 3.990 ;
        RECT 5.225 3.160 5.525 3.990 ;
        RECT 7.005 2.795 7.305 3.990 ;
        RECT 8.065 2.745 8.365 3.990 ;
        RECT 0.000 3.390 9.020 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.175 1.125 1.785 1.295 ;
        RECT 1.615 1.125 1.785 2.300 ;
        RECT 0.925 2.130 1.785 2.300 ;
        RECT 1.615 1.525 1.830 1.825 ;
        RECT 3.370 0.865 3.540 2.280 ;
        RECT 3.370 1.675 4.775 1.845 ;
        RECT 4.780 0.840 4.950 1.445 ;
        RECT 3.995 1.275 5.635 1.445 ;
        RECT 5.465 1.275 5.635 2.215 ;
        RECT 4.715 2.045 5.635 2.215 ;
        RECT 0.170 1.060 0.340 1.980 ;
        RECT 0.170 1.810 0.610 1.980 ;
        RECT 0.440 1.810 0.610 2.715 ;
        RECT 1.965 2.395 2.140 2.715 ;
        RECT 0.440 2.545 2.140 2.715 ;
        RECT 1.965 2.395 2.840 2.565 ;
        RECT 2.670 2.395 2.840 3.190 ;
        RECT 3.675 2.835 3.910 3.190 ;
        RECT 2.670 3.020 3.910 3.190 ;
        RECT 3.860 2.810 4.030 3.005 ;
        RECT 3.675 2.835 4.030 3.005 ;
        RECT 3.860 2.810 6.215 2.980 ;
        RECT 6.875 1.495 7.855 1.665 ;
        RECT 7.650 1.060 7.820 1.665 ;
        RECT 7.685 1.495 7.855 2.215 ;
        RECT 7.555 2.045 7.855 2.215 ;
        RECT 1.725 0.765 2.180 0.935 ;
        RECT 2.010 0.765 2.180 2.215 ;
        RECT 1.965 2.045 3.190 2.215 ;
        RECT 3.020 0.515 3.190 2.840 ;
        RECT 3.020 2.460 3.395 2.840 ;
        RECT 3.020 0.515 3.815 0.685 ;
        RECT 5.815 1.425 5.985 2.630 ;
        RECT 5.880 0.710 6.050 1.595 ;
        RECT 5.815 1.425 6.050 1.595 ;
        RECT 5.815 2.440 6.595 2.630 ;
        RECT 6.425 2.440 6.595 2.755 ;
        RECT 3.020 2.460 6.595 2.630 ;
        RECT 5.880 0.710 6.770 0.880 ;
        RECT 6.425 2.585 6.725 2.755 ;
        RECT 6.600 0.710 6.770 1.150 ;
        RECT 7.300 0.480 7.470 1.150 ;
        RECT 6.600 0.980 7.470 1.150 ;
        RECT 7.300 0.480 7.910 0.650 ;
        RECT 6.250 1.060 6.420 2.215 ;
        RECT 6.175 2.045 7.375 2.215 ;
        RECT 7.205 2.045 7.375 2.565 ;
        RECT 7.485 2.395 7.655 2.900 ;
        RECT 8.330 1.520 8.500 2.565 ;
        RECT 7.205 2.395 8.500 2.565 ;
  END 
END FFDHQHDMXHT

MACRO FFDHQHD3XHT
  CLASS  CORE ;
  FOREIGN FFDHQHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.120 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.630 0.720 11.800 1.405 ;
        RECT 11.630 1.980 11.800 2.960 ;
        RECT 11.630 1.235 12.840 1.405 ;
        RECT 11.630 2.150 12.840 2.360 ;
        RECT 12.670 0.720 12.840 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.280 1.110 3.620 1.800 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.600 -0.300 0.770 0.700 ;
        RECT 2.145 -0.300 2.445 0.745 ;
        RECT 3.170 -0.300 3.470 0.785 ;
        RECT 5.180 -0.300 5.480 0.595 ;
        RECT 6.240 -0.300 6.540 0.595 ;
        RECT 8.080 -0.300 8.380 1.035 ;
        RECT 9.940 -0.300 10.240 0.715 ;
        RECT 11.110 -0.300 11.280 1.120 ;
        RECT 12.085 -0.300 12.385 1.055 ;
        RECT 0.000 -0.300 13.120 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 1.500 1.525 2.015 1.950 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.605 2.935 0.905 3.990 ;
        RECT 1.995 2.935 2.295 3.990 ;
        RECT 3.160 2.790 3.330 3.990 ;
        RECT 5.160 3.095 5.460 3.990 ;
        RECT 6.240 3.095 6.540 3.990 ;
        RECT 8.080 2.745 8.380 3.990 ;
        RECT 9.975 2.805 10.145 3.990 ;
        RECT 11.045 2.975 11.345 3.990 ;
        RECT 12.085 2.635 12.385 3.990 ;
        RECT 0.000 3.390 13.120 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.595 1.125 2.365 1.295 ;
        RECT 2.195 1.125 2.365 2.300 ;
        RECT 1.455 2.130 2.365 2.300 ;
        RECT 2.195 1.525 2.575 1.825 ;
        RECT 4.210 0.850 4.510 1.020 ;
        RECT 4.340 0.850 4.510 2.215 ;
        RECT 4.210 2.045 4.510 2.215 ;
        RECT 4.340 1.675 5.710 1.845 ;
        RECT 0.970 1.125 1.140 2.650 ;
        RECT 1.150 0.720 1.320 1.295 ;
        RECT 0.105 1.125 1.385 1.295 ;
        RECT 2.780 2.395 2.960 2.650 ;
        RECT 0.970 2.480 2.960 2.650 ;
        RECT 2.780 2.395 3.680 2.565 ;
        RECT 3.510 2.395 3.680 2.915 ;
        RECT 3.510 2.745 7.165 2.915 ;
        RECT 6.980 2.745 7.165 3.195 ;
        RECT 6.980 3.025 7.620 3.195 ;
        RECT 4.930 1.275 6.060 1.445 ;
        RECT 5.730 1.125 6.030 1.445 ;
        RECT 5.890 1.275 6.060 2.215 ;
        RECT 5.710 2.045 6.060 2.215 ;
        RECT 5.890 1.585 8.555 1.755 ;
        RECT 2.755 1.060 2.925 2.215 ;
        RECT 2.545 2.045 4.030 2.215 ;
        RECT 3.860 0.480 4.030 2.565 ;
        RECT 3.860 1.595 4.095 1.895 ;
        RECT 3.860 0.480 4.860 0.650 ;
        RECT 4.690 0.480 4.860 0.945 ;
        RECT 6.730 0.480 6.900 0.945 ;
        RECT 4.690 0.775 6.900 0.945 ;
        RECT 6.730 0.480 7.620 0.650 ;
        RECT 3.860 2.395 9.570 2.565 ;
        RECT 9.400 2.395 9.570 3.005 ;
        RECT 9.770 1.590 10.725 1.760 ;
        RECT 10.555 1.060 10.725 2.280 ;
        RECT 7.225 1.060 7.395 1.405 ;
        RECT 7.225 1.235 9.235 1.405 ;
        RECT 9.065 1.060 9.235 2.215 ;
        RECT 7.160 2.045 10.375 2.215 ;
        RECT 10.205 2.045 10.375 2.630 ;
        RECT 10.375 2.460 10.545 2.820 ;
        RECT 11.195 1.590 11.365 2.630 ;
        RECT 10.205 2.460 11.365 2.630 ;
        RECT 11.195 1.590 12.465 1.760 ;
  END 
END FFDHQHD3XHT

MACRO FFDHQHD2XHT
  CLASS  CORE ;
  FOREIGN FFDHQHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.070 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.210 0.720 10.380 2.960 ;
        RECT 10.210 1.655 10.560 2.025 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.870 1.265 3.210 1.800 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.170 -0.300 0.340 1.205 ;
        RECT 1.725 -0.300 2.025 0.745 ;
        RECT 2.760 -0.300 3.060 0.785 ;
        RECT 4.770 -0.300 5.070 0.595 ;
        RECT 6.750 -0.300 7.050 1.015 ;
        RECT 8.675 -0.300 8.845 0.780 ;
        RECT 9.690 -0.300 9.860 0.780 ;
        RECT 10.665 -0.300 10.965 1.055 ;
        RECT 0.000 -0.300 11.070 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 1.180 1.525 1.655 1.950 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.935 0.925 3.990 ;
        RECT 1.645 2.830 1.945 3.990 ;
        RECT 2.750 2.790 2.920 3.990 ;
        RECT 4.750 3.095 5.050 3.990 ;
        RECT 6.750 2.800 7.050 3.990 ;
        RECT 8.675 2.830 8.845 3.990 ;
        RECT 9.625 2.975 9.925 3.990 ;
        RECT 10.665 2.295 10.965 3.990 ;
        RECT 0.000 3.390 11.070 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.175 1.125 2.010 1.295 ;
        RECT 1.840 1.125 2.010 2.300 ;
        RECT 1.175 2.130 2.010 2.300 ;
        RECT 1.840 1.525 2.165 1.825 ;
        RECT 3.800 0.850 4.100 1.020 ;
        RECT 3.930 0.850 4.100 2.215 ;
        RECT 3.800 2.045 4.100 2.215 ;
        RECT 3.930 1.675 5.300 1.845 ;
        RECT 0.690 0.720 0.860 2.650 ;
        RECT 2.370 2.395 2.550 2.650 ;
        RECT 0.690 2.480 2.550 2.650 ;
        RECT 2.370 2.395 3.270 2.565 ;
        RECT 3.100 2.395 3.270 2.915 ;
        RECT 5.190 2.745 5.360 2.930 ;
        RECT 3.100 2.745 5.360 2.915 ;
        RECT 5.190 2.760 6.310 2.930 ;
        RECT 6.010 2.760 6.310 3.210 ;
        RECT 4.520 1.275 5.650 1.445 ;
        RECT 5.320 1.125 5.620 1.445 ;
        RECT 5.480 1.275 5.650 2.215 ;
        RECT 5.300 2.045 5.650 2.215 ;
        RECT 5.480 1.585 7.225 1.755 ;
        RECT 2.345 1.060 2.515 2.215 ;
        RECT 2.215 2.045 3.620 2.215 ;
        RECT 3.450 0.480 3.620 2.565 ;
        RECT 3.450 1.605 3.685 1.905 ;
        RECT 3.450 0.480 4.450 0.650 ;
        RECT 4.280 0.480 4.450 0.945 ;
        RECT 5.525 0.480 5.695 0.945 ;
        RECT 4.280 0.775 5.695 0.945 ;
        RECT 5.540 2.395 5.710 2.580 ;
        RECT 3.450 2.395 5.710 2.565 ;
        RECT 5.525 0.480 6.310 0.650 ;
        RECT 5.540 2.410 8.185 2.580 ;
        RECT 8.015 2.410 8.185 2.795 ;
        RECT 8.440 1.590 9.395 1.760 ;
        RECT 9.225 1.060 9.395 2.280 ;
        RECT 5.895 1.060 6.065 1.405 ;
        RECT 5.895 1.235 7.935 1.405 ;
        RECT 7.765 1.060 7.935 2.230 ;
        RECT 5.830 2.060 9.045 2.230 ;
        RECT 8.875 2.060 9.045 2.630 ;
        RECT 9.045 2.460 9.215 2.820 ;
        RECT 9.860 1.525 10.030 2.630 ;
        RECT 8.875 2.460 10.030 2.630 ;
  END 
END FFDHQHD2XHT

MACRO FFDHQHD1XHT
  CLASS  CORE ;
  FOREIGN FFDHQHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.020 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.680 0.720 8.920 2.960 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.420 1.265 2.805 1.795 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 -0.300 0.860 1.060 ;
        RECT 2.380 -0.300 2.550 1.000 ;
        RECT 4.165 -0.300 4.465 0.525 ;
        RECT 5.225 -0.300 5.525 0.945 ;
        RECT 6.950 -0.300 7.120 0.780 ;
        RECT 8.160 -0.300 8.330 1.120 ;
        RECT 0.000 -0.300 9.020 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.850 1.525 1.340 1.950 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.385 2.895 1.685 3.990 ;
        RECT 2.320 2.760 2.490 3.990 ;
        RECT 4.255 3.160 4.555 3.990 ;
        RECT 5.225 3.160 5.525 3.990 ;
        RECT 7.005 2.795 7.305 3.990 ;
        RECT 8.095 2.975 8.395 3.990 ;
        RECT 0.000 3.390 9.020 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.175 1.125 1.785 1.295 ;
        RECT 1.615 1.125 1.785 2.300 ;
        RECT 0.925 2.130 1.785 2.300 ;
        RECT 1.615 1.525 1.830 1.825 ;
        RECT 3.370 0.865 3.540 2.280 ;
        RECT 3.370 1.675 4.775 1.845 ;
        RECT 4.780 0.840 4.950 1.445 ;
        RECT 3.995 1.275 5.635 1.445 ;
        RECT 5.465 1.275 5.635 2.215 ;
        RECT 4.715 2.045 5.635 2.215 ;
        RECT 0.170 1.060 0.340 1.980 ;
        RECT 0.170 1.810 0.610 1.980 ;
        RECT 0.440 1.810 0.610 2.715 ;
        RECT 1.965 2.395 2.140 2.715 ;
        RECT 0.440 2.545 2.140 2.715 ;
        RECT 1.965 2.395 2.840 2.565 ;
        RECT 2.670 2.395 2.840 3.170 ;
        RECT 3.675 2.835 3.910 3.170 ;
        RECT 3.675 2.835 4.030 3.005 ;
        RECT 2.670 3.000 3.910 3.170 ;
        RECT 3.860 2.810 4.030 3.005 ;
        RECT 3.860 2.810 6.085 2.980 ;
        RECT 5.915 2.810 6.085 3.195 ;
        RECT 5.915 3.025 6.215 3.195 ;
        RECT 6.875 1.495 7.855 1.665 ;
        RECT 7.650 1.060 7.820 1.665 ;
        RECT 7.685 1.495 7.855 2.215 ;
        RECT 7.555 2.045 7.855 2.215 ;
        RECT 1.725 0.765 2.180 0.935 ;
        RECT 2.010 0.765 2.180 2.215 ;
        RECT 1.965 2.045 3.190 2.215 ;
        RECT 3.020 0.515 3.190 2.820 ;
        RECT 3.020 2.460 3.395 2.820 ;
        RECT 3.020 0.515 3.815 0.685 ;
        RECT 5.815 0.710 5.985 2.630 ;
        RECT 5.815 2.440 6.595 2.630 ;
        RECT 5.815 0.710 6.760 0.880 ;
        RECT 6.425 2.440 6.595 2.755 ;
        RECT 3.020 2.460 6.595 2.630 ;
        RECT 6.425 2.585 6.725 2.755 ;
        RECT 6.590 0.710 6.760 1.150 ;
        RECT 7.300 0.480 7.470 1.150 ;
        RECT 6.590 0.980 7.470 1.150 ;
        RECT 7.300 0.480 7.910 0.650 ;
        RECT 6.230 1.060 6.400 2.215 ;
        RECT 6.165 2.045 7.375 2.215 ;
        RECT 7.205 2.045 7.375 2.565 ;
        RECT 7.485 2.395 7.655 2.900 ;
        RECT 8.330 1.520 8.500 2.565 ;
        RECT 7.205 2.395 8.500 2.565 ;
  END 
END FFDHQHD1XHT

MACRO FFDHDMXHT
  CLASS  CORE ;
  FOREIGN FFDHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.610 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.270 1.060 8.510 1.360 ;
        RECT 8.300 1.060 8.510 2.435 ;
        RECT 8.270 1.980 8.510 2.435 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.230 1.060 7.400 1.410 ;
        RECT 7.230 2.000 7.400 2.300 ;
        RECT 7.230 1.230 7.690 1.410 ;
        RECT 7.480 1.230 7.690 2.170 ;
        RECT 7.230 2.000 7.690 2.170 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.600 1.265 1.985 1.755 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.585 -0.300 0.885 0.745 ;
        RECT 1.535 -0.300 1.835 0.785 ;
        RECT 3.315 -0.300 3.615 0.605 ;
        RECT 4.295 -0.300 4.595 0.565 ;
        RECT 6.185 -0.300 6.485 0.470 ;
        RECT 7.715 -0.300 8.015 0.595 ;
        RECT 0.000 -0.300 8.610 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 2.745 0.865 3.990 ;
        RECT 1.500 2.760 1.670 3.990 ;
        RECT 3.435 3.160 3.735 3.990 ;
        RECT 4.295 3.160 4.595 3.990 ;
        RECT 6.195 2.830 6.495 3.990 ;
        RECT 7.685 2.925 7.985 3.990 ;
        RECT 0.000 3.390 8.610 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.550 0.865 2.720 2.280 ;
        RECT 2.550 1.675 3.955 1.845 ;
        RECT 3.930 0.840 4.100 1.445 ;
        RECT 3.175 1.275 4.705 1.445 ;
        RECT 4.535 1.275 4.705 2.215 ;
        RECT 3.865 2.045 4.705 2.215 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.195 0.965 2.365 ;
        RECT 0.795 1.125 0.965 2.565 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 2.395 2.020 2.565 ;
        RECT 1.850 2.395 2.020 3.075 ;
        RECT 2.855 2.810 3.155 3.075 ;
        RECT 1.850 2.905 3.155 3.075 ;
        RECT 2.855 2.810 5.175 2.980 ;
        RECT 1.210 1.060 1.400 1.360 ;
        RECT 1.230 1.060 1.400 2.215 ;
        RECT 1.145 2.045 2.370 2.215 ;
        RECT 2.200 0.515 2.370 2.725 ;
        RECT 2.200 2.460 2.575 2.725 ;
        RECT 2.200 0.515 2.995 0.685 ;
        RECT 4.885 0.525 5.055 2.630 ;
        RECT 4.885 0.525 5.285 0.695 ;
        RECT 4.885 2.440 5.755 2.630 ;
        RECT 2.200 2.460 5.755 2.630 ;
        RECT 5.945 1.220 7.050 1.390 ;
        RECT 6.720 0.785 6.890 1.390 ;
        RECT 6.880 1.220 7.050 2.215 ;
        RECT 6.625 2.045 7.050 2.215 ;
        RECT 6.880 1.590 7.300 1.760 ;
        RECT 5.300 0.875 5.470 2.215 ;
        RECT 5.235 2.045 5.535 2.215 ;
        RECT 6.275 1.675 6.445 2.650 ;
        RECT 5.300 1.675 6.700 1.845 ;
        RECT 7.920 1.520 8.090 2.650 ;
        RECT 6.275 2.480 8.090 2.650 ;
        RECT 7.920 1.520 8.110 1.820 ;
  END 
END FFDHDMXHT

MACRO FFDHD1XHT
  CLASS  CORE ;
  FOREIGN FFDHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.610 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.270 0.720 8.510 1.360 ;
        RECT 8.300 0.720 8.510 2.960 ;
        RECT 8.270 1.980 8.510 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 7.230 0.720 7.400 1.470 ;
        RECT 7.230 2.000 7.400 2.300 ;
        RECT 7.230 1.290 7.690 1.470 ;
        RECT 7.480 1.290 7.690 2.235 ;
        RECT 7.230 2.000 7.690 2.235 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.600 1.265 1.985 1.670 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 -0.300 0.895 0.745 ;
        RECT 1.535 -0.300 1.835 0.720 ;
        RECT 3.315 -0.300 3.615 0.525 ;
        RECT 4.295 -0.300 4.595 0.565 ;
        RECT 6.185 -0.300 6.485 0.470 ;
        RECT 7.685 -0.300 7.985 1.055 ;
        RECT 0.000 -0.300 8.610 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 2.745 0.865 3.990 ;
        RECT 1.500 2.760 1.670 3.990 ;
        RECT 3.435 3.160 3.735 3.990 ;
        RECT 4.295 3.160 4.595 3.990 ;
        RECT 6.195 2.830 6.495 3.990 ;
        RECT 7.685 2.975 7.985 3.990 ;
        RECT 0.000 3.390 8.610 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.550 0.840 2.720 2.280 ;
        RECT 2.550 1.675 3.955 1.845 ;
        RECT 3.930 0.840 4.100 1.445 ;
        RECT 3.175 1.275 4.705 1.445 ;
        RECT 4.535 1.275 4.705 2.215 ;
        RECT 3.865 2.045 4.705 2.215 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.195 0.965 2.365 ;
        RECT 0.795 1.125 0.965 2.565 ;
        RECT 0.795 1.525 1.040 1.825 ;
        RECT 0.795 2.395 2.020 2.565 ;
        RECT 1.850 2.395 2.020 3.170 ;
        RECT 2.855 2.810 3.090 3.170 ;
        RECT 1.850 3.000 3.090 3.170 ;
        RECT 2.855 2.810 3.155 3.005 ;
        RECT 2.855 2.810 5.285 2.980 ;
        RECT 1.210 0.995 1.400 1.295 ;
        RECT 1.230 0.995 1.400 2.215 ;
        RECT 1.145 2.045 2.370 2.215 ;
        RECT 2.200 0.490 2.370 2.820 ;
        RECT 2.200 2.460 2.525 2.820 ;
        RECT 2.200 0.490 2.995 0.660 ;
        RECT 4.885 1.425 5.055 2.630 ;
        RECT 4.950 0.500 5.120 1.595 ;
        RECT 4.885 1.425 5.120 1.595 ;
        RECT 4.950 0.500 5.285 0.670 ;
        RECT 4.885 2.440 5.730 2.630 ;
        RECT 2.200 2.460 5.730 2.630 ;
        RECT 5.560 2.440 5.730 2.770 ;
        RECT 5.945 1.220 7.050 1.390 ;
        RECT 6.720 0.785 6.890 1.390 ;
        RECT 6.880 1.220 7.050 2.215 ;
        RECT 6.625 2.045 7.050 2.215 ;
        RECT 6.880 1.650 7.275 1.820 ;
        RECT 5.300 0.875 5.470 2.215 ;
        RECT 5.235 2.045 6.445 2.215 ;
        RECT 6.275 1.675 6.445 2.650 ;
        RECT 6.275 1.675 6.700 1.845 ;
        RECT 7.920 1.520 8.090 2.650 ;
        RECT 6.275 2.480 8.090 2.650 ;
        RECT 7.920 1.520 8.110 1.820 ;
  END 
END FFDHD1XHT

MACRO FFDHD1XSPGHT
  CLASS  CORE ;
  FOREIGN FFDHD1XSPGHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.610 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 7.725 0.300 8.265 3.080 ;
      LAYER V7 ;
        RECT 7.815 0.435 8.175 0.795 ;
      LAYER M7 ;
        RECT 7.685 0.415 8.455 0.815 ;
      LAYER V6 ;
        RECT 7.900 0.520 8.090 0.710 ;
      LAYER M4 ;
        RECT 7.895 0.315 8.095 2.430 ;
      LAYER V3 ;
        RECT 7.900 1.750 8.090 1.940 ;
      LAYER M3 ;
        RECT 7.805 1.645 8.505 2.045 ;
      LAYER V2 ;
        RECT 8.310 1.750 8.500 1.940 ;
      LAYER M2 ;
        RECT 8.305 1.175 8.505 2.160 ;
      LAYER V1 ;
        RECT 8.310 1.750 8.500 1.940 ;
      LAYER M1 ;
        RECT 8.270 0.720 8.510 1.360 ;
        RECT 8.300 0.720 8.510 2.960 ;
        RECT 8.270 1.980 8.510 2.960 ;
      LAYER M6 ;
        RECT 7.895 0.300 8.095 2.090 ;
      LAYER V5 ;
        RECT 7.900 0.520 8.090 0.710 ;
      LAYER M5 ;
        RECT 7.685 0.515 8.455 0.715 ;
      LAYER V4 ;
        RECT 7.900 0.520 8.090 0.710 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 6.495 0.300 7.035 3.080 ;
      LAYER V7 ;
        RECT 6.585 0.435 6.945 0.795 ;
      LAYER M7 ;
        RECT 5.840 0.415 7.445 0.815 ;
      LAYER V6 ;
        RECT 6.670 0.520 6.860 0.710 ;
      LAYER M4 ;
        RECT 7.075 0.335 7.275 2.160 ;
      LAYER V3 ;
        RECT 7.080 0.930 7.270 1.120 ;
      LAYER M3 ;
        RECT 6.945 0.925 7.790 1.125 ;
      LAYER V2 ;
        RECT 7.490 0.930 7.680 1.120 ;
      LAYER M2 ;
        RECT 7.485 0.765 7.685 2.280 ;
      LAYER V1 ;
        RECT 7.490 1.750 7.680 1.940 ;
      LAYER M1 ;
        RECT 7.230 0.720 7.400 1.470 ;
        RECT 7.230 2.000 7.400 2.300 ;
        RECT 7.230 1.290 7.690 1.470 ;
        RECT 7.480 1.290 7.690 2.235 ;
        RECT 7.230 2.000 7.690 2.235 ;
      LAYER M6 ;
        RECT 6.665 0.300 6.865 2.090 ;
      LAYER V5 ;
        RECT 6.670 0.520 6.860 0.710 ;
      LAYER M5 ;
        RECT 5.840 0.515 7.445 0.715 ;
      LAYER V4 ;
        RECT 7.080 0.520 7.270 0.710 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 1.985 0.300 2.525 3.065 ;
      LAYER V7 ;
        RECT 2.075 0.435 2.435 0.795 ;
      LAYER M7 ;
        RECT 1.845 0.415 2.855 0.815 ;
      LAYER V6 ;
        RECT 2.160 0.520 2.350 0.710 ;
      LAYER M4 ;
        RECT 2.155 0.300 2.355 2.610 ;
      LAYER V3 ;
        RECT 2.160 2.160 2.350 2.350 ;
      LAYER M3 ;
        RECT 1.655 2.155 2.665 2.355 ;
      LAYER V2 ;
        RECT 1.750 2.160 1.940 2.350 ;
      LAYER M2 ;
        RECT 1.745 1.200 1.945 2.505 ;
      LAYER V1 ;
        RECT 1.750 1.340 1.940 1.530 ;
      LAYER M1 ;
        RECT 1.600 1.265 1.985 1.670 ;
      LAYER M6 ;
        RECT 2.155 0.300 2.355 2.090 ;
      LAYER V5 ;
        RECT 2.160 0.520 2.350 0.710 ;
      LAYER M5 ;
        RECT 1.845 0.515 2.855 0.715 ;
      LAYER V4 ;
        RECT 2.160 0.520 2.350 0.710 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.745 ;
        RECT 1.535 -0.300 1.835 0.720 ;
        RECT 3.315 -0.300 3.615 0.525 ;
        RECT 4.295 -0.300 4.595 0.565 ;
        RECT 6.185 -0.300 6.485 0.470 ;
        RECT 7.685 -0.300 7.985 1.055 ;
        RECT 0.000 -0.300 8.610 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M8 ;
        RECT 0.755 0.300 1.295 3.065 ;
      LAYER V7 ;
        RECT 0.845 0.435 1.205 0.795 ;
      LAYER M7 ;
        RECT 0.335 0.415 1.295 0.815 ;
      LAYER V6 ;
        RECT 0.930 0.520 1.120 0.710 ;
      LAYER M4 ;
        RECT 0.515 0.355 0.715 1.820 ;
      LAYER V3 ;
        RECT 0.520 1.340 0.710 1.530 ;
      LAYER M3 ;
        RECT 0.105 1.265 0.820 1.605 ;
      LAYER V2 ;
        RECT 0.110 1.340 0.300 1.530 ;
      LAYER M2 ;
        RECT 0.105 1.165 0.305 2.050 ;
      LAYER V1 ;
        RECT 0.110 1.750 0.300 1.940 ;
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
      LAYER M6 ;
        RECT 0.925 0.300 1.125 2.090 ;
      LAYER V5 ;
        RECT 0.930 0.520 1.120 0.710 ;
      LAYER M5 ;
        RECT 0.335 0.515 1.295 0.715 ;
      LAYER V4 ;
        RECT 0.520 0.520 0.710 0.710 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 2.810 0.865 3.990 ;
        RECT 1.500 2.760 1.670 3.990 ;
        RECT 3.435 3.160 3.735 3.990 ;
        RECT 4.295 3.160 4.595 3.990 ;
        RECT 6.195 2.830 6.495 3.990 ;
        RECT 7.685 2.975 7.985 3.990 ;
        RECT 0.000 3.390 8.610 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 2.550 0.865 2.720 2.280 ;
        RECT 2.550 1.675 3.955 1.845 ;
        RECT 3.930 0.840 4.100 1.445 ;
        RECT 3.175 1.275 4.705 1.445 ;
        RECT 4.535 1.275 4.705 2.215 ;
        RECT 3.865 2.045 4.705 2.215 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.195 0.965 2.365 ;
        RECT 0.795 1.125 0.965 2.565 ;
        RECT 0.795 1.525 1.030 1.825 ;
        RECT 0.795 2.395 2.020 2.565 ;
        RECT 1.850 2.395 2.020 3.170 ;
        RECT 2.855 2.810 3.090 3.170 ;
        RECT 1.850 3.000 3.090 3.170 ;
        RECT 2.855 2.810 3.155 3.005 ;
        RECT 2.855 2.810 5.285 2.980 ;
        RECT 1.210 0.995 1.400 1.295 ;
        RECT 1.230 0.995 1.400 2.215 ;
        RECT 1.145 2.045 2.370 2.215 ;
        RECT 2.200 0.515 2.370 2.820 ;
        RECT 2.200 2.460 2.575 2.820 ;
        RECT 2.200 0.515 2.995 0.685 ;
        RECT 4.885 1.425 5.055 2.630 ;
        RECT 4.950 0.500 5.120 1.595 ;
        RECT 4.885 1.425 5.120 1.595 ;
        RECT 4.950 0.500 5.285 0.670 ;
        RECT 4.885 2.440 5.665 2.630 ;
        RECT 5.495 2.440 5.665 2.705 ;
        RECT 2.200 2.460 5.665 2.630 ;
        RECT 5.495 2.535 5.795 2.705 ;
        RECT 6.655 0.850 7.050 1.020 ;
        RECT 5.945 1.220 7.050 1.390 ;
        RECT 6.880 0.850 7.050 2.215 ;
        RECT 6.625 2.045 7.050 2.215 ;
        RECT 6.880 1.650 7.275 1.820 ;
        RECT 5.300 0.875 5.470 2.215 ;
        RECT 5.235 2.045 5.535 2.215 ;
        RECT 6.275 1.675 6.445 2.650 ;
        RECT 5.300 1.675 6.700 1.845 ;
        RECT 7.920 1.520 8.090 2.650 ;
        RECT 6.275 2.480 8.090 2.650 ;
        RECT 7.920 1.520 8.110 1.820 ;
  END 
END FFDHD1XSPGHT

MACRO FFDCRHDMXHT
  CLASS  CORE ;
  FOREIGN FFDCRHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.430 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.090 1.060 9.330 2.280 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.080 1.060 8.510 1.360 ;
        RECT 8.300 1.060 8.510 2.280 ;
        RECT 8.080 1.980 8.510 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.680 1.265 2.080 1.780 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.380 1.265 2.770 1.780 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.670 -0.300 0.970 0.845 ;
        RECT 1.835 -0.300 2.135 0.735 ;
        RECT 4.215 -0.300 4.515 1.020 ;
        RECT 5.370 -0.300 5.540 0.730 ;
        RECT 7.150 -0.300 7.320 0.850 ;
        RECT 8.640 -0.300 8.810 0.660 ;
        RECT 0.000 -0.300 9.430 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 2.810 0.865 3.990 ;
        RECT 2.085 2.810 2.385 3.990 ;
        RECT 4.215 3.160 4.515 3.990 ;
        RECT 5.185 3.160 5.485 3.990 ;
        RECT 6.895 2.540 7.065 3.990 ;
        RECT 8.540 2.860 8.710 3.990 ;
        RECT 0.000 3.390 9.430 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.690 1.980 2.900 2.280 ;
        RECT 3.330 0.900 3.600 1.200 ;
        RECT 3.430 0.900 3.600 2.280 ;
        RECT 3.430 1.675 4.700 1.845 ;
        RECT 3.985 1.220 5.095 1.390 ;
        RECT 4.860 0.785 5.030 1.390 ;
        RECT 4.925 1.220 5.095 2.215 ;
        RECT 4.795 2.045 5.095 2.215 ;
        RECT 4.925 1.410 5.670 1.580 ;
        RECT 0.105 1.125 0.935 1.295 ;
        RECT 0.105 2.195 0.935 2.365 ;
        RECT 0.765 1.125 0.935 2.630 ;
        RECT 0.765 1.525 1.130 1.825 ;
        RECT 0.765 2.460 2.860 2.630 ;
        RECT 2.690 2.460 2.860 2.995 ;
        RECT 3.630 2.810 3.930 2.995 ;
        RECT 2.690 2.825 3.930 2.995 ;
        RECT 3.630 2.810 6.065 2.980 ;
        RECT 2.980 1.415 3.250 1.585 ;
        RECT 1.300 0.915 1.500 1.360 ;
        RECT 1.330 0.915 1.500 2.215 ;
        RECT 1.115 2.045 1.500 2.215 ;
        RECT 1.300 0.915 3.150 1.085 ;
        RECT 2.980 0.550 3.150 1.585 ;
        RECT 3.080 1.415 3.250 2.645 ;
        RECT 3.080 2.460 3.380 2.645 ;
        RECT 2.980 0.550 3.775 0.720 ;
        RECT 5.850 0.550 6.020 2.630 ;
        RECT 5.850 0.550 6.180 0.720 ;
        RECT 3.080 2.460 6.580 2.630 ;
        RECT 6.410 2.460 6.580 2.770 ;
        RECT 6.875 1.195 7.900 1.365 ;
        RECT 7.670 0.550 7.840 1.365 ;
        RECT 7.730 1.195 7.900 2.775 ;
        RECT 7.595 2.605 7.900 2.775 ;
        RECT 7.730 1.630 8.120 1.800 ;
        RECT 6.200 0.900 6.370 2.280 ;
        RECT 7.245 1.675 7.415 3.125 ;
        RECT 6.200 1.675 7.550 1.845 ;
        RECT 8.080 2.460 8.250 3.125 ;
        RECT 7.245 2.955 8.250 3.125 ;
        RECT 8.740 1.605 8.910 2.630 ;
        RECT 8.080 2.460 8.910 2.630 ;
  END 
END FFDCRHDMXHT

MACRO FFDCRHDLXHT
  CLASS  CORE ;
  FOREIGN FFDCRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.430 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.090 1.060 9.330 2.445 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.080 1.060 8.510 1.360 ;
        RECT 8.300 1.060 8.510 2.280 ;
        RECT 8.080 1.980 8.510 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.680 1.265 2.070 1.780 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.380 1.265 2.770 1.780 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.685 -0.300 0.985 0.945 ;
        RECT 1.835 -0.300 2.135 0.735 ;
        RECT 4.215 -0.300 4.515 0.970 ;
        RECT 5.305 -0.300 5.605 0.585 ;
        RECT 7.085 -0.300 7.385 0.785 ;
        RECT 8.575 -0.300 8.875 0.745 ;
        RECT 0.000 -0.300 9.430 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.445 2.640 0.615 3.990 ;
        RECT 2.205 2.810 2.505 3.990 ;
        RECT 4.215 3.160 4.515 3.990 ;
        RECT 5.185 3.160 5.485 3.990 ;
        RECT 6.895 2.540 7.065 3.990 ;
        RECT 8.475 2.810 8.775 3.990 ;
        RECT 0.000 3.390 9.430 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.690 1.980 2.900 2.280 ;
        RECT 3.330 1.030 3.600 1.200 ;
        RECT 3.330 0.900 3.500 1.200 ;
        RECT 3.430 1.030 3.600 2.280 ;
        RECT 3.430 1.675 4.725 1.845 ;
        RECT 3.985 1.220 5.095 1.390 ;
        RECT 4.860 0.735 5.030 1.390 ;
        RECT 4.925 1.220 5.095 2.215 ;
        RECT 4.795 2.045 5.095 2.215 ;
        RECT 4.925 1.410 5.670 1.580 ;
        RECT 0.105 1.125 0.965 1.295 ;
        RECT 0.105 2.195 0.965 2.365 ;
        RECT 0.795 1.125 0.965 2.985 ;
        RECT 0.795 1.525 1.130 1.825 ;
        RECT 1.810 2.460 1.980 2.985 ;
        RECT 0.795 2.815 1.980 2.985 ;
        RECT 1.810 2.460 2.860 2.630 ;
        RECT 2.690 2.460 2.860 2.980 ;
        RECT 2.690 2.810 6.065 2.980 ;
        RECT 2.980 1.415 3.250 1.585 ;
        RECT 1.330 0.915 1.500 2.635 ;
        RECT 1.145 2.465 1.500 2.635 ;
        RECT 1.330 0.915 3.150 1.085 ;
        RECT 2.980 0.550 3.150 1.585 ;
        RECT 3.080 1.415 3.250 2.630 ;
        RECT 2.980 0.550 3.775 0.720 ;
        RECT 5.850 0.535 6.020 2.630 ;
        RECT 5.850 0.535 6.180 0.705 ;
        RECT 3.080 2.460 6.645 2.630 ;
        RECT 6.875 1.195 7.900 1.365 ;
        RECT 7.730 0.550 7.900 2.775 ;
        RECT 7.595 2.605 7.900 2.775 ;
        RECT 7.730 1.630 8.120 1.800 ;
        RECT 6.200 0.900 6.370 2.280 ;
        RECT 7.245 1.675 7.415 3.125 ;
        RECT 6.200 1.675 7.550 1.845 ;
        RECT 8.080 2.460 8.250 3.125 ;
        RECT 7.245 2.955 8.250 3.125 ;
        RECT 8.740 1.610 8.910 2.630 ;
        RECT 8.080 2.460 8.910 2.630 ;
  END 
END FFDCRHDLXHT

MACRO FFDCRHD2XHT
  CLASS  CORE ;
  FOREIGN FFDCRHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.800 0.720 9.970 2.960 ;
        RECT 9.800 1.645 10.150 2.015 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.725 0.720 8.930 2.280 ;
        RECT 8.710 1.575 8.930 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.665 1.265 2.090 1.780 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.345 1.265 2.785 1.780 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.675 -0.300 0.975 0.995 ;
        RECT 1.800 -0.300 2.100 0.735 ;
        RECT 4.300 -0.300 4.600 1.020 ;
        RECT 5.285 -0.300 5.585 0.715 ;
        RECT 7.030 -0.300 7.200 0.780 ;
        RECT 8.375 -0.300 8.545 1.360 ;
        RECT 8.240 1.060 8.545 1.360 ;
        RECT 9.215 -0.300 9.515 1.055 ;
        RECT 10.255 -0.300 10.555 1.055 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.545 0.520 2.010 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 2.810 0.835 3.990 ;
        RECT 2.145 2.810 2.445 3.990 ;
        RECT 4.270 3.095 4.570 3.990 ;
        RECT 5.180 3.095 5.480 3.990 ;
        RECT 7.105 2.795 7.275 3.990 ;
        RECT 8.175 2.975 8.475 3.990 ;
        RECT 9.215 2.975 9.515 3.990 ;
        RECT 10.255 2.295 10.555 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.660 1.980 2.810 2.280 ;
        RECT 3.320 0.950 3.665 1.120 ;
        RECT 3.495 0.950 3.665 2.215 ;
        RECT 3.365 2.045 3.665 2.215 ;
        RECT 3.495 1.675 4.840 1.845 ;
        RECT 4.040 1.275 5.190 1.445 ;
        RECT 4.905 0.985 5.075 1.445 ;
        RECT 5.020 1.275 5.190 2.215 ;
        RECT 4.840 2.045 5.190 2.215 ;
        RECT 5.020 1.585 5.675 1.755 ;
        RECT 0.105 1.125 0.405 1.345 ;
        RECT 0.105 1.175 0.885 1.345 ;
        RECT 0.105 2.190 0.885 2.360 ;
        RECT 0.715 1.175 0.885 2.630 ;
        RECT 0.715 1.525 1.020 1.825 ;
        RECT 0.715 2.460 2.810 2.630 ;
        RECT 2.640 2.460 2.810 2.915 ;
        RECT 3.690 2.745 3.990 2.990 ;
        RECT 2.640 2.745 6.240 2.915 ;
        RECT 6.070 2.745 6.240 3.210 ;
        RECT 6.070 3.040 6.755 3.210 ;
        RECT 2.965 1.605 3.205 1.885 ;
        RECT 1.290 0.915 1.460 2.215 ;
        RECT 1.085 2.045 1.460 2.215 ;
        RECT 1.290 0.915 3.135 1.085 ;
        RECT 2.965 0.480 3.135 1.885 ;
        RECT 2.990 1.605 3.185 2.565 ;
        RECT 2.990 1.605 3.205 1.905 ;
        RECT 2.965 0.480 3.890 0.650 ;
        RECT 5.855 0.695 6.025 2.565 ;
        RECT 2.990 2.395 6.755 2.565 ;
        RECT 5.855 0.695 6.795 0.865 ;
        RECT 6.455 2.395 6.755 2.730 ;
        RECT 6.625 0.695 6.795 1.140 ;
        RECT 7.380 0.480 7.550 1.140 ;
        RECT 6.625 0.970 7.550 1.140 ;
        RECT 7.380 0.480 8.195 0.650 ;
        RECT 6.945 1.675 7.900 1.845 ;
        RECT 7.730 1.060 7.900 2.280 ;
        RECT 7.730 1.595 8.530 1.765 ;
        RECT 6.270 1.060 6.440 2.215 ;
        RECT 6.205 2.045 7.550 2.215 ;
        RECT 7.380 2.045 7.550 2.630 ;
        RECT 7.455 2.460 7.625 3.185 ;
        RECT 7.455 3.010 7.755 3.185 ;
        RECT 9.450 1.525 9.620 2.630 ;
        RECT 7.380 2.460 9.620 2.630 ;
  END 
END FFDCRHD2XHT

MACRO FFDCRHD1XHT
  CLASS  CORE ;
  FOREIGN FFDCRHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.840 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.500 0.720 9.740 2.960 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.460 0.720 8.630 1.480 ;
        RECT 8.460 1.300 8.920 1.480 ;
        RECT 8.710 1.300 8.920 2.215 ;
        RECT 8.395 2.045 8.920 2.215 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.680 1.290 2.105 1.780 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.435 1.265 2.820 1.780 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.670 -0.300 0.970 0.945 ;
        RECT 1.890 -0.300 2.190 0.735 ;
        RECT 4.270 -0.300 4.570 1.020 ;
        RECT 5.360 -0.300 5.660 1.075 ;
        RECT 7.260 -0.300 7.560 0.995 ;
        RECT 8.915 -0.300 9.215 1.055 ;
        RECT 0.000 -0.300 9.840 0.300 ;
    END
  END GND
  PIN CK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.525 0.550 2.015 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.580 2.810 0.880 3.990 ;
        RECT 2.190 2.810 2.490 3.990 ;
        RECT 4.270 3.160 4.570 3.990 ;
        RECT 5.360 3.160 5.660 3.990 ;
        RECT 7.260 2.810 7.560 3.990 ;
        RECT 8.915 2.975 9.215 3.990 ;
        RECT 0.000 3.390 9.840 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.705 1.980 2.915 2.280 ;
        RECT 3.385 1.030 3.615 1.200 ;
        RECT 3.385 0.900 3.555 1.200 ;
        RECT 3.445 1.030 3.615 2.280 ;
        RECT 3.445 1.675 4.755 1.845 ;
        RECT 4.850 0.850 5.150 1.020 ;
        RECT 4.040 1.220 5.150 1.390 ;
        RECT 4.980 0.850 5.150 2.215 ;
        RECT 4.850 2.045 5.150 2.215 ;
        RECT 4.980 1.535 5.845 1.705 ;
        RECT 0.105 1.125 0.950 1.295 ;
        RECT 0.105 2.195 0.950 2.365 ;
        RECT 0.780 1.125 0.950 2.630 ;
        RECT 0.780 1.525 1.085 1.825 ;
        RECT 0.780 2.460 2.915 2.630 ;
        RECT 2.745 2.460 2.915 3.075 ;
        RECT 3.680 2.810 3.900 3.075 ;
        RECT 2.745 2.905 3.900 3.075 ;
        RECT 3.680 2.810 6.370 2.980 ;
        RECT 3.035 1.415 3.265 1.585 ;
        RECT 1.265 0.915 1.435 2.215 ;
        RECT 1.130 2.045 1.435 2.215 ;
        RECT 1.265 0.915 1.500 1.360 ;
        RECT 1.265 0.915 3.205 1.085 ;
        RECT 3.035 0.480 3.205 1.585 ;
        RECT 3.095 1.415 3.265 2.725 ;
        RECT 3.095 2.460 3.410 2.725 ;
        RECT 3.035 0.480 3.830 0.650 ;
        RECT 6.025 0.535 6.195 2.630 ;
        RECT 6.025 0.535 6.360 0.705 ;
        RECT 3.095 2.460 6.795 2.630 ;
        RECT 6.625 2.460 6.795 2.770 ;
        RECT 7.050 1.195 8.120 1.365 ;
        RECT 7.860 0.760 8.030 1.365 ;
        RECT 7.950 1.195 8.120 2.280 ;
        RECT 7.950 1.660 8.530 1.830 ;
        RECT 6.375 0.900 6.545 2.280 ;
        RECT 6.375 1.675 7.725 1.845 ;
        RECT 7.555 1.675 7.725 2.630 ;
        RECT 9.150 1.610 9.320 2.630 ;
        RECT 7.555 2.460 9.320 2.630 ;
  END 
END FFDCRHD1XHT

MACRO FAHHDMXHT
  CLASS  CORE ;
  FOREIGN FAHHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.250 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.485 0.720 1.820 ;
        RECT 0.510 1.485 0.720 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.135 1.275 4.475 1.840 ;
    END
  END B
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.905 1.060 10.160 1.360 ;
        RECT 9.990 1.060 10.160 2.865 ;
        RECT 9.905 2.100 10.160 2.865 ;
    END
  END S
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.815 1.245 8.100 1.820 ;
    END
  END CI
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.955 ;
        RECT 3.950 -0.300 4.250 0.665 ;
        RECT 7.615 -0.300 7.915 0.550 ;
        RECT 9.370 -0.300 9.540 0.665 ;
        RECT 0.000 -0.300 10.250 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.985 0.955 3.990 ;
        RECT 3.825 2.985 4.125 3.990 ;
        RECT 7.645 3.095 7.945 3.990 ;
        RECT 9.290 2.905 9.590 3.990 ;
        RECT 0.000 3.390 10.250 3.990 ;
    END
  END VDD
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.710 1.060 8.960 2.215 ;
        RECT 8.710 2.045 9.050 2.215 ;
    END
  END CO
  OBS 
      LAYER M1 ;
        RECT 1.270 1.060 1.505 1.360 ;
        RECT 1.315 1.060 1.505 2.455 ;
        RECT 1.205 2.285 1.505 2.455 ;
        RECT 0.090 1.125 0.260 2.805 ;
        RECT 0.090 2.110 0.340 2.805 ;
        RECT 0.090 1.125 0.405 1.305 ;
        RECT 0.090 1.135 1.090 1.305 ;
        RECT 0.920 1.135 1.090 1.850 ;
        RECT 2.310 1.060 2.480 2.805 ;
        RECT 0.090 2.635 2.480 2.805 ;
        RECT 1.235 2.985 3.615 3.155 ;
        RECT 3.180 1.125 3.350 2.455 ;
        RECT 3.180 2.285 3.585 2.455 ;
        RECT 3.180 1.125 3.615 1.295 ;
        RECT 3.530 1.625 3.935 1.795 ;
        RECT 3.765 1.625 3.935 2.250 ;
        RECT 4.820 0.855 4.990 2.250 ;
        RECT 3.765 2.045 4.990 2.250 ;
        RECT 3.765 2.055 5.310 2.250 ;
        RECT 1.790 0.710 1.960 2.455 ;
        RECT 1.725 2.280 2.025 2.455 ;
        RECT 1.790 0.710 3.635 0.880 ;
        RECT 4.470 0.500 4.640 1.020 ;
        RECT 3.850 0.850 4.640 1.020 ;
        RECT 4.470 0.500 5.395 0.670 ;
        RECT 3.775 0.785 3.785 1.019 ;
        RECT 3.785 0.795 3.795 1.019 ;
        RECT 3.795 0.805 3.805 1.019 ;
        RECT 3.805 0.815 3.815 1.019 ;
        RECT 3.815 0.825 3.825 1.019 ;
        RECT 3.825 0.835 3.835 1.019 ;
        RECT 3.835 0.845 3.845 1.019 ;
        RECT 3.845 0.850 3.851 1.020 ;
        RECT 3.710 0.720 3.720 0.954 ;
        RECT 3.720 0.730 3.730 0.964 ;
        RECT 3.730 0.740 3.740 0.974 ;
        RECT 3.740 0.750 3.750 0.984 ;
        RECT 3.750 0.760 3.760 0.994 ;
        RECT 3.760 0.770 3.770 1.004 ;
        RECT 3.770 0.775 3.776 1.015 ;
        RECT 3.635 0.710 3.645 0.880 ;
        RECT 3.645 0.710 3.655 0.890 ;
        RECT 3.655 0.710 3.665 0.900 ;
        RECT 3.665 0.710 3.675 0.910 ;
        RECT 3.675 0.710 3.685 0.920 ;
        RECT 3.685 0.710 3.695 0.930 ;
        RECT 3.695 0.710 3.705 0.940 ;
        RECT 3.705 0.710 3.711 0.950 ;
        RECT 2.830 1.060 3.000 2.805 ;
        RECT 3.890 2.480 4.060 2.805 ;
        RECT 2.830 2.635 4.060 2.805 ;
        RECT 3.890 2.480 5.490 2.650 ;
        RECT 5.935 2.675 6.105 3.030 ;
        RECT 4.640 2.860 6.105 3.030 ;
        RECT 7.185 1.060 7.355 2.215 ;
        RECT 7.120 2.045 7.420 2.215 ;
        RECT 8.280 1.060 8.450 2.215 ;
        RECT 8.215 2.045 8.515 2.215 ;
        RECT 6.115 2.225 6.455 2.395 ;
        RECT 6.115 0.920 6.285 2.395 ;
        RECT 6.050 0.920 6.350 1.090 ;
        RECT 6.285 2.225 6.455 2.915 ;
        RECT 6.285 2.745 8.540 2.915 ;
        RECT 5.405 0.920 5.765 1.090 ;
        RECT 5.595 0.570 5.765 2.315 ;
        RECT 5.595 0.570 7.295 0.740 ;
        RECT 7.625 0.820 7.925 0.990 ;
        RECT 8.110 0.710 9.040 0.880 ;
        RECT 9.155 0.760 9.165 1.814 ;
        RECT 9.165 0.770 9.175 1.814 ;
        RECT 9.175 0.780 9.185 1.814 ;
        RECT 9.185 0.790 9.195 1.814 ;
        RECT 9.195 0.800 9.205 1.814 ;
        RECT 9.205 0.810 9.215 1.814 ;
        RECT 9.215 0.820 9.225 1.814 ;
        RECT 9.225 0.830 9.235 1.814 ;
        RECT 9.235 0.840 9.245 1.814 ;
        RECT 9.245 0.850 9.255 1.814 ;
        RECT 9.255 0.860 9.265 1.814 ;
        RECT 9.265 0.870 9.275 1.814 ;
        RECT 9.275 0.880 9.285 1.814 ;
        RECT 9.285 0.890 9.295 1.814 ;
        RECT 9.295 0.900 9.305 1.814 ;
        RECT 9.305 0.910 9.315 1.814 ;
        RECT 9.315 0.920 9.325 1.814 ;
        RECT 9.115 0.720 9.125 0.954 ;
        RECT 9.125 0.730 9.135 0.964 ;
        RECT 9.135 0.740 9.145 0.974 ;
        RECT 9.145 0.750 9.155 0.984 ;
        RECT 9.040 0.710 9.050 0.880 ;
        RECT 9.050 0.710 9.060 0.890 ;
        RECT 9.060 0.710 9.070 0.900 ;
        RECT 9.070 0.710 9.080 0.910 ;
        RECT 9.080 0.710 9.090 0.920 ;
        RECT 9.090 0.710 9.100 0.930 ;
        RECT 9.100 0.710 9.110 0.940 ;
        RECT 9.110 0.710 9.116 0.950 ;
        RECT 8.035 0.710 8.045 0.944 ;
        RECT 8.045 0.710 8.055 0.934 ;
        RECT 8.055 0.710 8.065 0.924 ;
        RECT 8.065 0.710 8.075 0.914 ;
        RECT 8.075 0.710 8.085 0.904 ;
        RECT 8.085 0.710 8.095 0.894 ;
        RECT 8.095 0.710 8.105 0.884 ;
        RECT 8.105 0.710 8.111 0.880 ;
        RECT 8.000 0.745 8.010 0.979 ;
        RECT 8.010 0.735 8.020 0.969 ;
        RECT 8.020 0.725 8.030 0.959 ;
        RECT 8.030 0.715 8.036 0.955 ;
        RECT 7.925 0.820 7.935 0.990 ;
        RECT 7.935 0.810 7.945 0.990 ;
        RECT 7.945 0.800 7.955 0.990 ;
        RECT 7.955 0.790 7.965 0.990 ;
        RECT 7.965 0.780 7.975 0.990 ;
        RECT 7.975 0.770 7.985 0.990 ;
        RECT 7.985 0.760 7.995 0.990 ;
        RECT 7.995 0.750 8.001 0.990 ;
        RECT 7.545 0.750 7.555 0.990 ;
        RECT 7.555 0.760 7.565 0.990 ;
        RECT 7.565 0.770 7.575 0.990 ;
        RECT 7.575 0.780 7.585 0.990 ;
        RECT 7.585 0.790 7.595 0.990 ;
        RECT 7.595 0.800 7.605 0.990 ;
        RECT 7.605 0.810 7.615 0.990 ;
        RECT 7.615 0.820 7.625 0.990 ;
        RECT 7.375 0.580 7.385 0.820 ;
        RECT 7.385 0.590 7.395 0.830 ;
        RECT 7.395 0.600 7.405 0.840 ;
        RECT 7.405 0.610 7.415 0.850 ;
        RECT 7.415 0.620 7.425 0.860 ;
        RECT 7.425 0.630 7.435 0.870 ;
        RECT 7.435 0.640 7.445 0.880 ;
        RECT 7.445 0.650 7.455 0.890 ;
        RECT 7.455 0.660 7.465 0.900 ;
        RECT 7.465 0.670 7.475 0.910 ;
        RECT 7.475 0.680 7.485 0.920 ;
        RECT 7.485 0.690 7.495 0.930 ;
        RECT 7.495 0.700 7.505 0.940 ;
        RECT 7.505 0.710 7.515 0.950 ;
        RECT 7.515 0.720 7.525 0.960 ;
        RECT 7.525 0.730 7.535 0.970 ;
        RECT 7.535 0.740 7.545 0.980 ;
        RECT 7.295 0.570 7.305 0.740 ;
        RECT 7.305 0.570 7.315 0.750 ;
        RECT 7.315 0.570 7.325 0.760 ;
        RECT 7.325 0.570 7.335 0.770 ;
        RECT 7.335 0.570 7.345 0.780 ;
        RECT 7.345 0.570 7.355 0.790 ;
        RECT 7.355 0.570 7.365 0.800 ;
        RECT 7.365 0.570 7.375 0.810 ;
        RECT 6.635 0.920 6.805 2.565 ;
        RECT 6.570 0.920 6.870 1.090 ;
        RECT 9.545 1.520 9.715 2.565 ;
        RECT 6.635 2.395 9.715 2.565 ;
        RECT 9.545 1.520 9.805 1.820 ;
  END 
END FAHHDMXHT

MACRO FAHHD2XHT
  CLASS  CORE ;
  FOREIGN FAHHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.480 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.485 0.720 1.820 ;
        RECT 0.510 1.485 0.720 2.045 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.135 1.285 4.485 1.840 ;
    END
  END B
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.285 2.560 10.655 2.770 ;
        RECT 10.455 0.720 10.655 2.960 ;
    END
  END S
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.760 1.265 8.100 1.820 ;
    END
  END CI
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.955 ;
        RECT 3.985 -0.300 4.285 0.665 ;
        RECT 7.680 -0.300 7.850 0.615 ;
        RECT 8.810 -0.300 9.110 0.660 ;
        RECT 9.880 -0.300 10.180 1.055 ;
        RECT 10.930 -0.300 11.230 1.055 ;
        RECT 0.000 -0.300 11.480 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.985 0.955 3.990 ;
        RECT 3.825 2.985 4.125 3.990 ;
        RECT 7.645 3.095 7.945 3.990 ;
        RECT 8.835 2.975 9.135 3.990 ;
        RECT 9.880 2.975 10.185 3.990 ;
        RECT 10.925 2.295 11.225 3.990 ;
        RECT 0.000 3.390 11.480 3.990 ;
    END
  END VDD
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.425 0.720 9.660 2.215 ;
        RECT 9.360 2.045 9.660 2.215 ;
        RECT 9.425 1.265 9.750 1.610 ;
    END
  END CO
  OBS 
      LAYER M1 ;
        RECT 1.270 1.060 1.505 1.360 ;
        RECT 1.315 1.060 1.505 2.455 ;
        RECT 1.205 2.285 1.505 2.455 ;
        RECT 0.090 1.125 0.260 2.805 ;
        RECT 0.090 2.110 0.340 2.805 ;
        RECT 0.090 1.125 0.445 1.305 ;
        RECT 0.090 1.135 1.090 1.305 ;
        RECT 0.920 1.135 1.090 1.850 ;
        RECT 2.310 1.060 2.480 2.805 ;
        RECT 0.090 2.635 2.480 2.805 ;
        RECT 3.180 1.125 3.350 2.455 ;
        RECT 3.180 1.125 3.585 1.295 ;
        RECT 3.180 2.285 3.585 2.455 ;
        RECT 1.235 2.985 3.615 3.155 ;
        RECT 3.530 1.625 3.935 1.795 ;
        RECT 3.765 1.625 3.935 2.230 ;
        RECT 4.815 0.935 4.985 2.230 ;
        RECT 3.765 2.045 4.985 2.230 ;
        RECT 3.765 2.055 5.310 2.230 ;
        RECT 5.010 2.055 5.310 2.315 ;
        RECT 1.790 0.635 1.960 2.455 ;
        RECT 1.725 2.285 2.025 2.455 ;
        RECT 1.790 0.635 3.535 0.805 ;
        RECT 4.465 0.480 4.635 1.025 ;
        RECT 3.830 0.855 4.635 1.025 ;
        RECT 4.465 0.480 5.395 0.650 ;
        RECT 3.755 0.790 3.765 1.024 ;
        RECT 3.765 0.800 3.775 1.024 ;
        RECT 3.775 0.810 3.785 1.024 ;
        RECT 3.785 0.820 3.795 1.024 ;
        RECT 3.795 0.830 3.805 1.024 ;
        RECT 3.805 0.840 3.815 1.024 ;
        RECT 3.815 0.850 3.825 1.024 ;
        RECT 3.825 0.855 3.831 1.025 ;
        RECT 3.610 0.645 3.620 0.879 ;
        RECT 3.620 0.655 3.630 0.889 ;
        RECT 3.630 0.665 3.640 0.899 ;
        RECT 3.640 0.675 3.650 0.909 ;
        RECT 3.650 0.685 3.660 0.919 ;
        RECT 3.660 0.695 3.670 0.929 ;
        RECT 3.670 0.705 3.680 0.939 ;
        RECT 3.680 0.715 3.690 0.949 ;
        RECT 3.690 0.725 3.700 0.959 ;
        RECT 3.700 0.735 3.710 0.969 ;
        RECT 3.710 0.745 3.720 0.979 ;
        RECT 3.720 0.755 3.730 0.989 ;
        RECT 3.730 0.765 3.740 0.999 ;
        RECT 3.740 0.775 3.750 1.009 ;
        RECT 3.750 0.780 3.756 1.020 ;
        RECT 3.535 0.635 3.545 0.805 ;
        RECT 3.545 0.635 3.555 0.815 ;
        RECT 3.555 0.635 3.565 0.825 ;
        RECT 3.565 0.635 3.575 0.835 ;
        RECT 3.575 0.635 3.585 0.845 ;
        RECT 3.585 0.635 3.595 0.855 ;
        RECT 3.595 0.635 3.605 0.865 ;
        RECT 3.605 0.635 3.611 0.875 ;
        RECT 2.830 1.060 3.000 2.805 ;
        RECT 2.830 2.635 5.490 2.805 ;
        RECT 5.190 2.635 5.490 2.840 ;
        RECT 4.905 2.985 5.075 3.190 ;
        RECT 4.640 2.985 5.075 3.155 ;
        RECT 5.670 2.970 5.840 3.190 ;
        RECT 4.905 3.020 5.840 3.190 ;
        RECT 5.670 2.970 6.170 3.140 ;
        RECT 7.185 1.060 7.355 2.215 ;
        RECT 7.120 2.045 7.420 2.215 ;
        RECT 8.280 1.060 8.455 2.215 ;
        RECT 8.195 2.045 8.495 2.215 ;
        RECT 6.115 0.935 6.285 2.420 ;
        RECT 6.560 2.745 8.525 2.915 ;
        RECT 6.480 2.675 6.490 2.915 ;
        RECT 6.490 2.685 6.500 2.915 ;
        RECT 6.500 2.695 6.510 2.915 ;
        RECT 6.510 2.705 6.520 2.915 ;
        RECT 6.520 2.715 6.530 2.915 ;
        RECT 6.530 2.725 6.540 2.915 ;
        RECT 6.540 2.735 6.550 2.915 ;
        RECT 6.550 2.745 6.560 2.915 ;
        RECT 6.455 2.650 6.465 2.890 ;
        RECT 6.465 2.660 6.475 2.900 ;
        RECT 6.475 2.665 6.481 2.909 ;
        RECT 6.285 2.250 6.295 2.720 ;
        RECT 6.295 2.250 6.305 2.730 ;
        RECT 6.305 2.250 6.315 2.740 ;
        RECT 6.315 2.250 6.325 2.750 ;
        RECT 6.325 2.250 6.335 2.760 ;
        RECT 6.335 2.250 6.345 2.770 ;
        RECT 6.345 2.250 6.355 2.780 ;
        RECT 6.355 2.250 6.365 2.790 ;
        RECT 6.365 2.250 6.375 2.800 ;
        RECT 6.375 2.250 6.385 2.810 ;
        RECT 6.385 2.250 6.395 2.820 ;
        RECT 6.395 2.250 6.405 2.830 ;
        RECT 6.405 2.250 6.415 2.840 ;
        RECT 6.415 2.250 6.425 2.850 ;
        RECT 6.425 2.250 6.435 2.860 ;
        RECT 6.435 2.250 6.445 2.870 ;
        RECT 6.445 2.250 6.455 2.880 ;
        RECT 5.400 1.000 5.765 1.170 ;
        RECT 5.595 0.585 5.765 2.395 ;
        RECT 5.595 0.585 7.310 0.755 ;
        RECT 7.625 0.820 7.925 0.990 ;
        RECT 8.145 0.675 8.495 0.845 ;
        RECT 8.900 1.525 9.245 1.825 ;
        RECT 8.730 0.845 8.740 1.825 ;
        RECT 8.740 0.855 8.750 1.825 ;
        RECT 8.750 0.865 8.760 1.825 ;
        RECT 8.760 0.875 8.770 1.825 ;
        RECT 8.770 0.885 8.780 1.825 ;
        RECT 8.780 0.895 8.790 1.825 ;
        RECT 8.790 0.905 8.800 1.825 ;
        RECT 8.800 0.915 8.810 1.825 ;
        RECT 8.810 0.925 8.820 1.825 ;
        RECT 8.820 0.935 8.830 1.825 ;
        RECT 8.830 0.945 8.840 1.825 ;
        RECT 8.840 0.955 8.850 1.825 ;
        RECT 8.850 0.965 8.860 1.825 ;
        RECT 8.860 0.975 8.870 1.825 ;
        RECT 8.870 0.985 8.880 1.825 ;
        RECT 8.880 0.995 8.890 1.825 ;
        RECT 8.890 1.005 8.900 1.825 ;
        RECT 8.570 0.685 8.580 0.919 ;
        RECT 8.580 0.695 8.590 0.929 ;
        RECT 8.590 0.705 8.600 0.939 ;
        RECT 8.600 0.715 8.610 0.949 ;
        RECT 8.610 0.725 8.620 0.959 ;
        RECT 8.620 0.735 8.630 0.969 ;
        RECT 8.630 0.745 8.640 0.979 ;
        RECT 8.640 0.755 8.650 0.989 ;
        RECT 8.650 0.765 8.660 0.999 ;
        RECT 8.660 0.775 8.670 1.009 ;
        RECT 8.670 0.785 8.680 1.019 ;
        RECT 8.680 0.795 8.690 1.029 ;
        RECT 8.690 0.805 8.700 1.039 ;
        RECT 8.700 0.815 8.710 1.049 ;
        RECT 8.710 0.825 8.720 1.059 ;
        RECT 8.720 0.835 8.730 1.069 ;
        RECT 8.495 0.675 8.505 0.845 ;
        RECT 8.505 0.675 8.515 0.855 ;
        RECT 8.515 0.675 8.525 0.865 ;
        RECT 8.525 0.675 8.535 0.875 ;
        RECT 8.535 0.675 8.545 0.885 ;
        RECT 8.545 0.675 8.555 0.895 ;
        RECT 8.555 0.675 8.565 0.905 ;
        RECT 8.565 0.675 8.571 0.915 ;
        RECT 8.070 0.675 8.080 0.909 ;
        RECT 8.080 0.675 8.090 0.899 ;
        RECT 8.090 0.675 8.100 0.889 ;
        RECT 8.100 0.675 8.110 0.879 ;
        RECT 8.110 0.675 8.120 0.869 ;
        RECT 8.120 0.675 8.130 0.859 ;
        RECT 8.130 0.675 8.140 0.849 ;
        RECT 8.140 0.675 8.146 0.845 ;
        RECT 8.000 0.745 8.010 0.979 ;
        RECT 8.010 0.735 8.020 0.969 ;
        RECT 8.020 0.725 8.030 0.959 ;
        RECT 8.030 0.715 8.040 0.949 ;
        RECT 8.040 0.705 8.050 0.939 ;
        RECT 8.050 0.695 8.060 0.929 ;
        RECT 8.060 0.685 8.070 0.919 ;
        RECT 7.925 0.820 7.935 0.990 ;
        RECT 7.935 0.810 7.945 0.990 ;
        RECT 7.945 0.800 7.955 0.990 ;
        RECT 7.955 0.790 7.965 0.990 ;
        RECT 7.965 0.780 7.975 0.990 ;
        RECT 7.975 0.770 7.985 0.990 ;
        RECT 7.985 0.760 7.995 0.990 ;
        RECT 7.995 0.750 8.001 0.990 ;
        RECT 7.545 0.750 7.555 0.990 ;
        RECT 7.555 0.760 7.565 0.990 ;
        RECT 7.565 0.770 7.575 0.990 ;
        RECT 7.575 0.780 7.585 0.990 ;
        RECT 7.585 0.790 7.595 0.990 ;
        RECT 7.595 0.800 7.605 0.990 ;
        RECT 7.605 0.810 7.615 0.990 ;
        RECT 7.615 0.820 7.625 0.990 ;
        RECT 7.390 0.595 7.400 0.835 ;
        RECT 7.400 0.605 7.410 0.845 ;
        RECT 7.410 0.615 7.420 0.855 ;
        RECT 7.420 0.625 7.430 0.865 ;
        RECT 7.430 0.635 7.440 0.875 ;
        RECT 7.440 0.645 7.450 0.885 ;
        RECT 7.450 0.655 7.460 0.895 ;
        RECT 7.460 0.665 7.470 0.905 ;
        RECT 7.470 0.675 7.480 0.915 ;
        RECT 7.480 0.685 7.490 0.925 ;
        RECT 7.490 0.695 7.500 0.935 ;
        RECT 7.500 0.705 7.510 0.945 ;
        RECT 7.510 0.715 7.520 0.955 ;
        RECT 7.520 0.725 7.530 0.965 ;
        RECT 7.530 0.735 7.540 0.975 ;
        RECT 7.540 0.740 7.546 0.984 ;
        RECT 7.310 0.585 7.320 0.755 ;
        RECT 7.320 0.585 7.330 0.765 ;
        RECT 7.330 0.585 7.340 0.775 ;
        RECT 7.340 0.585 7.350 0.785 ;
        RECT 7.350 0.585 7.360 0.795 ;
        RECT 7.360 0.585 7.370 0.805 ;
        RECT 7.370 0.585 7.380 0.815 ;
        RECT 7.380 0.585 7.390 0.825 ;
        RECT 6.635 0.935 6.805 2.565 ;
        RECT 9.935 1.610 10.105 2.565 ;
        RECT 6.635 2.395 10.105 2.565 ;
        RECT 9.935 1.610 10.270 1.910 ;
  END 
END FAHHD2XHT

MACRO FAHHD1XHT
  CLASS  CORE ;
  FOREIGN FAHHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.250 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.485 0.720 1.820 ;
        RECT 0.510 1.485 0.720 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.155 1.265 4.435 1.865 ;
    END
  END B
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.905 0.720 10.150 1.360 ;
        RECT 9.970 0.720 10.150 2.960 ;
        RECT 9.905 1.980 10.150 2.960 ;
    END
  END S
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.695 1.500 8.100 2.025 ;
    END
  END CI
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.955 ;
        RECT 4.015 -0.300 4.315 0.665 ;
        RECT 7.680 -0.300 7.850 0.615 ;
        RECT 9.355 -0.300 9.525 0.660 ;
        RECT 0.000 -0.300 10.250 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.985 0.955 3.990 ;
        RECT 3.825 2.985 4.125 3.990 ;
        RECT 7.645 3.095 7.945 3.990 ;
        RECT 9.320 2.975 9.620 3.990 ;
        RECT 0.000 3.390 10.250 3.990 ;
    END
  END VDD
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 8.710 1.530 8.960 1.700 ;
        RECT 8.790 1.060 8.945 2.215 ;
        RECT 8.710 1.060 8.945 1.700 ;
        RECT 8.790 1.530 8.960 2.215 ;
        RECT 8.790 2.045 9.115 2.215 ;
    END
  END CO
  OBS 
      LAYER M1 ;
        RECT 1.270 1.060 1.505 1.360 ;
        RECT 1.315 1.060 1.505 2.455 ;
        RECT 1.205 2.285 1.505 2.455 ;
        RECT 0.090 1.125 0.260 2.805 ;
        RECT 0.090 2.110 0.340 2.805 ;
        RECT 0.090 1.125 0.405 1.305 ;
        RECT 0.090 1.135 1.090 1.305 ;
        RECT 0.920 1.135 1.090 1.850 ;
        RECT 2.310 1.060 2.480 2.805 ;
        RECT 0.090 2.635 2.480 2.805 ;
        RECT 1.235 2.985 3.615 3.155 ;
        RECT 3.180 1.125 3.350 2.455 ;
        RECT 3.180 2.285 3.585 2.455 ;
        RECT 3.180 1.125 3.615 1.295 ;
        RECT 3.530 1.625 3.935 1.795 ;
        RECT 3.765 1.625 3.935 2.255 ;
        RECT 4.845 0.855 5.015 2.255 ;
        RECT 4.845 2.055 5.310 2.255 ;
        RECT 3.765 2.085 5.310 2.255 ;
        RECT 1.790 0.635 1.960 2.455 ;
        RECT 1.725 2.285 2.025 2.455 ;
        RECT 1.790 0.635 3.555 0.805 ;
        RECT 4.495 0.480 4.665 1.025 ;
        RECT 3.850 0.855 4.665 1.025 ;
        RECT 4.495 0.480 5.395 0.650 ;
        RECT 3.775 0.790 3.785 1.024 ;
        RECT 3.785 0.800 3.795 1.024 ;
        RECT 3.795 0.810 3.805 1.024 ;
        RECT 3.805 0.820 3.815 1.024 ;
        RECT 3.815 0.830 3.825 1.024 ;
        RECT 3.825 0.840 3.835 1.024 ;
        RECT 3.835 0.850 3.845 1.024 ;
        RECT 3.845 0.855 3.851 1.025 ;
        RECT 3.630 0.645 3.640 0.879 ;
        RECT 3.640 0.655 3.650 0.889 ;
        RECT 3.650 0.665 3.660 0.899 ;
        RECT 3.660 0.675 3.670 0.909 ;
        RECT 3.670 0.685 3.680 0.919 ;
        RECT 3.680 0.695 3.690 0.929 ;
        RECT 3.690 0.705 3.700 0.939 ;
        RECT 3.700 0.715 3.710 0.949 ;
        RECT 3.710 0.725 3.720 0.959 ;
        RECT 3.720 0.735 3.730 0.969 ;
        RECT 3.730 0.745 3.740 0.979 ;
        RECT 3.740 0.755 3.750 0.989 ;
        RECT 3.750 0.765 3.760 0.999 ;
        RECT 3.760 0.775 3.770 1.009 ;
        RECT 3.770 0.780 3.776 1.020 ;
        RECT 3.555 0.635 3.565 0.805 ;
        RECT 3.565 0.635 3.575 0.815 ;
        RECT 3.575 0.635 3.585 0.825 ;
        RECT 3.585 0.635 3.595 0.835 ;
        RECT 3.595 0.635 3.605 0.845 ;
        RECT 3.605 0.635 3.615 0.855 ;
        RECT 3.615 0.635 3.625 0.865 ;
        RECT 3.625 0.635 3.631 0.875 ;
        RECT 2.830 1.060 3.000 2.805 ;
        RECT 3.890 2.480 4.060 2.805 ;
        RECT 2.830 2.635 4.060 2.805 ;
        RECT 3.890 2.480 5.490 2.650 ;
        RECT 4.640 2.860 5.935 3.030 ;
        RECT 5.765 2.830 5.935 3.130 ;
        RECT 7.185 1.060 7.355 2.215 ;
        RECT 7.120 2.045 7.420 2.215 ;
        RECT 6.115 0.920 6.285 2.915 ;
        RECT 6.050 0.920 6.350 1.090 ;
        RECT 6.115 2.745 8.525 2.915 ;
        RECT 8.280 1.125 8.450 2.215 ;
        RECT 8.200 1.125 8.500 1.295 ;
        RECT 8.280 2.045 8.580 2.215 ;
        RECT 5.420 0.920 5.765 1.090 ;
        RECT 5.595 0.570 5.765 2.320 ;
        RECT 5.595 0.570 7.295 0.740 ;
        RECT 7.600 0.795 7.950 0.965 ;
        RECT 8.190 0.630 8.945 0.800 ;
        RECT 9.140 0.760 9.150 1.840 ;
        RECT 9.150 0.770 9.160 1.840 ;
        RECT 9.160 0.780 9.170 1.840 ;
        RECT 9.170 0.790 9.180 1.840 ;
        RECT 9.180 0.800 9.190 1.840 ;
        RECT 9.190 0.810 9.200 1.840 ;
        RECT 9.200 0.820 9.210 1.840 ;
        RECT 9.210 0.830 9.220 1.840 ;
        RECT 9.220 0.840 9.230 1.840 ;
        RECT 9.230 0.850 9.240 1.840 ;
        RECT 9.240 0.860 9.250 1.840 ;
        RECT 9.250 0.870 9.260 1.840 ;
        RECT 9.260 0.880 9.270 1.840 ;
        RECT 9.270 0.890 9.280 1.840 ;
        RECT 9.280 0.900 9.290 1.840 ;
        RECT 9.290 0.910 9.300 1.840 ;
        RECT 9.300 0.920 9.310 1.840 ;
        RECT 9.020 0.640 9.030 0.874 ;
        RECT 9.030 0.650 9.040 0.884 ;
        RECT 9.040 0.660 9.050 0.894 ;
        RECT 9.050 0.670 9.060 0.904 ;
        RECT 9.060 0.680 9.070 0.914 ;
        RECT 9.070 0.690 9.080 0.924 ;
        RECT 9.080 0.700 9.090 0.934 ;
        RECT 9.090 0.710 9.100 0.944 ;
        RECT 9.100 0.720 9.110 0.954 ;
        RECT 9.110 0.730 9.120 0.964 ;
        RECT 9.120 0.740 9.130 0.974 ;
        RECT 9.130 0.750 9.140 0.984 ;
        RECT 8.945 0.630 8.955 0.800 ;
        RECT 8.955 0.630 8.965 0.810 ;
        RECT 8.965 0.630 8.975 0.820 ;
        RECT 8.975 0.630 8.985 0.830 ;
        RECT 8.985 0.630 8.995 0.840 ;
        RECT 8.995 0.630 9.005 0.850 ;
        RECT 9.005 0.630 9.015 0.860 ;
        RECT 9.015 0.630 9.021 0.870 ;
        RECT 8.115 0.630 8.125 0.864 ;
        RECT 8.125 0.630 8.135 0.854 ;
        RECT 8.135 0.630 8.145 0.844 ;
        RECT 8.145 0.630 8.155 0.834 ;
        RECT 8.155 0.630 8.165 0.824 ;
        RECT 8.165 0.630 8.175 0.814 ;
        RECT 8.175 0.630 8.185 0.804 ;
        RECT 8.185 0.630 8.191 0.800 ;
        RECT 8.025 0.720 8.035 0.954 ;
        RECT 8.035 0.710 8.045 0.944 ;
        RECT 8.045 0.700 8.055 0.934 ;
        RECT 8.055 0.690 8.065 0.924 ;
        RECT 8.065 0.680 8.075 0.914 ;
        RECT 8.075 0.670 8.085 0.904 ;
        RECT 8.085 0.660 8.095 0.894 ;
        RECT 8.095 0.650 8.105 0.884 ;
        RECT 8.105 0.640 8.115 0.874 ;
        RECT 7.950 0.795 7.960 0.965 ;
        RECT 7.960 0.785 7.970 0.965 ;
        RECT 7.970 0.775 7.980 0.965 ;
        RECT 7.980 0.765 7.990 0.965 ;
        RECT 7.990 0.755 8.000 0.965 ;
        RECT 8.000 0.745 8.010 0.965 ;
        RECT 8.010 0.735 8.020 0.965 ;
        RECT 8.020 0.725 8.026 0.965 ;
        RECT 7.520 0.725 7.530 0.965 ;
        RECT 7.530 0.735 7.540 0.965 ;
        RECT 7.540 0.745 7.550 0.965 ;
        RECT 7.550 0.755 7.560 0.965 ;
        RECT 7.560 0.765 7.570 0.965 ;
        RECT 7.570 0.775 7.580 0.965 ;
        RECT 7.580 0.785 7.590 0.965 ;
        RECT 7.590 0.795 7.600 0.965 ;
        RECT 7.375 0.580 7.385 0.820 ;
        RECT 7.385 0.590 7.395 0.830 ;
        RECT 7.395 0.600 7.405 0.840 ;
        RECT 7.405 0.610 7.415 0.850 ;
        RECT 7.415 0.620 7.425 0.860 ;
        RECT 7.425 0.630 7.435 0.870 ;
        RECT 7.435 0.640 7.445 0.880 ;
        RECT 7.445 0.650 7.455 0.890 ;
        RECT 7.455 0.660 7.465 0.900 ;
        RECT 7.465 0.670 7.475 0.910 ;
        RECT 7.475 0.680 7.485 0.920 ;
        RECT 7.485 0.690 7.495 0.930 ;
        RECT 7.495 0.700 7.505 0.940 ;
        RECT 7.505 0.710 7.515 0.950 ;
        RECT 7.515 0.715 7.521 0.959 ;
        RECT 7.295 0.570 7.305 0.740 ;
        RECT 7.305 0.570 7.315 0.750 ;
        RECT 7.315 0.570 7.325 0.760 ;
        RECT 7.325 0.570 7.335 0.770 ;
        RECT 7.335 0.570 7.345 0.780 ;
        RECT 7.345 0.570 7.355 0.790 ;
        RECT 7.355 0.570 7.365 0.800 ;
        RECT 7.365 0.570 7.375 0.810 ;
        RECT 6.635 0.920 6.805 2.565 ;
        RECT 6.570 0.920 6.870 1.090 ;
        RECT 9.545 1.520 9.715 2.565 ;
        RECT 6.635 2.395 9.715 2.565 ;
        RECT 9.545 1.520 9.790 1.820 ;
  END 
END FAHHD1XHT

MACRO FAHDUXHT
  CLASS  CORE ;
  FOREIGN FAHDUXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.070 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.475 1.270 6.870 1.720 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.495 0.520 2.835 ;
    END
  END B
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.710 1.060 10.880 2.835 ;
        RECT 10.710 2.460 10.970 2.835 ;
    END
  END S
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.070 1.680 7.570 2.015 ;
    END
  END CI
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.350 -0.300 0.585 0.660 ;
        RECT 7.395 -0.300 7.695 0.435 ;
        RECT 10.185 -0.300 10.485 0.845 ;
        RECT 0.000 -0.300 11.070 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.490 3.015 0.790 3.990 ;
        RECT 7.875 3.255 8.175 3.990 ;
        RECT 10.250 2.915 10.420 3.990 ;
        RECT 0.000 3.390 11.070 3.990 ;
    END
  END VDD
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.530 0.855 9.840 1.195 ;
        RECT 9.670 0.855 9.840 2.280 ;
    END
  END CO
  OBS 
      LAYER M1 ;
        RECT 1.880 0.495 2.115 1.165 ;
        RECT 1.180 0.910 1.350 2.365 ;
        RECT 1.180 1.825 2.325 1.995 ;
        RECT 3.440 0.910 3.610 2.365 ;
        RECT 3.375 2.165 3.675 2.365 ;
        RECT 3.440 1.585 3.885 1.755 ;
        RECT 3.375 2.165 4.265 2.335 ;
        RECT 2.920 0.910 3.090 2.735 ;
        RECT 1.465 2.565 4.370 2.735 ;
        RECT 0.170 0.910 0.340 2.310 ;
        RECT 0.170 1.585 1.000 1.755 ;
        RECT 0.765 0.480 0.935 2.805 ;
        RECT 0.765 2.635 1.140 2.805 ;
        RECT 0.765 1.520 1.000 1.820 ;
        RECT 0.970 2.635 1.140 3.085 ;
        RECT 0.765 0.480 1.700 0.650 ;
        RECT 1.530 0.480 1.700 1.515 ;
        RECT 1.530 1.345 2.095 1.515 ;
        RECT 4.550 0.860 4.720 3.085 ;
        RECT 0.970 2.915 4.720 3.085 ;
        RECT 6.050 0.900 6.220 2.140 ;
        RECT 6.050 0.900 6.835 1.070 ;
        RECT 6.050 1.970 6.835 2.140 ;
        RECT 7.610 1.325 7.920 1.495 ;
        RECT 5.525 0.920 5.695 2.490 ;
        RECT 5.525 0.920 5.825 1.095 ;
        RECT 5.525 2.165 5.825 2.490 ;
        RECT 5.525 2.320 7.235 2.490 ;
        RECT 7.610 0.965 7.780 1.495 ;
        RECT 7.545 0.965 7.845 1.135 ;
        RECT 7.750 1.325 7.920 2.375 ;
        RECT 7.435 2.205 7.920 2.375 ;
        RECT 7.750 1.600 8.080 1.900 ;
        RECT 7.350 2.205 7.360 2.449 ;
        RECT 7.360 2.205 7.370 2.439 ;
        RECT 7.370 2.205 7.380 2.429 ;
        RECT 7.380 2.205 7.390 2.419 ;
        RECT 7.390 2.205 7.400 2.409 ;
        RECT 7.400 2.205 7.410 2.399 ;
        RECT 7.410 2.205 7.420 2.389 ;
        RECT 7.420 2.205 7.430 2.379 ;
        RECT 7.430 2.205 7.436 2.375 ;
        RECT 7.320 2.235 7.330 2.479 ;
        RECT 7.330 2.225 7.340 2.469 ;
        RECT 7.340 2.215 7.350 2.459 ;
        RECT 7.235 2.320 7.245 2.490 ;
        RECT 7.245 2.310 7.255 2.490 ;
        RECT 7.255 2.300 7.265 2.490 ;
        RECT 7.265 2.290 7.275 2.490 ;
        RECT 7.275 2.280 7.285 2.490 ;
        RECT 7.285 2.270 7.295 2.490 ;
        RECT 7.295 2.260 7.305 2.490 ;
        RECT 7.305 2.250 7.315 2.490 ;
        RECT 7.315 2.240 7.321 2.490 ;
        RECT 5.665 2.670 7.400 2.840 ;
        RECT 8.055 0.965 8.460 1.135 ;
        RECT 8.120 2.100 8.300 2.725 ;
        RECT 7.590 2.555 8.300 2.725 ;
        RECT 8.290 0.965 8.460 2.335 ;
        RECT 8.120 2.100 8.460 2.335 ;
        RECT 7.515 2.555 7.525 2.789 ;
        RECT 7.525 2.555 7.535 2.779 ;
        RECT 7.535 2.555 7.545 2.769 ;
        RECT 7.545 2.555 7.555 2.759 ;
        RECT 7.555 2.555 7.565 2.749 ;
        RECT 7.565 2.555 7.575 2.739 ;
        RECT 7.575 2.555 7.585 2.729 ;
        RECT 7.585 2.555 7.591 2.725 ;
        RECT 7.475 2.595 7.485 2.829 ;
        RECT 7.485 2.585 7.495 2.819 ;
        RECT 7.495 2.575 7.505 2.809 ;
        RECT 7.505 2.565 7.515 2.799 ;
        RECT 7.400 2.670 7.410 2.840 ;
        RECT 7.410 2.660 7.420 2.840 ;
        RECT 7.420 2.650 7.430 2.840 ;
        RECT 7.430 2.640 7.440 2.840 ;
        RECT 7.440 2.630 7.450 2.840 ;
        RECT 7.450 2.620 7.460 2.840 ;
        RECT 7.460 2.610 7.470 2.840 ;
        RECT 7.470 2.600 7.476 2.840 ;
        RECT 2.560 0.500 2.740 1.145 ;
        RECT 2.335 0.975 2.740 1.145 ;
        RECT 2.570 0.500 2.740 2.365 ;
        RECT 1.655 2.195 2.740 2.365 ;
        RECT 4.030 0.500 4.200 1.160 ;
        RECT 7.045 0.500 7.215 0.785 ;
        RECT 2.560 0.500 7.215 0.670 ;
        RECT 7.885 0.520 8.055 0.785 ;
        RECT 7.045 0.615 8.055 0.785 ;
        RECT 7.885 0.520 9.330 0.690 ;
        RECT 9.160 0.520 9.330 2.335 ;
        RECT 9.095 2.165 9.395 2.335 ;
        RECT 5.070 0.860 5.240 3.190 ;
        RECT 5.070 3.020 7.560 3.190 ;
        RECT 7.760 2.905 10.070 3.075 ;
        RECT 7.675 2.905 7.685 3.149 ;
        RECT 7.685 2.905 7.695 3.139 ;
        RECT 7.695 2.905 7.705 3.129 ;
        RECT 7.705 2.905 7.715 3.119 ;
        RECT 7.715 2.905 7.725 3.109 ;
        RECT 7.725 2.905 7.735 3.099 ;
        RECT 7.735 2.905 7.745 3.089 ;
        RECT 7.745 2.905 7.755 3.079 ;
        RECT 7.755 2.905 7.761 3.075 ;
        RECT 7.645 2.935 7.655 3.179 ;
        RECT 7.655 2.925 7.665 3.169 ;
        RECT 7.665 2.915 7.675 3.159 ;
        RECT 7.560 3.020 7.570 3.190 ;
        RECT 7.570 3.010 7.580 3.190 ;
        RECT 7.580 3.000 7.590 3.190 ;
        RECT 7.590 2.990 7.600 3.190 ;
        RECT 7.600 2.980 7.610 3.190 ;
        RECT 7.610 2.970 7.620 3.190 ;
        RECT 7.620 2.960 7.630 3.190 ;
        RECT 7.630 2.950 7.640 3.190 ;
        RECT 7.640 2.940 7.646 3.190 ;
        RECT 8.640 0.900 8.810 2.685 ;
        RECT 10.115 1.530 10.285 2.685 ;
        RECT 8.640 2.515 10.285 2.685 ;
        RECT 10.115 1.530 10.530 1.830 ;
  END 
END FAHDUXHT

MACRO FAHDMXHT
  CLASS  CORE ;
  FOREIGN FAHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.590 1.125 4.010 1.795 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 1.550 0.925 1.970 ;
    END
  END B
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.275 1.060 10.445 2.830 ;
        RECT 10.275 2.500 10.560 2.830 ;
    END
  END S
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.885 2.125 7.340 2.560 ;
    END
  END CI
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.075 ;
        RECT 1.175 -0.300 1.475 0.920 ;
        RECT 3.570 -0.300 3.870 0.460 ;
        RECT 7.375 -0.300 7.675 0.435 ;
        RECT 9.690 -0.300 9.990 1.295 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.465 0.405 3.990 ;
        RECT 1.135 3.070 1.435 3.990 ;
        RECT 3.585 3.025 3.885 3.990 ;
        RECT 6.930 3.090 7.230 3.990 ;
        RECT 9.660 2.810 9.960 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.120 0.860 9.330 2.280 ;
        RECT 9.120 0.860 9.405 1.360 ;
    END
  END CO
  OBS 
      LAYER M1 ;
        RECT 1.795 1.035 1.965 2.540 ;
        RECT 1.750 2.135 1.965 2.540 ;
        RECT 1.750 2.370 2.490 2.540 ;
        RECT 2.320 2.370 2.490 2.860 ;
        RECT 2.320 2.690 2.790 2.860 ;
        RECT 3.085 0.990 3.255 2.145 ;
        RECT 4.200 0.990 4.370 1.530 ;
        RECT 4.265 1.360 4.435 2.145 ;
        RECT 3.035 1.975 4.435 2.145 ;
        RECT 4.200 1.360 5.060 1.530 ;
        RECT 4.890 1.360 5.060 1.660 ;
        RECT 0.625 1.100 1.570 1.270 ;
        RECT 0.625 2.290 1.570 2.460 ;
        RECT 1.400 1.100 1.570 2.890 ;
        RECT 1.400 1.515 1.615 1.815 ;
        RECT 1.400 2.720 2.140 2.890 ;
        RECT 1.970 2.720 2.140 3.210 ;
        RECT 1.970 3.040 2.875 3.210 ;
        RECT 3.140 2.675 4.360 2.845 ;
        RECT 4.190 2.675 4.360 3.085 ;
        RECT 5.270 2.190 5.440 3.085 ;
        RECT 4.190 2.915 5.440 3.085 ;
        RECT 5.270 2.190 5.545 2.360 ;
        RECT 5.590 1.245 5.760 1.415 ;
        RECT 5.760 1.245 5.770 2.209 ;
        RECT 5.770 1.245 5.780 2.199 ;
        RECT 5.780 1.245 5.790 2.189 ;
        RECT 5.790 1.245 5.800 2.179 ;
        RECT 5.800 1.245 5.810 2.169 ;
        RECT 5.810 1.245 5.820 2.159 ;
        RECT 5.820 1.245 5.830 2.149 ;
        RECT 5.830 1.245 5.840 2.139 ;
        RECT 5.840 1.245 5.850 2.129 ;
        RECT 5.850 1.245 5.860 2.119 ;
        RECT 5.860 1.245 5.870 2.109 ;
        RECT 5.870 1.245 5.880 2.099 ;
        RECT 5.880 1.245 5.890 2.089 ;
        RECT 5.890 1.245 5.900 2.079 ;
        RECT 5.900 1.245 5.910 2.069 ;
        RECT 5.910 1.245 5.920 2.059 ;
        RECT 5.920 1.245 5.930 2.049 ;
        RECT 5.620 2.115 5.630 2.349 ;
        RECT 5.630 2.105 5.640 2.339 ;
        RECT 5.640 2.095 5.650 2.329 ;
        RECT 5.650 2.085 5.660 2.319 ;
        RECT 5.660 2.075 5.670 2.309 ;
        RECT 5.670 2.065 5.680 2.299 ;
        RECT 5.680 2.055 5.690 2.289 ;
        RECT 5.690 2.045 5.700 2.279 ;
        RECT 5.700 2.035 5.710 2.269 ;
        RECT 5.710 2.025 5.720 2.259 ;
        RECT 5.720 2.015 5.730 2.249 ;
        RECT 5.730 2.005 5.740 2.239 ;
        RECT 5.740 1.995 5.750 2.229 ;
        RECT 5.750 1.985 5.760 2.219 ;
        RECT 5.545 2.190 5.555 2.360 ;
        RECT 5.555 2.180 5.565 2.360 ;
        RECT 5.565 2.170 5.575 2.360 ;
        RECT 5.575 2.160 5.585 2.360 ;
        RECT 5.585 2.150 5.595 2.360 ;
        RECT 5.595 2.140 5.605 2.360 ;
        RECT 5.605 2.130 5.615 2.360 ;
        RECT 5.615 2.120 5.621 2.360 ;
        RECT 2.970 2.675 2.980 3.179 ;
        RECT 2.980 2.675 2.990 3.169 ;
        RECT 2.990 2.675 3.000 3.159 ;
        RECT 3.000 2.675 3.010 3.149 ;
        RECT 3.010 2.675 3.020 3.139 ;
        RECT 3.020 2.675 3.030 3.129 ;
        RECT 3.030 2.675 3.040 3.119 ;
        RECT 3.040 2.675 3.050 3.109 ;
        RECT 3.050 2.675 3.060 3.099 ;
        RECT 3.060 2.675 3.070 3.089 ;
        RECT 3.070 2.675 3.080 3.079 ;
        RECT 3.080 2.675 3.090 3.069 ;
        RECT 3.090 2.675 3.100 3.059 ;
        RECT 3.100 2.675 3.110 3.049 ;
        RECT 3.110 2.675 3.120 3.039 ;
        RECT 3.120 2.675 3.130 3.029 ;
        RECT 3.130 2.675 3.140 3.019 ;
        RECT 2.950 2.965 2.960 3.199 ;
        RECT 2.960 2.955 2.970 3.189 ;
        RECT 2.875 3.040 2.885 3.210 ;
        RECT 2.885 3.030 2.895 3.210 ;
        RECT 2.895 3.020 2.905 3.210 ;
        RECT 2.905 3.010 2.915 3.210 ;
        RECT 2.915 3.000 2.925 3.210 ;
        RECT 2.925 2.990 2.935 3.210 ;
        RECT 2.935 2.980 2.945 3.210 ;
        RECT 2.945 2.970 2.951 3.210 ;
        RECT 6.705 1.245 6.800 1.935 ;
        RECT 6.705 1.245 6.930 1.415 ;
        RECT 6.705 1.765 7.620 1.935 ;
        RECT 6.630 1.245 6.640 2.395 ;
        RECT 6.640 1.245 6.650 2.385 ;
        RECT 6.650 1.245 6.660 2.375 ;
        RECT 6.660 1.245 6.670 2.365 ;
        RECT 6.670 1.245 6.680 2.355 ;
        RECT 6.680 1.245 6.690 2.345 ;
        RECT 6.690 1.245 6.700 2.335 ;
        RECT 6.700 1.245 6.706 2.329 ;
        RECT 6.535 1.765 6.545 2.489 ;
        RECT 6.545 1.765 6.555 2.479 ;
        RECT 6.555 1.765 6.565 2.469 ;
        RECT 6.565 1.765 6.575 2.459 ;
        RECT 6.575 1.765 6.585 2.449 ;
        RECT 6.585 1.765 6.595 2.439 ;
        RECT 6.595 1.765 6.605 2.429 ;
        RECT 6.605 1.765 6.615 2.419 ;
        RECT 6.615 1.765 6.625 2.409 ;
        RECT 6.625 1.765 6.631 2.405 ;
        RECT 6.480 2.310 6.490 2.544 ;
        RECT 6.490 2.300 6.500 2.534 ;
        RECT 6.500 2.290 6.510 2.524 ;
        RECT 6.510 2.280 6.520 2.514 ;
        RECT 6.520 2.270 6.530 2.504 ;
        RECT 6.530 2.260 6.536 2.500 ;
        RECT 6.310 2.480 6.320 2.780 ;
        RECT 6.320 2.470 6.330 2.780 ;
        RECT 6.330 2.460 6.340 2.780 ;
        RECT 6.340 2.450 6.350 2.780 ;
        RECT 6.350 2.440 6.360 2.780 ;
        RECT 6.360 2.430 6.370 2.780 ;
        RECT 6.370 2.420 6.380 2.780 ;
        RECT 6.380 2.410 6.390 2.780 ;
        RECT 6.390 2.400 6.400 2.780 ;
        RECT 6.400 2.390 6.410 2.780 ;
        RECT 6.410 2.380 6.420 2.780 ;
        RECT 6.420 2.370 6.430 2.780 ;
        RECT 6.430 2.360 6.440 2.780 ;
        RECT 6.440 2.350 6.450 2.780 ;
        RECT 6.450 2.340 6.460 2.780 ;
        RECT 6.460 2.330 6.470 2.780 ;
        RECT 6.470 2.320 6.480 2.780 ;
        RECT 2.560 1.470 2.855 1.640 ;
        RECT 2.560 0.990 2.730 1.640 ;
        RECT 2.685 1.470 2.855 2.495 ;
        RECT 4.750 1.840 4.920 2.495 ;
        RECT 2.685 2.325 4.920 2.495 ;
        RECT 5.240 0.875 5.410 2.010 ;
        RECT 4.750 1.840 5.410 2.010 ;
        RECT 5.240 1.600 5.580 1.900 ;
        RECT 5.240 0.875 6.985 1.045 ;
        RECT 7.585 2.115 7.755 2.500 ;
        RECT 7.255 1.070 7.970 1.240 ;
        RECT 7.800 1.070 7.970 2.285 ;
        RECT 7.585 2.115 7.970 2.285 ;
        RECT 7.180 1.005 7.190 1.239 ;
        RECT 7.190 1.015 7.200 1.239 ;
        RECT 7.200 1.025 7.210 1.239 ;
        RECT 7.210 1.035 7.220 1.239 ;
        RECT 7.220 1.045 7.230 1.239 ;
        RECT 7.230 1.055 7.240 1.239 ;
        RECT 7.240 1.065 7.250 1.239 ;
        RECT 7.250 1.070 7.256 1.240 ;
        RECT 7.060 0.885 7.070 1.119 ;
        RECT 7.070 0.895 7.080 1.129 ;
        RECT 7.080 0.905 7.090 1.139 ;
        RECT 7.090 0.915 7.100 1.149 ;
        RECT 7.100 0.925 7.110 1.159 ;
        RECT 7.110 0.935 7.120 1.169 ;
        RECT 7.120 0.945 7.130 1.179 ;
        RECT 7.130 0.955 7.140 1.189 ;
        RECT 7.140 0.965 7.150 1.199 ;
        RECT 7.150 0.975 7.160 1.209 ;
        RECT 7.160 0.985 7.170 1.219 ;
        RECT 7.170 0.995 7.180 1.229 ;
        RECT 6.985 0.875 6.995 1.045 ;
        RECT 6.995 0.875 7.005 1.055 ;
        RECT 7.005 0.875 7.015 1.065 ;
        RECT 7.015 0.875 7.025 1.075 ;
        RECT 7.025 0.875 7.035 1.085 ;
        RECT 7.035 0.875 7.045 1.095 ;
        RECT 7.045 0.875 7.055 1.105 ;
        RECT 7.055 0.875 7.061 1.115 ;
        RECT 2.205 0.640 2.375 2.190 ;
        RECT 2.205 2.020 2.505 2.190 ;
        RECT 2.205 0.640 4.890 0.810 ;
        RECT 4.720 0.525 4.890 1.170 ;
        RECT 4.720 0.525 7.135 0.695 ;
        RECT 7.345 0.660 8.895 0.830 ;
        RECT 8.725 0.660 8.895 2.435 ;
        RECT 8.560 2.265 8.895 2.435 ;
        RECT 7.270 0.595 7.280 0.829 ;
        RECT 7.280 0.605 7.290 0.829 ;
        RECT 7.290 0.615 7.300 0.829 ;
        RECT 7.300 0.625 7.310 0.829 ;
        RECT 7.310 0.635 7.320 0.829 ;
        RECT 7.320 0.645 7.330 0.829 ;
        RECT 7.330 0.655 7.340 0.829 ;
        RECT 7.340 0.660 7.346 0.830 ;
        RECT 7.210 0.535 7.220 0.769 ;
        RECT 7.220 0.545 7.230 0.779 ;
        RECT 7.230 0.555 7.240 0.789 ;
        RECT 7.240 0.565 7.250 0.799 ;
        RECT 7.250 0.575 7.260 0.809 ;
        RECT 7.260 0.585 7.270 0.819 ;
        RECT 7.135 0.525 7.145 0.695 ;
        RECT 7.145 0.525 7.155 0.705 ;
        RECT 7.155 0.525 7.165 0.715 ;
        RECT 7.165 0.525 7.175 0.725 ;
        RECT 7.175 0.525 7.185 0.735 ;
        RECT 7.185 0.525 7.195 0.745 ;
        RECT 7.195 0.525 7.205 0.755 ;
        RECT 7.205 0.525 7.211 0.765 ;
        RECT 5.725 2.545 5.960 2.715 ;
        RECT 6.110 1.245 6.175 1.415 ;
        RECT 6.345 1.245 6.410 1.415 ;
        RECT 6.130 2.960 6.555 3.130 ;
        RECT 6.850 2.740 7.860 2.910 ;
        RECT 7.690 2.740 7.860 3.135 ;
        RECT 7.690 2.965 9.480 3.135 ;
        RECT 6.775 2.740 6.785 2.974 ;
        RECT 6.785 2.740 6.795 2.964 ;
        RECT 6.795 2.740 6.805 2.954 ;
        RECT 6.805 2.740 6.815 2.944 ;
        RECT 6.815 2.740 6.825 2.934 ;
        RECT 6.825 2.740 6.835 2.924 ;
        RECT 6.835 2.740 6.845 2.914 ;
        RECT 6.845 2.740 6.851 2.910 ;
        RECT 6.630 2.885 6.640 3.119 ;
        RECT 6.640 2.875 6.650 3.109 ;
        RECT 6.650 2.865 6.660 3.099 ;
        RECT 6.660 2.855 6.670 3.089 ;
        RECT 6.670 2.845 6.680 3.079 ;
        RECT 6.680 2.835 6.690 3.069 ;
        RECT 6.690 2.825 6.700 3.059 ;
        RECT 6.700 2.815 6.710 3.049 ;
        RECT 6.710 2.805 6.720 3.039 ;
        RECT 6.720 2.795 6.730 3.029 ;
        RECT 6.730 2.785 6.740 3.019 ;
        RECT 6.740 2.775 6.750 3.009 ;
        RECT 6.750 2.765 6.760 2.999 ;
        RECT 6.760 2.755 6.770 2.989 ;
        RECT 6.770 2.745 6.776 2.985 ;
        RECT 6.555 2.960 6.565 3.130 ;
        RECT 6.565 2.950 6.575 3.130 ;
        RECT 6.575 2.940 6.585 3.130 ;
        RECT 6.585 2.930 6.595 3.130 ;
        RECT 6.595 2.920 6.605 3.130 ;
        RECT 6.605 2.910 6.615 3.130 ;
        RECT 6.615 2.900 6.625 3.130 ;
        RECT 6.625 2.890 6.631 3.130 ;
        RECT 6.175 1.245 6.185 2.325 ;
        RECT 6.185 1.245 6.195 2.315 ;
        RECT 6.195 1.245 6.205 2.305 ;
        RECT 6.205 1.245 6.215 2.295 ;
        RECT 6.215 1.245 6.225 2.285 ;
        RECT 6.225 1.245 6.235 2.275 ;
        RECT 6.235 1.245 6.245 2.265 ;
        RECT 6.245 1.245 6.255 2.255 ;
        RECT 6.255 1.245 6.265 2.245 ;
        RECT 6.265 1.245 6.275 2.235 ;
        RECT 6.275 1.245 6.285 2.225 ;
        RECT 6.285 1.245 6.295 2.215 ;
        RECT 6.295 1.245 6.305 2.205 ;
        RECT 6.305 1.245 6.315 2.195 ;
        RECT 6.315 1.245 6.325 2.185 ;
        RECT 6.325 1.245 6.335 2.175 ;
        RECT 6.335 1.245 6.345 2.165 ;
        RECT 6.130 2.135 6.140 2.369 ;
        RECT 6.140 2.125 6.150 2.359 ;
        RECT 6.150 2.115 6.160 2.349 ;
        RECT 6.160 2.105 6.170 2.339 ;
        RECT 6.170 2.095 6.176 2.335 ;
        RECT 5.960 2.305 5.970 3.129 ;
        RECT 5.970 2.295 5.980 3.129 ;
        RECT 5.980 2.285 5.990 3.129 ;
        RECT 5.990 2.275 6.000 3.129 ;
        RECT 6.000 2.265 6.010 3.129 ;
        RECT 6.010 2.255 6.020 3.129 ;
        RECT 6.020 2.245 6.030 3.129 ;
        RECT 6.030 2.235 6.040 3.129 ;
        RECT 6.040 2.225 6.050 3.129 ;
        RECT 6.050 2.215 6.060 3.129 ;
        RECT 6.060 2.205 6.070 3.129 ;
        RECT 6.070 2.195 6.080 3.129 ;
        RECT 6.080 2.185 6.090 3.129 ;
        RECT 6.090 2.175 6.100 3.129 ;
        RECT 6.100 2.165 6.110 3.129 ;
        RECT 6.110 2.155 6.120 3.129 ;
        RECT 6.120 2.145 6.130 3.129 ;
        RECT 8.205 1.010 8.375 2.785 ;
        RECT 8.040 2.465 8.375 2.785 ;
        RECT 9.135 2.460 9.305 2.785 ;
        RECT 8.040 2.615 9.305 2.785 ;
        RECT 9.135 2.460 10.095 2.630 ;
        RECT 9.925 1.545 10.095 2.630 ;
  END 
END FAHDMXHT

MACRO DEL4HDMXHT
  CLASS  CORE ;
  FOREIGN DEL4HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 2.470 0.510 2.890 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 2.765 -0.300 3.065 0.785 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.350 0.700 3.520 2.580 ;
        RECT 3.350 1.250 3.590 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.100 0.860 3.990 ;
        RECT 2.765 2.675 3.065 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.605 1.390 1.775 ;
        RECT 1.630 1.060 1.800 2.280 ;
        RECT 1.630 1.605 2.465 1.775 ;
        RECT 1.825 0.615 2.370 0.785 ;
        RECT 2.200 0.615 2.370 1.265 ;
        RECT 2.290 2.160 2.460 2.845 ;
        RECT 1.820 2.675 2.460 2.845 ;
        RECT 2.200 1.095 3.170 1.265 ;
        RECT 3.000 1.095 3.170 2.330 ;
        RECT 2.290 2.160 3.170 2.330 ;
  END 
END DEL4HDMXHT

MACRO FFDNSRHDLXHT
  CLASS  CORE ;
  FOREIGN FFDNSRHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.890 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN CKN
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.605 0.550 2.060 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.540 1.060 11.715 2.430 ;
        RECT 11.540 2.070 11.790 2.430 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.440 1.125 10.970 1.295 ;
        RECT 10.760 1.125 10.970 2.280 ;
        RECT 10.440 1.980 10.970 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.655 1.330 2.050 1.785 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.380 1.580 3.850 2.035 ;
    END
  END RN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.855 ;
        RECT 1.655 -0.300 1.955 0.730 ;
        RECT 3.435 -0.300 3.735 1.160 ;
        RECT 6.175 -0.300 6.475 0.730 ;
        RECT 8.005 -0.300 8.305 0.730 ;
        RECT 10.050 -0.300 10.350 0.785 ;
        RECT 11.020 -0.300 11.320 0.745 ;
        RECT 0.000 -0.300 11.890 0.300 ;
    END
  END GND
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 9.530 1.635 9.910 2.020 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.785 2.810 1.765 3.990 ;
        RECT 3.600 3.025 4.580 3.990 ;
        RECT 6.160 3.025 6.460 3.990 ;
        RECT 8.130 2.365 8.430 3.990 ;
        RECT 9.875 2.945 10.175 3.990 ;
        RECT 10.925 2.945 11.225 3.990 ;
        RECT 0.000 3.390 11.890 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.210 0.980 1.380 2.280 ;
        RECT 2.135 0.620 2.305 1.150 ;
        RECT 1.210 0.980 2.305 1.150 ;
        RECT 2.135 0.620 3.135 0.790 ;
        RECT 2.965 0.620 3.135 2.085 ;
        RECT 2.775 1.915 3.135 2.085 ;
        RECT 4.020 0.925 4.220 1.225 ;
        RECT 4.050 0.925 4.220 2.145 ;
        RECT 4.050 1.470 4.845 1.770 ;
        RECT 2.425 1.565 2.595 2.495 ;
        RECT 2.485 0.990 2.655 1.735 ;
        RECT 2.425 1.565 2.655 1.735 ;
        RECT 2.485 0.990 2.785 1.160 ;
        RECT 2.425 2.295 2.815 2.495 ;
        RECT 4.400 1.950 4.570 2.495 ;
        RECT 2.425 2.325 4.570 2.495 ;
        RECT 5.025 1.550 5.195 2.120 ;
        RECT 4.400 1.950 5.195 2.120 ;
        RECT 5.025 1.550 5.360 1.850 ;
        RECT 4.465 0.990 4.765 1.230 ;
        RECT 4.465 1.060 5.740 1.230 ;
        RECT 5.570 1.060 5.740 1.360 ;
        RECT 5.045 0.560 5.345 0.825 ;
        RECT 4.095 0.560 5.665 0.730 ;
        RECT 5.540 1.590 5.710 2.215 ;
        RECT 5.410 2.045 5.710 2.215 ;
        RECT 5.540 1.590 5.920 1.760 ;
        RECT 6.090 1.590 6.495 1.760 ;
        RECT 5.920 0.740 5.930 1.760 ;
        RECT 5.930 0.750 5.940 1.760 ;
        RECT 5.940 0.760 5.950 1.760 ;
        RECT 5.950 0.770 5.960 1.760 ;
        RECT 5.960 0.780 5.970 1.760 ;
        RECT 5.970 0.790 5.980 1.760 ;
        RECT 5.980 0.800 5.990 1.760 ;
        RECT 5.990 0.810 6.000 1.760 ;
        RECT 6.000 0.820 6.010 1.760 ;
        RECT 6.010 0.830 6.020 1.760 ;
        RECT 6.020 0.840 6.030 1.760 ;
        RECT 6.030 0.850 6.040 1.760 ;
        RECT 6.040 0.860 6.050 1.760 ;
        RECT 6.050 0.870 6.060 1.760 ;
        RECT 6.060 0.880 6.070 1.760 ;
        RECT 6.070 0.890 6.080 1.760 ;
        RECT 6.080 0.900 6.090 1.760 ;
        RECT 5.750 0.570 5.760 0.814 ;
        RECT 5.760 0.580 5.770 0.824 ;
        RECT 5.770 0.590 5.780 0.834 ;
        RECT 5.780 0.600 5.790 0.844 ;
        RECT 5.790 0.610 5.800 0.854 ;
        RECT 5.800 0.620 5.810 0.864 ;
        RECT 5.810 0.630 5.820 0.874 ;
        RECT 5.820 0.640 5.830 0.884 ;
        RECT 5.830 0.650 5.840 0.894 ;
        RECT 5.840 0.660 5.850 0.904 ;
        RECT 5.850 0.670 5.860 0.914 ;
        RECT 5.860 0.680 5.870 0.924 ;
        RECT 5.870 0.690 5.880 0.934 ;
        RECT 5.880 0.700 5.890 0.944 ;
        RECT 5.890 0.710 5.900 0.954 ;
        RECT 5.900 0.720 5.910 0.964 ;
        RECT 5.910 0.730 5.920 0.974 ;
        RECT 5.665 0.560 5.675 0.730 ;
        RECT 5.675 0.560 5.685 0.740 ;
        RECT 5.685 0.560 5.695 0.750 ;
        RECT 5.695 0.560 5.705 0.760 ;
        RECT 5.705 0.560 5.715 0.770 ;
        RECT 5.715 0.560 5.725 0.780 ;
        RECT 5.725 0.560 5.735 0.790 ;
        RECT 5.735 0.560 5.745 0.800 ;
        RECT 5.745 0.560 5.751 0.810 ;
        RECT 0.105 1.125 1.030 1.295 ;
        RECT 0.105 2.245 1.030 2.415 ;
        RECT 0.860 1.125 1.030 2.630 ;
        RECT 0.860 2.460 2.170 2.630 ;
        RECT 2.000 2.460 2.170 2.845 ;
        RECT 4.750 2.395 4.920 2.845 ;
        RECT 2.000 2.675 4.920 2.845 ;
        RECT 4.750 2.395 5.785 2.565 ;
        RECT 5.960 2.295 6.700 2.465 ;
        RECT 6.875 2.395 7.385 2.565 ;
        RECT 7.215 2.395 7.385 2.695 ;
        RECT 6.800 2.330 6.810 2.564 ;
        RECT 6.810 2.340 6.820 2.564 ;
        RECT 6.820 2.350 6.830 2.564 ;
        RECT 6.830 2.360 6.840 2.564 ;
        RECT 6.840 2.370 6.850 2.564 ;
        RECT 6.850 2.380 6.860 2.564 ;
        RECT 6.860 2.390 6.870 2.564 ;
        RECT 6.870 2.395 6.876 2.565 ;
        RECT 6.775 2.305 6.785 2.539 ;
        RECT 6.785 2.315 6.795 2.549 ;
        RECT 6.795 2.320 6.801 2.560 ;
        RECT 6.700 2.295 6.710 2.465 ;
        RECT 6.710 2.295 6.720 2.475 ;
        RECT 6.720 2.295 6.730 2.485 ;
        RECT 6.730 2.295 6.740 2.495 ;
        RECT 6.740 2.295 6.750 2.505 ;
        RECT 6.750 2.295 6.760 2.515 ;
        RECT 6.760 2.295 6.770 2.525 ;
        RECT 6.770 2.295 6.776 2.535 ;
        RECT 5.885 2.295 5.895 2.529 ;
        RECT 5.895 2.295 5.905 2.519 ;
        RECT 5.905 2.295 5.915 2.509 ;
        RECT 5.915 2.295 5.925 2.499 ;
        RECT 5.925 2.295 5.935 2.489 ;
        RECT 5.935 2.295 5.945 2.479 ;
        RECT 5.945 2.295 5.955 2.469 ;
        RECT 5.955 2.295 5.961 2.465 ;
        RECT 5.860 2.320 5.870 2.554 ;
        RECT 5.870 2.310 5.880 2.544 ;
        RECT 5.880 2.300 5.886 2.540 ;
        RECT 5.785 2.395 5.795 2.565 ;
        RECT 5.795 2.385 5.805 2.565 ;
        RECT 5.805 2.375 5.815 2.565 ;
        RECT 5.815 2.365 5.825 2.565 ;
        RECT 5.825 2.355 5.835 2.565 ;
        RECT 5.835 2.345 5.845 2.565 ;
        RECT 5.845 2.335 5.855 2.565 ;
        RECT 5.855 2.325 5.861 2.565 ;
        RECT 5.100 2.795 5.270 3.210 ;
        RECT 4.765 3.040 5.270 3.210 ;
        RECT 5.100 2.795 5.890 2.965 ;
        RECT 6.115 2.645 6.510 2.815 ;
        RECT 6.610 2.645 6.625 2.915 ;
        RECT 6.725 2.745 6.950 2.915 ;
        RECT 6.780 2.745 6.950 3.120 ;
        RECT 7.380 1.230 7.735 1.530 ;
        RECT 7.565 1.230 7.735 3.120 ;
        RECT 6.780 2.950 7.735 3.120 ;
        RECT 6.625 2.655 6.635 2.915 ;
        RECT 6.635 2.665 6.645 2.915 ;
        RECT 6.645 2.675 6.655 2.915 ;
        RECT 6.655 2.685 6.665 2.915 ;
        RECT 6.665 2.695 6.675 2.915 ;
        RECT 6.675 2.705 6.685 2.915 ;
        RECT 6.685 2.715 6.695 2.915 ;
        RECT 6.695 2.725 6.705 2.915 ;
        RECT 6.705 2.735 6.715 2.915 ;
        RECT 6.715 2.745 6.725 2.915 ;
        RECT 6.510 2.645 6.520 2.815 ;
        RECT 6.520 2.645 6.530 2.825 ;
        RECT 6.530 2.645 6.540 2.835 ;
        RECT 6.540 2.645 6.550 2.845 ;
        RECT 6.550 2.645 6.560 2.855 ;
        RECT 6.560 2.645 6.570 2.865 ;
        RECT 6.570 2.645 6.580 2.875 ;
        RECT 6.580 2.645 6.590 2.885 ;
        RECT 6.590 2.645 6.600 2.895 ;
        RECT 6.600 2.645 6.610 2.905 ;
        RECT 6.040 2.645 6.050 2.879 ;
        RECT 6.050 2.645 6.060 2.869 ;
        RECT 6.060 2.645 6.070 2.859 ;
        RECT 6.070 2.645 6.080 2.849 ;
        RECT 6.080 2.645 6.090 2.839 ;
        RECT 6.090 2.645 6.100 2.829 ;
        RECT 6.100 2.645 6.110 2.819 ;
        RECT 6.110 2.645 6.116 2.815 ;
        RECT 5.965 2.720 5.975 2.954 ;
        RECT 5.975 2.710 5.985 2.944 ;
        RECT 5.985 2.700 5.995 2.934 ;
        RECT 5.995 2.690 6.005 2.924 ;
        RECT 6.005 2.680 6.015 2.914 ;
        RECT 6.015 2.670 6.025 2.904 ;
        RECT 6.025 2.660 6.035 2.894 ;
        RECT 6.035 2.650 6.041 2.890 ;
        RECT 5.890 2.795 5.900 2.965 ;
        RECT 5.900 2.785 5.910 2.965 ;
        RECT 5.910 2.775 5.920 2.965 ;
        RECT 5.920 2.765 5.930 2.965 ;
        RECT 5.930 2.755 5.940 2.965 ;
        RECT 5.940 2.745 5.950 2.965 ;
        RECT 5.950 2.735 5.960 2.965 ;
        RECT 5.960 2.725 5.966 2.965 ;
        RECT 8.570 0.775 8.740 1.295 ;
        RECT 8.430 1.125 8.740 1.295 ;
        RECT 9.470 0.655 9.770 0.945 ;
        RECT 8.570 0.775 9.770 0.945 ;
        RECT 8.265 1.495 8.435 1.795 ;
        RECT 9.010 1.125 9.310 1.295 ;
        RECT 8.265 1.625 9.310 1.795 ;
        RECT 9.135 1.125 9.310 2.415 ;
        RECT 10.090 1.480 10.260 2.415 ;
        RECT 9.135 2.245 10.260 2.415 ;
        RECT 10.090 1.480 10.580 1.780 ;
        RECT 6.980 0.880 7.150 2.215 ;
        RECT 6.955 2.045 7.255 2.215 ;
        RECT 6.980 0.880 7.810 1.050 ;
        RECT 8.085 1.975 8.945 2.145 ;
        RECT 8.775 1.975 8.945 2.765 ;
        RECT 9.085 2.595 9.385 2.905 ;
        RECT 11.190 1.530 11.360 2.765 ;
        RECT 8.775 2.595 11.360 2.765 ;
        RECT 7.915 0.910 7.925 2.144 ;
        RECT 7.925 0.920 7.935 2.144 ;
        RECT 7.935 0.930 7.945 2.144 ;
        RECT 7.945 0.940 7.955 2.144 ;
        RECT 7.955 0.950 7.965 2.144 ;
        RECT 7.965 0.960 7.975 2.144 ;
        RECT 7.975 0.970 7.985 2.144 ;
        RECT 7.985 0.980 7.995 2.144 ;
        RECT 7.995 0.990 8.005 2.144 ;
        RECT 8.005 1.000 8.015 2.144 ;
        RECT 8.015 1.010 8.025 2.144 ;
        RECT 8.025 1.020 8.035 2.144 ;
        RECT 8.035 1.030 8.045 2.144 ;
        RECT 8.045 1.040 8.055 2.144 ;
        RECT 8.055 1.050 8.065 2.144 ;
        RECT 8.065 1.060 8.075 2.144 ;
        RECT 8.075 1.070 8.085 2.144 ;
        RECT 7.895 0.890 7.905 1.134 ;
        RECT 7.905 0.900 7.915 1.144 ;
        RECT 7.810 0.880 7.820 1.050 ;
        RECT 7.820 0.880 7.830 1.060 ;
        RECT 7.830 0.880 7.840 1.070 ;
        RECT 7.840 0.880 7.850 1.080 ;
        RECT 7.850 0.880 7.860 1.090 ;
        RECT 7.860 0.880 7.870 1.100 ;
        RECT 7.870 0.880 7.880 1.110 ;
        RECT 7.880 0.880 7.890 1.120 ;
        RECT 7.890 0.880 7.896 1.130 ;
  END 
END FFDNSRHDLXHT

MACRO FAHD1XHT
  CLASS  CORE ;
  FOREIGN FAHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.590 1.125 4.010 1.795 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 1.550 0.925 1.970 ;
    END
  END B
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 10.185 0.720 10.355 2.960 ;
        RECT 10.185 2.500 10.560 2.960 ;
    END
  END S
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.885 2.125 7.340 2.560 ;
    END
  END CI
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.075 ;
        RECT 1.175 -0.300 1.475 0.920 ;
        RECT 3.570 -0.300 3.870 0.460 ;
        RECT 7.375 -0.300 7.675 0.435 ;
        RECT 9.600 -0.300 9.900 1.055 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.465 0.405 3.990 ;
        RECT 1.135 3.070 1.435 3.990 ;
        RECT 3.585 3.025 3.885 3.990 ;
        RECT 6.930 3.090 7.230 3.990 ;
        RECT 9.600 2.975 9.900 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 9.120 0.480 9.330 2.280 ;
    END
  END CO
  OBS 
      LAYER M1 ;
        RECT 1.795 1.035 1.965 2.540 ;
        RECT 1.750 2.135 1.965 2.540 ;
        RECT 1.750 2.370 2.490 2.540 ;
        RECT 2.320 2.370 2.490 2.860 ;
        RECT 2.320 2.690 2.790 2.860 ;
        RECT 3.085 0.990 3.255 2.145 ;
        RECT 4.200 0.990 4.370 1.530 ;
        RECT 4.265 1.360 4.435 2.145 ;
        RECT 3.035 1.975 4.435 2.145 ;
        RECT 4.200 1.360 5.060 1.530 ;
        RECT 4.890 1.360 5.060 1.660 ;
        RECT 0.625 1.100 1.570 1.270 ;
        RECT 0.625 2.290 1.570 2.460 ;
        RECT 1.400 1.100 1.570 2.890 ;
        RECT 1.400 1.515 1.615 1.815 ;
        RECT 1.400 2.720 2.140 2.890 ;
        RECT 1.970 2.720 2.140 3.210 ;
        RECT 1.970 3.040 2.875 3.210 ;
        RECT 3.140 2.675 4.360 2.845 ;
        RECT 4.190 2.675 4.360 3.085 ;
        RECT 5.270 2.190 5.440 3.085 ;
        RECT 4.190 2.915 5.440 3.085 ;
        RECT 5.270 2.190 5.545 2.360 ;
        RECT 5.590 1.245 5.760 1.415 ;
        RECT 5.760 1.245 5.770 2.209 ;
        RECT 5.770 1.245 5.780 2.199 ;
        RECT 5.780 1.245 5.790 2.189 ;
        RECT 5.790 1.245 5.800 2.179 ;
        RECT 5.800 1.245 5.810 2.169 ;
        RECT 5.810 1.245 5.820 2.159 ;
        RECT 5.820 1.245 5.830 2.149 ;
        RECT 5.830 1.245 5.840 2.139 ;
        RECT 5.840 1.245 5.850 2.129 ;
        RECT 5.850 1.245 5.860 2.119 ;
        RECT 5.860 1.245 5.870 2.109 ;
        RECT 5.870 1.245 5.880 2.099 ;
        RECT 5.880 1.245 5.890 2.089 ;
        RECT 5.890 1.245 5.900 2.079 ;
        RECT 5.900 1.245 5.910 2.069 ;
        RECT 5.910 1.245 5.920 2.059 ;
        RECT 5.920 1.245 5.930 2.049 ;
        RECT 5.620 2.115 5.630 2.349 ;
        RECT 5.630 2.105 5.640 2.339 ;
        RECT 5.640 2.095 5.650 2.329 ;
        RECT 5.650 2.085 5.660 2.319 ;
        RECT 5.660 2.075 5.670 2.309 ;
        RECT 5.670 2.065 5.680 2.299 ;
        RECT 5.680 2.055 5.690 2.289 ;
        RECT 5.690 2.045 5.700 2.279 ;
        RECT 5.700 2.035 5.710 2.269 ;
        RECT 5.710 2.025 5.720 2.259 ;
        RECT 5.720 2.015 5.730 2.249 ;
        RECT 5.730 2.005 5.740 2.239 ;
        RECT 5.740 1.995 5.750 2.229 ;
        RECT 5.750 1.985 5.760 2.219 ;
        RECT 5.545 2.190 5.555 2.360 ;
        RECT 5.555 2.180 5.565 2.360 ;
        RECT 5.565 2.170 5.575 2.360 ;
        RECT 5.575 2.160 5.585 2.360 ;
        RECT 5.585 2.150 5.595 2.360 ;
        RECT 5.595 2.140 5.605 2.360 ;
        RECT 5.605 2.130 5.615 2.360 ;
        RECT 5.615 2.120 5.621 2.360 ;
        RECT 2.970 2.675 2.980 3.179 ;
        RECT 2.980 2.675 2.990 3.169 ;
        RECT 2.990 2.675 3.000 3.159 ;
        RECT 3.000 2.675 3.010 3.149 ;
        RECT 3.010 2.675 3.020 3.139 ;
        RECT 3.020 2.675 3.030 3.129 ;
        RECT 3.030 2.675 3.040 3.119 ;
        RECT 3.040 2.675 3.050 3.109 ;
        RECT 3.050 2.675 3.060 3.099 ;
        RECT 3.060 2.675 3.070 3.089 ;
        RECT 3.070 2.675 3.080 3.079 ;
        RECT 3.080 2.675 3.090 3.069 ;
        RECT 3.090 2.675 3.100 3.059 ;
        RECT 3.100 2.675 3.110 3.049 ;
        RECT 3.110 2.675 3.120 3.039 ;
        RECT 3.120 2.675 3.130 3.029 ;
        RECT 3.130 2.675 3.140 3.019 ;
        RECT 2.950 2.965 2.960 3.199 ;
        RECT 2.960 2.955 2.970 3.189 ;
        RECT 2.875 3.040 2.885 3.210 ;
        RECT 2.885 3.030 2.895 3.210 ;
        RECT 2.895 3.020 2.905 3.210 ;
        RECT 2.905 3.010 2.915 3.210 ;
        RECT 2.915 3.000 2.925 3.210 ;
        RECT 2.925 2.990 2.935 3.210 ;
        RECT 2.935 2.980 2.945 3.210 ;
        RECT 2.945 2.970 2.951 3.210 ;
        RECT 6.705 1.245 6.800 1.935 ;
        RECT 6.705 1.245 6.930 1.415 ;
        RECT 6.705 1.765 7.620 1.935 ;
        RECT 6.630 1.245 6.640 2.395 ;
        RECT 6.640 1.245 6.650 2.385 ;
        RECT 6.650 1.245 6.660 2.375 ;
        RECT 6.660 1.245 6.670 2.365 ;
        RECT 6.670 1.245 6.680 2.355 ;
        RECT 6.680 1.245 6.690 2.345 ;
        RECT 6.690 1.245 6.700 2.335 ;
        RECT 6.700 1.245 6.706 2.329 ;
        RECT 6.535 1.765 6.545 2.489 ;
        RECT 6.545 1.765 6.555 2.479 ;
        RECT 6.555 1.765 6.565 2.469 ;
        RECT 6.565 1.765 6.575 2.459 ;
        RECT 6.575 1.765 6.585 2.449 ;
        RECT 6.585 1.765 6.595 2.439 ;
        RECT 6.595 1.765 6.605 2.429 ;
        RECT 6.605 1.765 6.615 2.419 ;
        RECT 6.615 1.765 6.625 2.409 ;
        RECT 6.625 1.765 6.631 2.405 ;
        RECT 6.480 2.310 6.490 2.544 ;
        RECT 6.490 2.300 6.500 2.534 ;
        RECT 6.500 2.290 6.510 2.524 ;
        RECT 6.510 2.280 6.520 2.514 ;
        RECT 6.520 2.270 6.530 2.504 ;
        RECT 6.530 2.260 6.536 2.500 ;
        RECT 6.310 2.480 6.320 2.780 ;
        RECT 6.320 2.470 6.330 2.780 ;
        RECT 6.330 2.460 6.340 2.780 ;
        RECT 6.340 2.450 6.350 2.780 ;
        RECT 6.350 2.440 6.360 2.780 ;
        RECT 6.360 2.430 6.370 2.780 ;
        RECT 6.370 2.420 6.380 2.780 ;
        RECT 6.380 2.410 6.390 2.780 ;
        RECT 6.390 2.400 6.400 2.780 ;
        RECT 6.400 2.390 6.410 2.780 ;
        RECT 6.410 2.380 6.420 2.780 ;
        RECT 6.420 2.370 6.430 2.780 ;
        RECT 6.430 2.360 6.440 2.780 ;
        RECT 6.440 2.350 6.450 2.780 ;
        RECT 6.450 2.340 6.460 2.780 ;
        RECT 6.460 2.330 6.470 2.780 ;
        RECT 6.470 2.320 6.480 2.780 ;
        RECT 2.560 1.470 2.855 1.640 ;
        RECT 2.560 0.990 2.730 1.640 ;
        RECT 2.685 1.470 2.855 2.495 ;
        RECT 4.750 1.840 4.920 2.495 ;
        RECT 2.685 2.325 4.920 2.495 ;
        RECT 5.240 0.875 5.410 2.010 ;
        RECT 4.750 1.840 5.410 2.010 ;
        RECT 5.240 1.600 5.580 1.900 ;
        RECT 5.240 0.875 6.985 1.045 ;
        RECT 7.585 2.115 7.755 2.500 ;
        RECT 7.225 1.040 7.970 1.210 ;
        RECT 7.800 1.040 7.970 2.285 ;
        RECT 7.585 2.115 7.970 2.285 ;
        RECT 7.150 0.975 7.160 1.209 ;
        RECT 7.160 0.985 7.170 1.209 ;
        RECT 7.170 0.995 7.180 1.209 ;
        RECT 7.180 1.005 7.190 1.209 ;
        RECT 7.190 1.015 7.200 1.209 ;
        RECT 7.200 1.025 7.210 1.209 ;
        RECT 7.210 1.035 7.220 1.209 ;
        RECT 7.220 1.040 7.226 1.210 ;
        RECT 7.060 0.885 7.070 1.119 ;
        RECT 7.070 0.895 7.080 1.129 ;
        RECT 7.080 0.905 7.090 1.139 ;
        RECT 7.090 0.915 7.100 1.149 ;
        RECT 7.100 0.925 7.110 1.159 ;
        RECT 7.110 0.935 7.120 1.169 ;
        RECT 7.120 0.945 7.130 1.179 ;
        RECT 7.130 0.955 7.140 1.189 ;
        RECT 7.140 0.965 7.150 1.199 ;
        RECT 6.985 0.875 6.995 1.045 ;
        RECT 6.995 0.875 7.005 1.055 ;
        RECT 7.005 0.875 7.015 1.065 ;
        RECT 7.015 0.875 7.025 1.075 ;
        RECT 7.025 0.875 7.035 1.085 ;
        RECT 7.035 0.875 7.045 1.095 ;
        RECT 7.045 0.875 7.055 1.105 ;
        RECT 7.055 0.875 7.061 1.115 ;
        RECT 2.205 0.640 2.375 2.190 ;
        RECT 2.205 2.020 2.505 2.190 ;
        RECT 2.205 0.640 4.890 0.810 ;
        RECT 4.720 0.525 4.890 1.170 ;
        RECT 7.145 0.620 8.895 0.705 ;
        RECT 7.155 0.620 8.895 0.715 ;
        RECT 7.165 0.620 8.895 0.725 ;
        RECT 7.175 0.620 8.895 0.735 ;
        RECT 7.185 0.620 8.895 0.745 ;
        RECT 7.195 0.620 8.895 0.755 ;
        RECT 7.205 0.620 8.895 0.765 ;
        RECT 4.720 0.525 7.211 0.695 ;
        RECT 7.210 0.620 8.895 0.769 ;
        RECT 4.720 0.535 7.220 0.695 ;
        RECT 7.220 0.620 8.895 0.779 ;
        RECT 4.720 0.545 7.230 0.695 ;
        RECT 4.720 0.555 7.240 0.695 ;
        RECT 4.720 0.565 7.250 0.695 ;
        RECT 4.720 0.575 7.260 0.695 ;
        RECT 4.720 0.585 7.270 0.695 ;
        RECT 4.720 0.595 7.280 0.695 ;
        RECT 4.720 0.605 7.290 0.695 ;
        RECT 7.230 0.620 8.895 0.789 ;
        RECT 4.720 0.615 7.300 0.695 ;
        RECT 7.300 0.620 8.895 0.790 ;
        RECT 8.725 0.620 8.895 2.435 ;
        RECT 8.560 2.265 8.895 2.435 ;
        RECT 5.725 2.545 5.960 2.715 ;
        RECT 6.110 1.245 6.175 1.415 ;
        RECT 6.345 1.245 6.410 1.415 ;
        RECT 6.130 2.960 6.555 3.130 ;
        RECT 6.850 2.740 7.860 2.910 ;
        RECT 7.690 2.740 7.860 3.150 ;
        RECT 7.690 2.980 9.090 3.150 ;
        RECT 8.790 2.980 9.090 3.210 ;
        RECT 6.775 2.740 6.785 2.974 ;
        RECT 6.785 2.740 6.795 2.964 ;
        RECT 6.795 2.740 6.805 2.954 ;
        RECT 6.805 2.740 6.815 2.944 ;
        RECT 6.815 2.740 6.825 2.934 ;
        RECT 6.825 2.740 6.835 2.924 ;
        RECT 6.835 2.740 6.845 2.914 ;
        RECT 6.845 2.740 6.851 2.910 ;
        RECT 6.630 2.885 6.640 3.119 ;
        RECT 6.640 2.875 6.650 3.109 ;
        RECT 6.650 2.865 6.660 3.099 ;
        RECT 6.660 2.855 6.670 3.089 ;
        RECT 6.670 2.845 6.680 3.079 ;
        RECT 6.680 2.835 6.690 3.069 ;
        RECT 6.690 2.825 6.700 3.059 ;
        RECT 6.700 2.815 6.710 3.049 ;
        RECT 6.710 2.805 6.720 3.039 ;
        RECT 6.720 2.795 6.730 3.029 ;
        RECT 6.730 2.785 6.740 3.019 ;
        RECT 6.740 2.775 6.750 3.009 ;
        RECT 6.750 2.765 6.760 2.999 ;
        RECT 6.760 2.755 6.770 2.989 ;
        RECT 6.770 2.745 6.776 2.985 ;
        RECT 6.555 2.960 6.565 3.130 ;
        RECT 6.565 2.950 6.575 3.130 ;
        RECT 6.575 2.940 6.585 3.130 ;
        RECT 6.585 2.930 6.595 3.130 ;
        RECT 6.595 2.920 6.605 3.130 ;
        RECT 6.605 2.910 6.615 3.130 ;
        RECT 6.615 2.900 6.625 3.130 ;
        RECT 6.625 2.890 6.631 3.130 ;
        RECT 6.175 1.245 6.185 2.325 ;
        RECT 6.185 1.245 6.195 2.315 ;
        RECT 6.195 1.245 6.205 2.305 ;
        RECT 6.205 1.245 6.215 2.295 ;
        RECT 6.215 1.245 6.225 2.285 ;
        RECT 6.225 1.245 6.235 2.275 ;
        RECT 6.235 1.245 6.245 2.265 ;
        RECT 6.245 1.245 6.255 2.255 ;
        RECT 6.255 1.245 6.265 2.245 ;
        RECT 6.265 1.245 6.275 2.235 ;
        RECT 6.275 1.245 6.285 2.225 ;
        RECT 6.285 1.245 6.295 2.215 ;
        RECT 6.295 1.245 6.305 2.205 ;
        RECT 6.305 1.245 6.315 2.195 ;
        RECT 6.315 1.245 6.325 2.185 ;
        RECT 6.325 1.245 6.335 2.175 ;
        RECT 6.335 1.245 6.345 2.165 ;
        RECT 6.130 2.135 6.140 2.369 ;
        RECT 6.140 2.125 6.150 2.359 ;
        RECT 6.150 2.115 6.160 2.349 ;
        RECT 6.160 2.105 6.170 2.339 ;
        RECT 6.170 2.095 6.176 2.335 ;
        RECT 5.960 2.305 5.970 3.129 ;
        RECT 5.970 2.295 5.980 3.129 ;
        RECT 5.980 2.285 5.990 3.129 ;
        RECT 5.990 2.275 6.000 3.129 ;
        RECT 6.000 2.265 6.010 3.129 ;
        RECT 6.010 2.255 6.020 3.129 ;
        RECT 6.020 2.245 6.030 3.129 ;
        RECT 6.030 2.235 6.040 3.129 ;
        RECT 6.040 2.225 6.050 3.129 ;
        RECT 6.050 2.215 6.060 3.129 ;
        RECT 6.060 2.205 6.070 3.129 ;
        RECT 6.070 2.195 6.080 3.129 ;
        RECT 6.080 2.185 6.090 3.129 ;
        RECT 6.090 2.175 6.100 3.129 ;
        RECT 6.100 2.165 6.110 3.129 ;
        RECT 6.110 2.155 6.120 3.129 ;
        RECT 6.120 2.145 6.130 3.129 ;
        RECT 8.205 1.010 8.375 2.800 ;
        RECT 8.105 2.490 8.375 2.800 ;
        RECT 9.135 2.460 9.305 2.800 ;
        RECT 8.105 2.630 9.305 2.800 ;
        RECT 9.135 2.460 10.005 2.630 ;
        RECT 9.835 1.545 10.005 2.630 ;
  END 
END FAHD1XHT

MACRO DEL4HDMXSPGHT
  CLASS  CORE ;
  FOREIGN DEL4HDMXSPGHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 0.755 0.425 1.295 3.065 ;
      LAYER V7 ;
        RECT 0.845 1.255 1.205 1.615 ;
      LAYER M7 ;
        RECT 0.290 1.245 1.350 1.625 ;
      LAYER V6 ;
        RECT 0.930 1.340 1.120 1.530 ;
      LAYER M4 ;
        RECT 0.515 1.210 0.715 2.440 ;
      LAYER V3 ;
        RECT 0.520 2.160 0.710 2.350 ;
      LAYER M3 ;
        RECT 0.105 2.070 0.815 2.440 ;
      LAYER V2 ;
        RECT 0.110 2.160 0.300 2.350 ;
      LAYER M2 ;
        RECT 0.105 2.070 0.305 2.890 ;
      LAYER V1 ;
        RECT 0.110 2.570 0.300 2.760 ;
      LAYER M1 ;
        RECT 0.095 2.470 0.510 2.890 ;
      LAYER M6 ;
        RECT 0.925 0.425 1.125 2.375 ;
      LAYER V5 ;
        RECT 0.930 1.340 1.120 1.530 ;
      LAYER M5 ;
        RECT 0.290 1.335 1.350 1.535 ;
      LAYER V4 ;
        RECT 0.520 1.340 0.710 1.530 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 -0.300 0.860 1.360 ;
        RECT 2.830 -0.300 3.000 0.850 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 2.395 0.325 2.935 3.060 ;
      LAYER V7 ;
        RECT 2.485 0.435 2.845 0.795 ;
      LAYER M7 ;
        RECT 2.390 0.425 3.175 0.805 ;
      LAYER V6 ;
        RECT 2.570 0.520 2.760 0.710 ;
      LAYER M4 ;
        RECT 2.975 0.440 3.175 1.210 ;
      LAYER V3 ;
        RECT 2.980 0.930 3.170 1.120 ;
      LAYER M3 ;
        RECT 2.795 0.840 3.585 1.210 ;
      LAYER V2 ;
        RECT 3.390 0.930 3.580 1.120 ;
      LAYER M2 ;
        RECT 3.385 0.855 3.585 1.600 ;
      LAYER V1 ;
        RECT 3.390 1.340 3.580 1.530 ;
      LAYER M1 ;
        RECT 3.350 0.700 3.520 2.580 ;
        RECT 3.350 1.250 3.590 1.600 ;
      LAYER M6 ;
        RECT 2.565 0.325 2.765 2.375 ;
      LAYER V5 ;
        RECT 2.570 0.520 2.760 0.710 ;
      LAYER M5 ;
        RECT 2.390 0.515 3.245 0.715 ;
      LAYER V4 ;
        RECT 2.980 0.520 3.170 0.710 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.100 0.860 3.990 ;
        RECT 2.765 2.675 3.065 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.540 1.200 1.840 ;
        RECT 1.630 1.060 1.800 2.280 ;
        RECT 1.630 1.585 2.465 1.755 ;
        RECT 1.825 0.615 2.370 0.785 ;
        RECT 2.200 0.615 2.370 1.265 ;
        RECT 2.290 2.160 2.460 2.845 ;
        RECT 1.820 2.675 2.460 2.845 ;
        RECT 2.200 1.095 3.170 1.265 ;
        RECT 3.000 1.095 3.170 2.330 ;
        RECT 2.290 2.160 3.170 2.330 ;
  END 
END DEL4HDMXSPGHT

MACRO DEL4HD1XHT
  CLASS  CORE ;
  FOREIGN DEL4HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.510 2.885 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 2.765 -0.300 3.065 0.785 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.350 0.720 3.520 2.960 ;
        RECT 3.350 1.250 3.590 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.100 0.860 3.990 ;
        RECT 2.765 2.790 3.065 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.605 1.380 1.775 ;
        RECT 1.630 1.060 1.800 2.280 ;
        RECT 1.630 1.605 2.465 1.775 ;
        RECT 1.825 0.615 2.370 0.785 ;
        RECT 2.200 0.615 2.370 1.210 ;
        RECT 2.290 2.335 2.460 2.845 ;
        RECT 1.820 2.675 2.460 2.845 ;
        RECT 2.200 1.040 3.170 1.210 ;
        RECT 3.000 1.040 3.170 2.505 ;
        RECT 2.290 2.335 3.170 2.505 ;
  END 
END DEL4HD1XHT

MACRO DEL3HDMXHT
  CLASS  CORE ;
  FOREIGN DEL3HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.510 2.840 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 2.355 -0.300 2.655 0.785 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.940 0.700 3.110 2.580 ;
        RECT 2.940 1.250 3.180 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.100 0.860 3.990 ;
        RECT 2.355 2.675 2.655 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.605 1.265 1.775 ;
        RECT 1.490 1.060 1.660 2.280 ;
        RECT 1.490 1.585 2.195 1.755 ;
        RECT 1.555 0.615 2.130 0.785 ;
        RECT 1.960 0.615 2.130 1.240 ;
        RECT 2.005 2.060 2.175 2.845 ;
        RECT 1.555 2.675 2.175 2.845 ;
        RECT 1.960 1.070 2.760 1.240 ;
        RECT 2.590 1.070 2.760 2.230 ;
        RECT 2.005 2.060 2.760 2.230 ;
  END 
END DEL3HDMXHT

MACRO DEL3HD1XHT
  CLASS  CORE ;
  FOREIGN DEL3HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.510 2.870 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 2.355 -0.300 2.655 0.785 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.940 0.720 3.110 2.960 ;
        RECT 2.940 1.250 3.180 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.100 0.860 3.990 ;
        RECT 2.355 2.790 2.655 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.605 1.265 1.775 ;
        RECT 1.490 1.060 1.660 2.280 ;
        RECT 1.490 1.585 2.195 1.755 ;
        RECT 1.555 0.615 2.175 0.785 ;
        RECT 2.005 0.615 2.175 1.215 ;
        RECT 2.005 2.335 2.175 2.845 ;
        RECT 1.555 2.675 2.175 2.845 ;
        RECT 2.005 1.045 2.760 1.215 ;
        RECT 2.590 1.045 2.760 2.505 ;
        RECT 2.005 2.335 2.760 2.505 ;
  END 
END DEL3HD1XHT

MACRO DEL2HDMXHT
  CLASS  CORE ;
  FOREIGN DEL2HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 2.470 0.510 2.865 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 2.355 -0.300 2.655 0.805 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.940 0.720 3.110 2.470 ;
        RECT 2.940 1.250 3.180 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.100 0.860 3.990 ;
        RECT 2.355 2.565 2.655 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.540 1.170 1.840 ;
        RECT 1.350 1.060 1.520 2.280 ;
        RECT 1.350 1.520 2.250 1.820 ;
        RECT 1.760 0.570 1.930 1.220 ;
        RECT 1.760 2.055 1.930 2.800 ;
        RECT 1.760 1.050 2.760 1.220 ;
        RECT 2.590 1.050 2.760 2.225 ;
        RECT 1.760 2.055 2.760 2.225 ;
  END 
END DEL2HDMXHT

MACRO DEL1HDMXHT
  CLASS  CORE ;
  FOREIGN DEL1HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 2.470 0.510 2.860 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 1.945 -0.300 2.245 0.785 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.530 0.700 2.700 2.580 ;
        RECT 2.530 1.250 2.770 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.100 0.860 3.990 ;
        RECT 1.945 2.675 2.245 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.540 1.030 1.840 ;
        RECT 1.210 1.060 1.380 2.280 ;
        RECT 1.210 1.585 1.905 1.755 ;
        RECT 1.425 0.615 1.765 0.785 ;
        RECT 1.595 0.615 1.765 1.245 ;
        RECT 1.595 2.290 1.765 2.845 ;
        RECT 1.425 2.675 1.765 2.845 ;
        RECT 1.595 1.075 2.350 1.245 ;
        RECT 2.180 1.075 2.350 2.460 ;
        RECT 1.595 2.290 2.350 2.460 ;
  END 
END DEL1HDMXHT

MACRO DEL2HD1XHT
  CLASS  CORE ;
  FOREIGN DEL2HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.510 2.855 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 -0.300 0.860 1.360 ;
        RECT 2.120 -0.300 2.420 0.785 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.705 0.720 2.875 2.960 ;
        RECT 2.705 1.250 3.185 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.100 0.860 3.990 ;
        RECT 2.120 2.790 2.420 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.540 1.170 1.840 ;
        RECT 1.350 1.060 1.520 2.280 ;
        RECT 1.350 1.585 1.940 1.755 ;
        RECT 1.460 0.615 1.940 0.785 ;
        RECT 1.770 0.615 1.940 1.215 ;
        RECT 1.770 2.335 1.940 2.845 ;
        RECT 1.460 2.675 1.940 2.845 ;
        RECT 1.770 1.045 2.525 1.215 ;
        RECT 2.355 1.045 2.525 2.505 ;
        RECT 1.770 2.335 2.525 2.505 ;
  END 
END DEL2HD1XHT

MACRO DEL1HDMXSPGHT
  CLASS  CORE ;
  FOREIGN DEL1HDMXSPGHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 0.325 0.425 0.905 3.075 ;
      LAYER V7 ;
        RECT 0.435 0.845 0.795 1.205 ;
      LAYER M7 ;
        RECT 0.225 0.835 1.015 1.215 ;
      LAYER V6 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M4 ;
        RECT 0.515 0.815 0.715 2.010 ;
      LAYER V3 ;
        RECT 0.520 1.750 0.710 1.940 ;
      LAYER M3 ;
        RECT 0.105 1.680 0.835 2.010 ;
      LAYER V2 ;
        RECT 0.110 1.750 0.300 1.940 ;
      LAYER M2 ;
        RECT 0.105 1.670 0.305 2.905 ;
      LAYER V1 ;
        RECT 0.110 2.570 0.300 2.760 ;
      LAYER M1 ;
        RECT 0.095 2.470 0.510 2.860 ;
      LAYER M6 ;
        RECT 0.515 0.425 0.715 2.305 ;
      LAYER V5 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M5 ;
        RECT 0.225 0.925 1.015 1.125 ;
      LAYER V4 ;
        RECT 0.520 0.930 0.710 1.120 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 -0.300 0.860 1.360 ;
        RECT 1.945 -0.300 2.245 0.785 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 1.965 0.330 2.545 3.070 ;
      LAYER V7 ;
        RECT 2.075 0.435 2.435 0.795 ;
      LAYER M7 ;
        RECT 1.755 0.425 2.675 0.805 ;
      LAYER V6 ;
        RECT 2.160 0.520 2.350 0.710 ;
      LAYER M4 ;
        RECT 2.155 0.405 2.355 1.325 ;
      LAYER V3 ;
        RECT 2.160 0.930 2.350 1.120 ;
      LAYER M3 ;
        RECT 2.140 0.840 2.765 1.210 ;
      LAYER V2 ;
        RECT 2.570 0.930 2.760 1.120 ;
      LAYER M2 ;
        RECT 2.565 0.850 2.765 1.670 ;
      LAYER V1 ;
        RECT 2.570 1.340 2.760 1.530 ;
      LAYER M1 ;
        RECT 2.530 0.700 2.700 2.580 ;
        RECT 2.530 1.250 2.770 1.600 ;
      LAYER M6 ;
        RECT 2.155 0.330 2.355 2.405 ;
      LAYER V5 ;
        RECT 2.160 0.520 2.350 0.710 ;
      LAYER M5 ;
        RECT 1.755 0.515 2.675 0.715 ;
      LAYER V4 ;
        RECT 2.160 0.520 2.350 0.710 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.100 0.860 3.990 ;
        RECT 1.945 2.675 2.245 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.540 1.030 1.840 ;
        RECT 1.210 1.060 1.380 2.280 ;
        RECT 1.210 1.585 1.905 1.755 ;
        RECT 1.425 0.615 1.765 0.785 ;
        RECT 1.595 0.615 1.765 1.245 ;
        RECT 1.595 2.290 1.765 2.845 ;
        RECT 1.425 2.675 1.765 2.845 ;
        RECT 1.595 1.075 2.350 1.245 ;
        RECT 2.180 1.075 2.350 2.460 ;
        RECT 1.595 2.290 2.350 2.460 ;
  END 
END DEL1HDMXSPGHT

MACRO DEL1HD1XHT
  CLASS  CORE ;
  FOREIGN DEL1HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.510 2.885 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 1.945 -0.300 2.245 0.785 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.530 0.720 2.700 2.960 ;
        RECT 2.530 1.250 2.770 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.100 0.860 3.990 ;
        RECT 1.945 2.795 2.245 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.540 1.030 1.840 ;
        RECT 1.210 1.060 1.380 2.280 ;
        RECT 1.210 1.585 1.905 1.755 ;
        RECT 1.425 0.615 1.765 0.785 ;
        RECT 1.595 0.615 1.765 1.245 ;
        RECT 1.595 2.290 1.765 2.845 ;
        RECT 1.425 2.675 1.765 2.845 ;
        RECT 1.595 1.075 2.350 1.245 ;
        RECT 2.180 1.075 2.350 2.460 ;
        RECT 1.595 2.290 2.350 2.460 ;
  END 
END DEL1HD1XHT

MACRO BUFTSHDUXHT
  CLASS  CORE ;
  FOREIGN BUFTSHDUXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.540 1.265 1.130 1.845 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.240 2.360 2.015 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.685 -0.300 0.985 1.085 ;
        RECT 1.720 -0.300 1.955 0.850 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 1.720 1.060 1.950 2.280 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.685 2.045 0.985 3.990 ;
        RECT 1.655 2.490 1.955 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.920 ;
        RECT 2.235 0.615 2.710 0.785 ;
        RECT 2.410 2.555 2.580 3.210 ;
        RECT 2.540 0.615 2.710 2.725 ;
        RECT 2.235 2.555 2.710 2.725 ;
  END 
END BUFTSHDUXHT

MACRO BUFTSHDMXHT
  CLASS  CORE ;
  FOREIGN BUFTSHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.470 0.520 2.835 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.370 1.520 2.770 2.015 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 -0.300 0.835 0.745 ;
        RECT 2.465 -0.300 2.765 0.745 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 1.260 2.150 1.690 2.360 ;
        RECT 1.520 1.060 1.690 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 3.095 0.835 3.990 ;
        RECT 2.465 2.875 2.765 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.060 0.345 1.755 ;
        RECT 0.170 1.585 1.085 1.755 ;
        RECT 1.885 1.120 2.065 2.380 ;
        RECT 1.885 1.120 2.265 1.300 ;
        RECT 1.885 2.200 2.265 2.380 ;
  END 
END BUFTSHDMXHT

MACRO LATHD2XHT
  CLASS  CORE ;
  FOREIGN LATHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.970 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 6.110 0.720 6.280 2.960 ;
        RECT 6.110 1.260 6.460 1.600 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.050 0.720 5.240 1.195 ;
        RECT 5.020 0.850 5.240 1.195 ;
        RECT 5.070 0.720 5.240 2.280 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.945 1.585 2.445 1.950 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.495 0.510 2.950 ;
    END
  END G
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.565 -0.300 0.865 0.745 ;
        RECT 1.780 -0.300 1.950 1.040 ;
        RECT 3.495 -0.300 3.795 1.295 ;
        RECT 4.485 -0.300 4.785 0.715 ;
        RECT 5.525 -0.300 5.825 1.055 ;
        RECT 6.565 -0.300 6.865 1.060 ;
        RECT 0.000 -0.300 6.970 0.300 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.280 0.860 3.990 ;
        RECT 1.715 2.635 2.015 3.990 ;
        RECT 3.465 2.895 3.765 3.990 ;
        RECT 4.485 2.975 4.785 3.990 ;
        RECT 5.525 2.975 5.825 3.990 ;
        RECT 6.565 2.295 6.865 3.990 ;
        RECT 0.000 3.390 6.970 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.520 1.000 1.820 ;
        RECT 1.180 0.525 1.350 2.305 ;
        RECT 1.180 1.980 1.380 2.305 ;
        RECT 1.180 0.525 1.560 0.695 ;
        RECT 1.180 2.135 2.440 2.305 ;
        RECT 2.270 2.135 2.440 3.095 ;
        RECT 2.270 2.925 3.185 3.095 ;
        RECT 1.530 1.230 1.700 1.820 ;
        RECT 2.195 0.515 2.365 1.400 ;
        RECT 1.530 1.230 2.365 1.400 ;
        RECT 2.195 0.515 3.185 0.685 ;
        RECT 3.315 1.825 3.615 1.995 ;
        RECT 3.445 1.825 3.615 2.365 ;
        RECT 4.015 1.125 4.840 1.295 ;
        RECT 4.670 1.125 4.840 2.365 ;
        RECT 3.445 2.195 4.840 2.365 ;
        RECT 2.670 1.060 2.840 2.715 ;
        RECT 2.670 1.475 4.135 1.645 ;
        RECT 3.835 1.475 4.135 1.665 ;
        RECT 5.760 1.520 5.930 2.715 ;
        RECT 2.670 2.545 5.930 2.715 ;
  END 
END LATHD2XHT

MACRO BUFTSHD2XHT
  CLASS  CORE ;
  FOREIGN BUFTSHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.375 1.650 4.820 2.015 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.310 2.015 ;
        RECT 0.100 1.520 0.520 1.820 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.945 ;
        RECT 2.955 -0.300 3.255 1.015 ;
        RECT 3.995 -0.300 4.295 0.995 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 2.500 1.060 2.670 1.360 ;
        RECT 2.500 1.195 3.710 1.360 ;
        RECT 2.560 1.060 2.670 2.760 ;
        RECT 2.500 2.120 2.670 2.760 ;
        RECT 2.560 1.195 2.770 2.430 ;
        RECT 2.500 2.120 2.770 2.430 ;
        RECT 2.500 2.260 3.775 2.430 ;
        RECT 3.540 1.060 3.710 1.365 ;
        RECT 2.560 1.195 3.710 1.365 ;
        RECT 3.475 2.260 3.775 2.770 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.705 2.460 1.005 3.990 ;
        RECT 2.955 2.705 3.255 3.990 ;
        RECT 3.995 2.705 4.295 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.455 2.145 1.100 2.280 ;
        RECT 0.465 2.135 0.495 2.365 ;
        RECT 0.445 2.155 1.100 2.280 ;
        RECT 0.475 2.125 0.495 2.365 ;
        RECT 0.435 2.165 1.100 2.280 ;
        RECT 0.485 2.115 0.495 2.365 ;
        RECT 0.425 2.175 1.100 2.280 ;
        RECT 0.105 2.195 0.495 2.365 ;
        RECT 0.105 2.195 0.505 2.354 ;
        RECT 0.105 2.195 0.515 2.344 ;
        RECT 0.105 2.195 0.525 2.334 ;
        RECT 0.105 2.195 0.535 2.324 ;
        RECT 0.105 2.195 0.545 2.314 ;
        RECT 0.105 2.195 0.555 2.304 ;
        RECT 0.105 2.195 0.565 2.294 ;
        RECT 0.105 2.195 0.575 2.284 ;
        RECT 0.105 1.125 1.100 1.295 ;
        RECT 0.490 2.110 1.100 2.280 ;
        RECT 0.415 2.185 1.100 2.280 ;
        RECT 0.930 1.125 1.100 2.280 ;
        RECT 1.320 1.680 1.490 2.620 ;
        RECT 1.800 1.060 1.970 1.850 ;
        RECT 1.320 1.680 1.970 1.850 ;
        RECT 1.320 2.415 2.305 2.620 ;
        RECT 1.280 0.710 1.450 1.360 ;
        RECT 1.280 0.710 2.320 0.880 ;
        RECT 2.150 0.710 2.320 2.215 ;
        RECT 1.805 2.045 2.320 2.215 ;
        RECT 3.240 1.750 3.410 2.080 ;
        RECT 3.240 1.910 4.125 2.080 ;
        RECT 3.955 1.910 4.125 2.365 ;
        RECT 3.955 2.195 4.750 2.365 ;
        RECT 4.580 2.195 4.750 2.835 ;
        RECT 3.890 1.300 4.060 1.730 ;
        RECT 4.580 0.720 4.750 1.470 ;
        RECT 3.890 1.300 4.750 1.470 ;
  END 
END BUFTSHD2XHT

MACRO BUFTSHD1XHT
  CLASS  CORE ;
  FOREIGN BUFTSHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.490 1.460 0.720 2.015 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 2.710 1.210 3.180 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.595 ;
        RECT 3.155 -0.300 3.455 1.025 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 2.115 1.125 2.415 2.555 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.440 3.010 0.610 3.990 ;
        RECT 3.155 2.545 3.455 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.085 1.125 1.460 1.295 ;
        RECT 1.290 1.125 1.460 2.375 ;
        RECT 1.085 2.205 1.460 2.375 ;
        RECT 0.105 1.110 0.275 2.685 ;
        RECT 0.105 2.175 0.405 2.685 ;
        RECT 0.715 0.775 0.885 1.280 ;
        RECT 0.105 1.110 0.885 1.280 ;
        RECT 1.290 0.480 1.460 0.945 ;
        RECT 0.715 0.775 1.460 0.945 ;
        RECT 1.660 2.140 1.830 3.120 ;
        RECT 2.700 2.110 2.870 3.120 ;
        RECT 1.660 2.950 2.870 3.120 ;
        RECT 2.700 2.110 3.910 2.280 ;
        RECT 3.740 2.110 3.910 3.120 ;
        RECT 1.660 0.775 1.830 1.080 ;
        RECT 1.660 0.775 2.870 0.945 ;
        RECT 2.700 0.775 2.870 1.375 ;
        RECT 3.740 1.060 3.910 1.375 ;
        RECT 2.700 1.205 3.910 1.375 ;
  END 
END BUFTSHD1XHT

MACRO BUFTSHDLXHT
  CLASS  CORE ;
  FOREIGN BUFTSHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.510 2.015 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.335 1.495 2.770 2.015 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.635 -0.300 0.935 0.655 ;
        RECT 2.465 -0.300 2.765 1.295 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 1.480 1.060 1.670 2.835 ;
        RECT 1.325 2.495 1.670 2.835 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.635 3.075 0.935 3.990 ;
        RECT 2.465 2.325 2.765 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.510 0.340 1.205 ;
        RECT 0.170 2.225 0.340 2.950 ;
        RECT 0.170 1.035 1.000 1.205 ;
        RECT 0.830 1.035 1.000 2.395 ;
        RECT 0.170 2.225 1.000 2.395 ;
        RECT 1.865 1.120 2.045 2.380 ;
        RECT 1.865 1.120 2.245 1.300 ;
        RECT 1.865 2.200 2.245 2.380 ;
  END 
END BUFTSHDLXHT

MACRO BUFTSHD8XHT
  CLASS  CORE ;
  FOREIGN BUFTSHD8XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.250 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 8.520 1.575 9.745 1.745 ;
        RECT 9.520 1.575 9.745 2.015 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.095 1.610 0.635 2.015 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.695 -0.300 0.995 0.715 ;
        RECT 3.735 -0.300 4.035 1.055 ;
        RECT 4.775 -0.300 5.075 1.055 ;
        RECT 5.815 -0.300 6.115 1.055 ;
        RECT 6.855 -0.300 7.155 1.055 ;
        RECT 8.635 -0.300 8.935 0.715 ;
        RECT 9.675 -0.300 9.975 1.055 ;
        RECT 0.000 -0.300 10.250 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 3.280 0.720 3.450 2.965 ;
        RECT 4.255 0.785 4.555 2.895 ;
        RECT 5.295 0.785 5.595 2.895 ;
        RECT 6.335 0.785 6.635 2.895 ;
        RECT 3.280 1.360 7.610 2.090 ;
        RECT 7.440 0.720 7.610 2.960 ;
        RECT 7.430 1.360 7.610 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.695 2.975 0.995 3.990 ;
        RECT 3.735 2.290 4.035 3.990 ;
        RECT 4.775 2.290 5.075 3.990 ;
        RECT 5.815 2.290 6.115 3.990 ;
        RECT 6.855 2.290 7.155 3.990 ;
        RECT 8.635 2.630 8.935 3.990 ;
        RECT 9.675 2.295 9.975 3.990 ;
        RECT 0.000 3.390 10.250 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.090 0.480 0.410 0.650 ;
        RECT 0.240 0.480 0.410 1.360 ;
        RECT 0.240 1.190 1.060 1.360 ;
        RECT 0.890 1.190 1.060 2.390 ;
        RECT 0.175 2.215 1.060 2.390 ;
        RECT 0.890 2.040 1.730 2.210 ;
        RECT 1.560 2.040 1.730 2.340 ;
        RECT 1.280 0.720 1.450 1.690 ;
        RECT 1.955 1.490 2.125 2.700 ;
        RECT 1.825 2.530 2.125 2.700 ;
        RECT 2.340 1.085 2.645 1.690 ;
        RECT 2.340 1.390 2.720 1.690 ;
        RECT 1.280 1.490 2.720 1.690 ;
        RECT 1.280 2.520 1.450 3.170 ;
        RECT 1.890 0.705 2.060 1.020 ;
        RECT 2.410 2.040 2.580 3.170 ;
        RECT 1.280 2.990 2.580 3.170 ;
        RECT 1.890 0.705 3.080 0.905 ;
        RECT 2.910 0.705 3.080 2.210 ;
        RECT 2.410 2.040 3.080 2.210 ;
        RECT 7.810 1.770 7.980 2.380 ;
        RECT 8.180 2.200 8.350 3.180 ;
        RECT 7.810 2.200 9.395 2.380 ;
        RECT 9.215 2.200 9.395 3.180 ;
        RECT 7.810 1.195 7.980 1.570 ;
        RECT 8.180 0.720 8.350 1.375 ;
        RECT 9.215 0.720 9.395 1.375 ;
        RECT 7.810 1.195 9.395 1.375 ;
  END 
END BUFTSHD8XHT

MACRO BUFTSHD7XHT
  CLASS  CORE ;
  FOREIGN BUFTSHD7XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.660 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 8.435 1.585 10.560 1.755 ;
        RECT 10.350 1.585 10.560 2.015 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.580 0.510 2.015 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.995 ;
        RECT 1.695 -0.300 1.995 0.995 ;
        RECT 4.465 -0.300 4.765 1.055 ;
        RECT 5.505 -0.300 5.805 1.055 ;
        RECT 6.545 -0.300 6.845 1.055 ;
        RECT 7.585 -0.300 7.820 1.120 ;
        RECT 8.095 -0.300 8.395 0.835 ;
        RECT 9.135 -0.300 9.435 0.835 ;
        RECT 10.175 -0.300 10.475 0.835 ;
        RECT 0.000 -0.300 10.660 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 4.010 0.480 4.245 3.210 ;
        RECT 4.985 0.720 5.285 2.965 ;
        RECT 4.010 1.290 5.430 2.045 ;
        RECT 6.025 0.720 6.325 2.960 ;
        RECT 4.010 1.295 7.365 2.045 ;
        RECT 7.065 0.720 7.365 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.745 0.955 3.990 ;
        RECT 1.695 2.745 1.995 3.990 ;
        RECT 4.465 2.295 4.765 3.990 ;
        RECT 5.505 2.295 5.805 3.990 ;
        RECT 6.545 2.295 6.845 3.990 ;
        RECT 7.585 2.230 7.820 3.990 ;
        RECT 8.095 2.405 8.395 3.990 ;
        RECT 9.135 2.405 9.435 3.990 ;
        RECT 10.175 2.405 10.475 3.990 ;
        RECT 0.000 3.390 10.660 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 1.360 ;
        RECT 0.170 1.190 1.020 1.360 ;
        RECT 0.850 1.190 1.020 2.375 ;
        RECT 0.105 2.205 1.020 2.375 ;
        RECT 0.850 1.815 2.455 1.985 ;
        RECT 1.240 1.060 1.410 1.560 ;
        RECT 1.240 1.390 2.960 1.560 ;
        RECT 2.790 1.060 2.960 2.740 ;
        RECT 1.240 2.340 1.410 2.980 ;
        RECT 1.240 2.340 2.440 2.510 ;
        RECT 2.270 0.710 2.440 1.160 ;
        RECT 2.270 2.340 2.440 3.090 ;
        RECT 2.270 0.710 3.480 0.880 ;
        RECT 3.310 0.710 3.480 3.090 ;
        RECT 2.270 2.920 3.480 3.090 ;
        RECT 3.310 2.070 3.810 2.370 ;
        RECT 8.020 1.770 8.190 2.225 ;
        RECT 8.680 2.055 8.850 2.780 ;
        RECT 8.020 2.055 9.890 2.225 ;
        RECT 9.720 2.055 9.890 2.780 ;
        RECT 8.020 1.030 8.190 1.570 ;
        RECT 8.680 0.900 8.850 1.200 ;
        RECT 9.720 0.900 9.890 1.200 ;
        RECT 8.020 1.030 9.890 1.200 ;
  END 
END BUFTSHD7XHT

MACRO BUFTSHD6XHT
  CLASS  CORE ;
  FOREIGN BUFTSHD6XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.200 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 7.085 1.585 8.100 1.755 ;
        RECT 7.890 1.585 8.100 2.015 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.540 0.560 2.015 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.585 -0.300 0.885 0.715 ;
        RECT 2.950 -0.300 3.185 1.120 ;
        RECT 3.925 -0.300 4.225 1.055 ;
        RECT 4.965 -0.300 5.265 1.055 ;
        RECT 6.005 -0.300 6.240 1.120 ;
        RECT 6.745 -0.300 7.045 1.055 ;
        RECT 7.785 -0.300 8.085 1.055 ;
        RECT 0.000 -0.300 8.200 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 3.405 0.720 3.705 2.965 ;
        RECT 4.445 0.720 4.745 2.960 ;
        RECT 3.405 1.295 5.785 2.045 ;
        RECT 5.485 0.720 5.785 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.615 2.975 0.915 3.990 ;
        RECT 2.950 2.230 3.185 3.990 ;
        RECT 3.925 2.295 4.225 3.990 ;
        RECT 4.965 2.295 5.265 3.990 ;
        RECT 6.005 2.230 6.240 3.990 ;
        RECT 6.745 2.295 7.045 3.990 ;
        RECT 7.785 2.295 8.085 3.990 ;
        RECT 0.000 3.390 8.200 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.090 0.480 0.390 0.650 ;
        RECT 0.220 0.480 0.390 1.360 ;
        RECT 0.220 1.190 0.910 1.360 ;
        RECT 0.740 1.190 0.910 2.375 ;
        RECT 0.155 2.205 0.910 2.375 ;
        RECT 0.740 2.040 1.650 2.210 ;
        RECT 1.480 2.040 1.650 2.340 ;
        RECT 1.200 1.060 1.370 1.600 ;
        RECT 1.895 1.430 2.065 2.800 ;
        RECT 1.685 2.630 2.065 2.800 ;
        RECT 1.895 1.840 2.195 2.010 ;
        RECT 2.240 1.060 2.410 1.600 ;
        RECT 1.200 1.430 2.410 1.600 ;
        RECT 1.200 2.520 1.370 3.160 ;
        RECT 1.720 0.710 1.890 1.210 ;
        RECT 2.270 2.225 2.440 3.160 ;
        RECT 1.200 2.990 2.440 3.160 ;
        RECT 1.720 0.710 2.760 0.880 ;
        RECT 2.515 2.095 2.760 2.395 ;
        RECT 2.590 0.710 2.760 2.395 ;
        RECT 2.270 2.225 2.760 2.395 ;
        RECT 6.440 1.770 6.610 2.115 ;
        RECT 6.440 1.945 7.500 2.115 ;
        RECT 7.330 1.945 7.500 2.960 ;
        RECT 6.440 1.235 6.610 1.570 ;
        RECT 7.330 0.720 7.500 1.405 ;
        RECT 6.440 1.235 7.500 1.405 ;
  END 
END BUFTSHD6XHT

MACRO BUFTSHD5XHT
  CLASS  CORE ;
  FOREIGN BUFTSHD5XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.380 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 6.025 1.585 6.870 1.755 ;
        RECT 6.660 1.585 6.870 2.015 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.555 0.570 2.015 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.595 -0.300 0.895 0.745 ;
        RECT 3.045 -0.300 3.345 1.055 ;
        RECT 4.085 -0.300 4.385 1.055 ;
        RECT 5.125 -0.300 5.425 1.055 ;
        RECT 5.685 -0.300 5.985 0.795 ;
        RECT 6.725 -0.300 7.025 1.135 ;
        RECT 0.000 -0.300 7.380 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 2.590 0.720 2.825 2.965 ;
        RECT 3.565 0.720 3.865 2.960 ;
        RECT 2.590 1.295 4.905 2.045 ;
        RECT 4.605 0.720 4.905 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.975 0.925 3.990 ;
        RECT 3.045 2.295 3.345 3.990 ;
        RECT 4.085 2.295 4.385 3.990 ;
        RECT 5.125 2.295 5.425 3.990 ;
        RECT 5.685 2.525 5.985 3.990 ;
        RECT 6.725 2.525 7.025 3.990 ;
        RECT 0.000 3.390 7.380 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.100 0.480 0.400 0.650 ;
        RECT 0.230 0.480 0.400 1.360 ;
        RECT 0.230 1.190 0.920 1.360 ;
        RECT 0.750 1.190 0.920 2.375 ;
        RECT 0.165 2.205 0.920 2.375 ;
        RECT 0.750 2.040 1.660 2.210 ;
        RECT 1.490 2.040 1.660 2.340 ;
        RECT 1.210 0.720 1.380 1.600 ;
        RECT 1.210 1.430 2.040 1.600 ;
        RECT 1.870 1.430 2.040 2.795 ;
        RECT 1.695 2.625 2.040 2.795 ;
        RECT 1.210 2.520 1.380 3.160 ;
        RECT 1.730 0.560 1.900 1.200 ;
        RECT 1.730 1.030 2.390 1.200 ;
        RECT 2.220 1.030 2.390 3.160 ;
        RECT 1.210 2.990 2.390 3.160 ;
        RECT 5.640 1.835 5.810 2.150 ;
        RECT 5.405 1.835 5.810 2.005 ;
        RECT 5.640 1.980 6.440 2.150 ;
        RECT 6.270 1.980 6.440 2.960 ;
        RECT 5.640 1.190 5.810 1.505 ;
        RECT 5.405 1.335 5.810 1.505 ;
        RECT 5.640 1.190 6.440 1.360 ;
        RECT 6.270 0.720 6.440 1.360 ;
  END 
END BUFTSHD5XHT

MACRO BUFTSHD4XHT
  CLASS  CORE ;
  FOREIGN BUFTSHD4XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.970 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 5.770 1.575 6.870 1.745 ;
        RECT 6.660 1.575 6.870 2.015 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.355 1.670 0.890 2.010 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.855 -0.300 1.155 0.895 ;
        RECT 3.335 -0.300 3.635 0.935 ;
        RECT 4.375 -0.300 4.675 0.935 ;
        RECT 5.415 -0.300 5.715 0.895 ;
        RECT 6.455 -0.300 6.755 1.235 ;
        RECT 0.000 -0.300 6.970 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 2.880 0.720 3.050 1.360 ;
        RECT 2.880 2.150 3.050 3.140 ;
        RECT 3.500 1.145 3.710 2.320 ;
        RECT 2.880 2.150 4.150 2.320 ;
        RECT 3.920 2.150 4.150 3.130 ;
        RECT 3.855 0.785 4.155 1.315 ;
        RECT 3.920 2.410 5.230 2.580 ;
        RECT 4.960 0.675 5.130 1.315 ;
        RECT 2.880 1.145 5.130 1.315 ;
        RECT 4.960 2.410 5.230 3.050 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.855 2.635 1.155 3.990 ;
        RECT 3.335 2.565 3.635 3.990 ;
        RECT 4.375 2.895 4.675 3.990 ;
        RECT 5.415 2.555 5.715 3.990 ;
        RECT 6.455 2.215 6.755 3.990 ;
        RECT 0.000 3.390 6.970 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.320 0.480 0.490 1.490 ;
        RECT 0.255 0.480 0.555 0.650 ;
        RECT 0.320 1.320 1.250 1.490 ;
        RECT 1.080 1.320 1.250 2.360 ;
        RECT 0.255 2.190 1.250 2.360 ;
        RECT 1.080 2.115 1.955 2.285 ;
        RECT 1.440 1.015 1.610 1.600 ;
        RECT 1.440 1.430 2.330 1.600 ;
        RECT 2.100 1.430 2.330 1.730 ;
        RECT 2.160 1.430 2.330 2.655 ;
        RECT 1.925 2.485 2.330 2.655 ;
        RECT 1.375 2.615 1.675 3.125 ;
        RECT 1.895 1.080 2.680 1.250 ;
        RECT 2.510 1.080 2.680 3.020 ;
        RECT 1.375 2.835 2.680 3.020 ;
        RECT 4.735 1.845 5.375 2.195 ;
        RECT 4.735 2.025 6.170 2.195 ;
        RECT 6.000 2.025 6.170 3.130 ;
        RECT 5.335 1.225 5.505 1.665 ;
        RECT 3.905 1.495 5.505 1.665 ;
        RECT 6.000 0.720 6.175 1.395 ;
        RECT 5.335 1.225 6.175 1.395 ;
  END 
END BUFTSHD4XHT

MACRO BUFTSHD3XHT
  CLASS  CORE ;
  FOREIGN BUFTSHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.740 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 4.945 1.585 5.385 1.995 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.520 2.020 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.945 ;
        RECT 2.520 -0.300 2.690 1.340 ;
        RECT 3.495 -0.300 3.795 1.275 ;
        RECT 4.565 -0.300 4.865 1.055 ;
        RECT 0.000 -0.300 5.740 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 2.970 1.260 3.210 1.610 ;
        RECT 2.970 1.455 4.250 1.610 ;
        RECT 3.040 0.720 3.210 2.815 ;
        RECT 3.040 1.455 3.215 2.430 ;
        RECT 3.040 2.260 4.315 2.430 ;
        RECT 4.080 0.720 4.250 1.625 ;
        RECT 3.040 1.455 4.250 1.625 ;
        RECT 4.015 2.260 4.315 2.770 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.705 2.605 1.005 3.990 ;
        RECT 2.520 2.400 2.690 3.990 ;
        RECT 3.495 2.805 3.795 3.990 ;
        RECT 4.565 2.635 4.865 3.990 ;
        RECT 0.000 3.390 5.740 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 1.085 1.295 ;
        RECT 0.915 1.125 1.085 2.370 ;
        RECT 0.105 2.200 1.085 2.370 ;
        RECT 1.320 1.680 1.490 2.695 ;
        RECT 1.800 1.060 1.970 1.850 ;
        RECT 1.320 1.680 1.970 1.850 ;
        RECT 1.320 2.395 2.320 2.695 ;
        RECT 1.280 0.710 1.450 1.220 ;
        RECT 1.280 0.710 2.340 0.880 ;
        RECT 2.170 0.710 2.340 2.215 ;
        RECT 1.805 2.045 2.340 2.215 ;
        RECT 3.545 1.815 4.185 2.080 ;
        RECT 3.545 1.910 4.715 2.080 ;
        RECT 4.545 1.910 4.715 2.345 ;
        RECT 4.545 2.175 5.320 2.345 ;
        RECT 5.150 2.175 5.320 3.155 ;
        RECT 4.430 1.235 4.600 1.730 ;
        RECT 5.150 0.720 5.320 1.405 ;
        RECT 4.430 1.235 5.320 1.405 ;
  END 
END BUFTSHD3XHT

MACRO BUFTSHD20XHT
  CLASS  CORE ;
  FOREIGN BUFTSHD20XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.910 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 17.290 1.575 20.465 1.745 ;
        RECT 20.125 1.575 20.465 1.950 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.610 0.485 2.015 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.055 ;
        RECT 1.705 -0.300 2.005 1.145 ;
        RECT 2.745 -0.300 3.045 1.145 ;
        RECT 6.325 -0.300 6.625 1.055 ;
        RECT 7.365 -0.300 7.665 1.055 ;
        RECT 8.405 -0.300 8.705 1.055 ;
        RECT 9.445 -0.300 9.745 1.055 ;
        RECT 10.485 -0.300 10.785 1.055 ;
        RECT 11.525 -0.300 11.825 1.055 ;
        RECT 12.565 -0.300 12.865 1.055 ;
        RECT 13.605 -0.300 13.905 1.055 ;
        RECT 14.645 -0.300 14.945 1.055 ;
        RECT 15.685 -0.300 15.985 1.055 ;
        RECT 17.375 -0.300 17.675 0.715 ;
        RECT 18.415 -0.300 18.715 0.715 ;
        RECT 19.455 -0.300 19.755 0.715 ;
        RECT 20.495 -0.300 20.795 1.055 ;
        RECT 0.000 -0.300 20.910 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 5.870 0.720 6.040 2.960 ;
        RECT 6.845 0.785 7.145 2.895 ;
        RECT 7.885 0.785 8.185 2.895 ;
        RECT 8.925 0.785 9.225 2.895 ;
        RECT 9.965 0.785 10.265 2.895 ;
        RECT 11.005 0.785 11.305 2.895 ;
        RECT 12.045 0.785 12.345 2.895 ;
        RECT 13.085 0.765 13.385 2.895 ;
        RECT 14.125 0.785 14.425 2.895 ;
        RECT 15.165 0.765 15.465 2.895 ;
        RECT 16.240 0.720 16.440 2.015 ;
        RECT 5.870 1.370 16.440 2.015 ;
        RECT 16.260 0.720 16.440 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.290 0.405 3.990 ;
        RECT 1.705 2.535 2.005 3.990 ;
        RECT 2.790 2.545 3.090 3.990 ;
        RECT 6.325 2.295 6.625 3.990 ;
        RECT 7.365 2.295 7.665 3.990 ;
        RECT 8.405 2.295 8.705 3.990 ;
        RECT 9.445 2.295 9.745 3.990 ;
        RECT 10.485 2.295 10.785 3.990 ;
        RECT 11.525 2.295 11.825 3.990 ;
        RECT 12.565 2.295 12.865 3.990 ;
        RECT 13.605 2.295 13.905 3.990 ;
        RECT 14.645 2.295 14.945 3.990 ;
        RECT 15.685 2.295 15.985 3.990 ;
        RECT 17.375 2.635 17.675 3.990 ;
        RECT 18.415 2.635 18.715 3.990 ;
        RECT 19.455 2.635 19.755 3.990 ;
        RECT 20.495 2.295 20.795 3.990 ;
        RECT 0.000 3.390 20.910 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.685 0.480 0.875 2.960 ;
        RECT 0.685 1.270 1.140 1.950 ;
        RECT 3.725 1.780 3.895 1.985 ;
        RECT 0.685 1.780 3.895 1.950 ;
        RECT 3.725 1.815 4.365 1.985 ;
        RECT 1.185 0.635 1.525 0.805 ;
        RECT 1.355 0.635 1.525 1.580 ;
        RECT 2.225 0.785 2.525 1.580 ;
        RECT 3.265 0.785 3.565 1.580 ;
        RECT 3.905 2.185 4.205 2.695 ;
        RECT 4.305 1.125 4.605 1.580 ;
        RECT 3.905 2.185 5.320 2.355 ;
        RECT 1.355 1.410 5.320 1.580 ;
        RECT 5.140 1.410 5.320 2.695 ;
        RECT 4.945 2.185 5.320 2.695 ;
        RECT 1.185 2.150 1.485 3.045 ;
        RECT 2.225 2.150 2.525 3.000 ;
        RECT 1.185 2.150 3.650 2.320 ;
        RECT 3.350 2.150 3.650 3.065 ;
        RECT 3.785 0.520 4.085 1.055 ;
        RECT 4.425 2.765 4.725 3.065 ;
        RECT 3.785 0.520 5.125 0.700 ;
        RECT 4.825 0.520 5.125 1.055 ;
        RECT 4.825 0.865 5.680 1.055 ;
        RECT 5.500 0.865 5.680 3.065 ;
        RECT 3.350 2.895 5.680 3.065 ;
        RECT 16.635 1.180 16.815 1.570 ;
        RECT 16.905 0.480 17.105 1.360 ;
        RECT 17.945 0.720 18.145 1.360 ;
        RECT 18.985 0.720 19.185 1.360 ;
        RECT 20.030 0.720 20.210 1.360 ;
        RECT 16.635 1.180 20.210 1.360 ;
        RECT 16.635 1.770 16.815 2.160 ;
        RECT 16.855 1.980 17.155 3.055 ;
        RECT 17.895 1.980 18.195 2.900 ;
        RECT 16.635 1.980 19.170 2.160 ;
        RECT 18.990 1.980 19.170 2.965 ;
        RECT 18.990 2.265 20.275 2.435 ;
        RECT 19.975 2.265 20.275 3.145 ;
  END 
END BUFTSHD20XHT

MACRO BUFTSHD12XHT
  CLASS  CORE ;
  FOREIGN BUFTSHD12XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.120 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 11.525 1.575 13.020 1.745 ;
        RECT 12.810 1.575 13.020 2.015 ;
    END
  END A
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.675 0.630 2.015 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.120 ;
        RECT 1.695 -0.300 1.995 1.120 ;
        RECT 4.660 -0.300 4.960 1.055 ;
        RECT 5.700 -0.300 6.000 1.055 ;
        RECT 6.740 -0.300 7.040 1.055 ;
        RECT 7.780 -0.300 8.080 1.055 ;
        RECT 8.820 -0.300 9.120 1.055 ;
        RECT 9.860 -0.300 10.160 1.055 ;
        RECT 11.640 -0.300 11.940 0.715 ;
        RECT 12.680 -0.300 12.980 1.055 ;
        RECT 0.000 -0.300 13.120 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER M1 ;
        RECT 4.205 0.720 4.375 2.960 ;
        RECT 5.180 0.785 5.480 2.895 ;
        RECT 5.180 1.300 6.520 2.005 ;
        RECT 6.220 0.785 6.520 2.895 ;
        RECT 7.260 0.785 7.560 2.895 ;
        RECT 7.260 1.300 8.600 2.005 ;
        RECT 8.300 0.785 8.600 2.895 ;
        RECT 9.340 0.765 9.640 2.895 ;
        RECT 4.205 1.365 10.615 1.980 ;
        RECT 10.445 0.715 10.615 2.960 ;
        RECT 10.435 1.365 10.615 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.545 0.955 3.990 ;
        RECT 1.695 2.885 1.995 3.990 ;
        RECT 4.660 2.295 4.960 3.990 ;
        RECT 5.700 2.295 6.000 3.990 ;
        RECT 6.740 2.295 7.040 3.990 ;
        RECT 7.780 2.295 8.080 3.990 ;
        RECT 8.820 2.295 9.120 3.990 ;
        RECT 9.860 2.295 10.160 3.990 ;
        RECT 11.640 2.635 11.940 3.990 ;
        RECT 12.680 2.295 12.980 3.990 ;
        RECT 0.000 3.390 13.120 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.995 0.340 1.495 ;
        RECT 0.105 2.195 0.405 2.705 ;
        RECT 0.170 1.325 1.060 1.495 ;
        RECT 0.880 1.325 1.060 2.365 ;
        RECT 0.105 2.195 1.060 2.365 ;
        RECT 0.880 1.840 2.505 2.010 ;
        RECT 1.240 1.430 3.620 1.600 ;
        RECT 1.240 0.655 1.410 1.600 ;
        RECT 2.790 1.060 2.960 2.480 ;
        RECT 1.240 1.400 2.960 1.600 ;
        RECT 2.780 1.430 2.980 2.480 ;
        RECT 2.780 1.430 3.620 1.730 ;
        RECT 1.240 2.190 1.410 2.830 ;
        RECT 1.240 2.190 2.440 2.360 ;
        RECT 2.270 2.190 2.440 2.830 ;
        RECT 2.205 0.520 2.505 1.055 ;
        RECT 2.205 0.520 3.545 0.700 ;
        RECT 3.310 2.180 3.480 2.830 ;
        RECT 2.270 2.660 3.480 2.830 ;
        RECT 3.245 0.520 3.545 1.120 ;
        RECT 3.245 0.940 4.005 1.120 ;
        RECT 3.835 0.940 4.005 2.350 ;
        RECT 3.310 2.180 4.005 2.350 ;
        RECT 10.810 1.770 10.990 2.160 ;
        RECT 11.185 1.980 11.355 2.960 ;
        RECT 10.810 1.980 12.400 2.160 ;
        RECT 12.220 1.980 12.400 2.960 ;
        RECT 10.810 1.195 10.990 1.570 ;
        RECT 11.170 0.720 11.370 1.375 ;
        RECT 12.220 0.720 12.400 1.375 ;
        RECT 10.810 1.195 12.400 1.375 ;
  END 
END BUFTSHD12XHT

MACRO BUFHDUXHT
  CLASS  CORE ;
  FOREIGN BUFHDUXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.550 2.020 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.685 -0.300 0.985 0.855 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.300 1.060 1.540 2.280 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.685 2.565 0.985 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 1.100 1.295 ;
        RECT 0.930 1.125 1.100 2.370 ;
        RECT 0.105 2.200 1.100 2.370 ;
  END 
END BUFHDUXHT

MACRO BUFHD7XHT
  CLASS  CORE ;
  FOREIGN BUFHD7XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.310 2.075 ;
        RECT 0.100 1.585 1.085 1.755 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.055 ;
        RECT 1.180 -0.300 1.480 1.055 ;
        RECT 2.245 -0.300 2.545 1.055 ;
        RECT 3.285 -0.300 3.585 1.055 ;
        RECT 4.325 -0.300 4.625 1.055 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.725 0.720 2.025 1.405 ;
        RECT 1.725 1.980 2.025 2.960 ;
        RECT 2.765 0.720 3.065 1.405 ;
        RECT 2.765 1.980 3.065 2.960 ;
        RECT 1.725 1.235 5.145 1.405 ;
        RECT 3.805 0.720 4.105 2.960 ;
        RECT 3.405 1.235 5.145 2.405 ;
        RECT 1.725 1.980 5.145 2.405 ;
        RECT 4.845 0.720 5.145 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.635 0.405 3.990 ;
        RECT 1.180 2.295 1.480 3.990 ;
        RECT 2.245 2.635 2.545 3.990 ;
        RECT 3.285 2.635 3.585 3.990 ;
        RECT 4.325 2.635 4.625 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 0.720 0.860 1.405 ;
        RECT 0.690 1.945 0.860 2.960 ;
        RECT 0.690 1.235 1.465 1.405 ;
        RECT 1.295 1.235 1.465 2.115 ;
        RECT 0.690 1.945 1.465 2.115 ;
        RECT 1.295 1.585 3.205 1.755 ;
  END 
END BUFHD7XHT

MACRO BUFHD2XHT
  CLASS  CORE ;
  FOREIGN BUFHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.595 0.555 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.490 -0.300 0.790 0.455 ;
        RECT 1.605 -0.300 1.905 1.055 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.150 0.720 1.320 1.415 ;
        RECT 1.085 1.980 1.385 2.905 ;
        RECT 1.150 1.235 1.950 1.415 ;
        RECT 1.740 1.235 1.950 2.150 ;
        RECT 1.085 1.980 1.950 2.150 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.490 3.125 0.790 3.990 ;
        RECT 1.605 2.635 1.905 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.195 0.405 2.745 ;
        RECT 0.105 1.125 0.905 1.295 ;
        RECT 0.735 1.125 0.905 2.365 ;
        RECT 0.105 2.195 0.905 2.365 ;
        RECT 0.735 1.595 1.375 1.765 ;
  END 
END BUFHD2XHT

MACRO BUFHD20XHT
  CLASS  CORE ;
  FOREIGN BUFHD20XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.350 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.410 1.605 0.820 1.950 ;
        RECT 0.410 1.605 2.595 1.775 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.255 -0.300 0.555 1.055 ;
        RECT 1.295 -0.300 1.595 1.055 ;
        RECT 2.335 -0.300 2.635 1.055 ;
        RECT 3.375 -0.300 3.675 1.055 ;
        RECT 4.415 -0.300 4.715 0.715 ;
        RECT 5.455 -0.300 5.755 0.715 ;
        RECT 6.495 -0.300 6.795 0.715 ;
        RECT 7.535 -0.300 7.835 0.715 ;
        RECT 8.575 -0.300 8.875 0.715 ;
        RECT 9.615 -0.300 9.915 0.715 ;
        RECT 10.655 -0.300 10.955 0.715 ;
        RECT 11.695 -0.300 11.995 0.715 ;
        RECT 12.735 -0.300 13.035 0.715 ;
        RECT 13.775 -0.300 14.075 1.055 ;
        RECT 0.000 -0.300 14.350 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.895 0.785 4.195 1.385 ;
        RECT 3.895 1.995 4.195 2.895 ;
        RECT 4.935 0.785 5.235 1.385 ;
        RECT 4.935 1.990 5.235 2.895 ;
        RECT 5.975 0.785 6.275 1.385 ;
        RECT 5.975 1.995 6.275 2.895 ;
        RECT 7.080 0.720 7.250 1.385 ;
        RECT 7.015 1.990 7.315 2.895 ;
        RECT 8.055 0.785 8.355 1.385 ;
        RECT 3.895 0.915 8.355 1.385 ;
        RECT 8.055 1.995 8.355 2.895 ;
        RECT 9.160 0.720 9.330 1.385 ;
        RECT 9.095 1.990 9.395 2.895 ;
        RECT 9.160 0.915 13.555 1.385 ;
        RECT 3.895 0.920 13.555 1.385 ;
        RECT 10.135 0.785 10.435 2.895 ;
        RECT 11.175 0.745 11.475 2.895 ;
        RECT 12.280 0.720 12.450 2.895 ;
        RECT 12.215 0.915 12.515 2.895 ;
        RECT 9.820 0.915 13.555 2.415 ;
        RECT 3.890 1.995 13.555 2.415 ;
        RECT 13.255 0.785 13.555 2.895 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.255 2.295 0.555 3.990 ;
        RECT 1.295 2.635 1.595 3.990 ;
        RECT 2.335 2.635 2.635 3.990 ;
        RECT 3.375 2.295 3.675 3.990 ;
        RECT 4.415 2.635 4.715 3.990 ;
        RECT 5.455 2.635 5.755 3.990 ;
        RECT 6.495 2.635 6.795 3.990 ;
        RECT 7.535 2.635 7.835 3.990 ;
        RECT 8.575 2.635 8.875 3.990 ;
        RECT 9.615 2.635 9.915 3.990 ;
        RECT 10.655 2.635 10.955 3.990 ;
        RECT 11.695 2.635 11.995 3.990 ;
        RECT 12.735 2.635 13.035 3.990 ;
        RECT 13.775 2.295 14.075 3.990 ;
        RECT 0.000 3.390 14.350 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.840 0.720 1.010 1.405 ;
        RECT 0.840 2.170 1.010 3.150 ;
        RECT 1.880 0.720 2.050 1.405 ;
        RECT 1.880 2.170 2.050 3.150 ;
        RECT 0.840 1.235 3.090 1.405 ;
        RECT 0.840 2.170 3.090 2.340 ;
        RECT 2.920 0.720 3.090 2.960 ;
        RECT 2.920 1.605 9.150 1.775 ;
  END 
END BUFHD20XHT

MACRO BUFHD8XHT
  CLASS  CORE ;
  FOREIGN BUFHD8XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.560 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.675 1.195 1.950 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.790 -0.300 1.090 1.055 ;
        RECT 1.830 -0.300 2.130 1.055 ;
        RECT 2.870 -0.300 3.170 1.055 ;
        RECT 3.910 -0.300 4.210 1.055 ;
        RECT 4.950 -0.300 5.250 1.055 ;
        RECT 5.990 -0.300 6.290 1.055 ;
        RECT 0.000 -0.300 6.560 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.355 2.075 5.775 2.315 ;
        RECT 2.350 2.230 5.775 2.315 ;
        RECT 2.350 0.785 2.650 1.450 ;
        RECT 2.355 1.980 2.650 2.895 ;
        RECT 2.350 2.230 2.650 2.895 ;
        RECT 3.390 0.785 3.690 1.450 ;
        RECT 3.390 1.980 3.690 2.895 ;
        RECT 4.430 0.785 4.730 1.450 ;
        RECT 4.430 1.980 4.730 2.895 ;
        RECT 2.350 1.235 5.770 1.450 ;
        RECT 4.760 1.235 5.770 2.315 ;
        RECT 5.470 0.785 5.770 2.895 ;
        RECT 2.355 1.980 5.770 2.315 ;
        RECT 5.470 2.075 5.775 2.895 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.790 2.495 1.090 3.990 ;
        RECT 1.830 2.165 2.130 3.990 ;
        RECT 2.870 2.635 3.170 3.990 ;
        RECT 3.910 2.635 4.210 3.990 ;
        RECT 4.950 2.635 5.250 3.990 ;
        RECT 5.990 2.295 6.290 3.990 ;
        RECT 0.000 3.390 6.560 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.335 0.620 0.505 1.495 ;
        RECT 0.335 2.130 0.505 2.770 ;
        RECT 0.335 1.325 1.545 1.495 ;
        RECT 0.335 2.130 1.545 2.300 ;
        RECT 1.375 0.620 1.545 2.965 ;
        RECT 1.375 1.630 4.515 1.800 ;
  END 
END BUFHD8XHT

MACRO BUFHDLXHT
  CLASS  CORE ;
  FOREIGN BUFHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 2.460 0.510 2.865 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.295 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.210 1.060 1.380 2.280 ;
        RECT 1.210 1.265 1.545 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.690 2.100 0.860 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 2.280 ;
        RECT 0.170 1.585 1.030 1.755 ;
        RECT 0.860 1.520 1.030 1.820 ;
  END 
END BUFHDLXHT

MACRO BUFHD8XSPGHT
  CLASS  CORE ;
  FOREIGN BUFHD8XSPGHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.560 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 1.165 0.345 1.705 3.080 ;
      LAYER V7 ;
        RECT 1.255 1.255 1.615 1.615 ;
      LAYER M7 ;
        RECT 0.730 1.245 1.870 1.625 ;
      LAYER V6 ;
        RECT 1.340 1.340 1.530 1.530 ;
      LAYER M4 ;
        RECT 0.925 0.825 1.125 1.640 ;
      LAYER V3 ;
        RECT 0.930 0.930 1.120 1.120 ;
      LAYER M3 ;
        RECT 0.360 0.925 1.220 1.125 ;
      LAYER V2 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M2 ;
        RECT 0.515 0.825 0.715 2.045 ;
      LAYER V1 ;
        RECT 0.520 1.750 0.710 1.940 ;
      LAYER M1 ;
        RECT 0.390 1.675 1.030 1.950 ;
      LAYER M6 ;
        RECT 1.335 0.805 1.535 1.925 ;
      LAYER V5 ;
        RECT 1.340 1.340 1.530 1.530 ;
      LAYER M5 ;
        RECT 0.730 1.335 1.705 1.535 ;
      LAYER V4 ;
        RECT 0.930 1.340 1.120 1.530 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.055 ;
        RECT 1.665 -0.300 1.965 1.055 ;
        RECT 2.705 -0.300 3.005 1.055 ;
        RECT 3.745 -0.300 4.045 1.055 ;
        RECT 4.785 -0.300 5.085 1.055 ;
        RECT 5.825 -0.300 6.125 1.055 ;
        RECT 0.000 -0.300 6.560 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 4.855 0.355 5.395 3.085 ;
      LAYER V7 ;
        RECT 4.945 2.075 5.305 2.435 ;
      LAYER M7 ;
        RECT 4.455 2.065 5.485 2.445 ;
      LAYER V6 ;
        RECT 5.030 2.160 5.220 2.350 ;
      LAYER M4 ;
        RECT 4.615 1.175 4.815 2.490 ;
      LAYER V3 ;
        RECT 4.620 1.340 4.810 1.530 ;
      LAYER M3 ;
        RECT 4.455 1.335 5.355 1.535 ;
      LAYER V2 ;
        RECT 5.030 1.340 5.220 1.530 ;
      LAYER M2 ;
        RECT 5.025 0.955 5.225 2.105 ;
      LAYER V1 ;
        RECT 5.030 1.750 5.220 1.940 ;
      LAYER M1 ;
        RECT 2.190 2.075 5.610 2.315 ;
        RECT 2.185 2.230 5.610 2.315 ;
        RECT 2.185 0.785 2.485 1.450 ;
        RECT 2.190 1.980 2.485 2.895 ;
        RECT 2.185 2.230 2.485 2.895 ;
        RECT 3.225 0.785 3.525 1.450 ;
        RECT 3.225 1.980 3.525 2.895 ;
        RECT 4.265 0.785 4.565 1.450 ;
        RECT 4.265 1.980 4.565 2.895 ;
        RECT 2.185 1.235 5.605 1.450 ;
        RECT 4.595 1.235 5.605 2.315 ;
        RECT 5.305 0.785 5.605 2.895 ;
        RECT 2.190 1.980 5.605 2.315 ;
        RECT 5.305 2.075 5.610 2.895 ;
      LAYER M6 ;
        RECT 5.025 0.805 5.225 2.715 ;
      LAYER V5 ;
        RECT 5.030 2.160 5.220 2.350 ;
      LAYER M5 ;
        RECT 4.455 2.155 5.485 2.355 ;
      LAYER V4 ;
        RECT 4.620 2.160 4.810 2.350 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.495 0.925 3.990 ;
        RECT 1.665 2.165 1.965 3.990 ;
        RECT 2.705 2.635 3.005 3.990 ;
        RECT 3.745 2.635 4.045 3.990 ;
        RECT 4.785 2.635 5.085 3.990 ;
        RECT 5.825 2.295 6.125 3.990 ;
        RECT 0.000 3.390 6.560 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.620 0.340 1.495 ;
        RECT 0.170 2.130 0.340 2.770 ;
        RECT 0.170 1.325 1.380 1.495 ;
        RECT 0.170 2.130 1.380 2.300 ;
        RECT 1.210 0.620 1.380 2.965 ;
        RECT 1.210 1.630 4.350 1.800 ;
  END 
END BUFHD8XSPGHT

MACRO BUFHD6XHT
  CLASS  CORE ;
  FOREIGN BUFHD6XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.310 2.015 ;
        RECT 0.100 1.585 1.085 1.755 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 0.935 ;
        RECT 1.175 -0.300 1.475 1.055 ;
        RECT 2.245 -0.300 2.545 1.055 ;
        RECT 3.285 -0.300 3.585 1.055 ;
        RECT 4.325 -0.300 4.625 1.055 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.725 0.720 2.025 1.405 ;
        RECT 1.725 1.980 2.025 2.960 ;
        RECT 1.725 1.235 4.105 1.405 ;
        RECT 1.725 1.980 3.070 2.415 ;
        RECT 2.765 0.720 3.065 1.405 ;
        RECT 3.065 1.235 3.070 2.960 ;
        RECT 2.765 1.980 3.070 2.960 ;
        RECT 3.065 1.235 4.105 2.400 ;
        RECT 1.725 1.980 4.105 2.400 ;
        RECT 3.805 0.720 4.105 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.325 0.405 3.990 ;
        RECT 1.175 2.295 1.475 3.990 ;
        RECT 2.245 2.635 2.545 3.990 ;
        RECT 3.285 2.635 3.585 3.990 ;
        RECT 4.325 2.295 4.625 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 1.060 0.860 1.405 ;
        RECT 0.690 1.945 0.860 2.620 ;
        RECT 0.690 1.235 1.465 1.405 ;
        RECT 1.295 1.235 1.465 2.115 ;
        RECT 0.690 1.945 1.465 2.115 ;
        RECT 1.295 1.585 2.865 1.755 ;
  END 
END BUFHD6XHT

MACRO BUFHD5XHT
  CLASS  CORE ;
  FOREIGN BUFHD5XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.510 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.310 2.015 ;
        RECT 0.100 1.585 1.085 1.755 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.005 ;
        RECT 1.205 -0.300 1.505 1.055 ;
        RECT 2.245 -0.300 2.545 1.055 ;
        RECT 3.285 -0.300 3.585 1.055 ;
        RECT 0.000 -0.300 4.510 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.725 0.720 2.025 1.405 ;
        RECT 1.725 1.980 2.025 2.960 ;
        RECT 1.725 1.235 4.105 1.405 ;
        RECT 2.765 0.720 3.065 2.960 ;
        RECT 2.765 1.235 3.070 2.960 ;
        RECT 2.765 1.235 4.105 2.440 ;
        RECT 1.725 1.980 4.105 2.440 ;
        RECT 3.805 0.720 4.105 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.225 0.405 3.990 ;
        RECT 1.205 2.295 1.505 3.990 ;
        RECT 2.245 2.635 2.545 3.990 ;
        RECT 3.285 2.635 3.585 3.990 ;
        RECT 0.000 3.390 4.510 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 1.060 0.860 1.405 ;
        RECT 0.690 1.945 0.860 2.620 ;
        RECT 0.690 1.235 1.465 1.405 ;
        RECT 1.295 1.235 1.465 2.115 ;
        RECT 0.690 1.945 1.465 2.115 ;
        RECT 1.295 1.585 2.525 1.755 ;
  END 
END BUFHD5XHT

MACRO BUFHD4XHT
  CLASS  CORE ;
  FOREIGN BUFHD4XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.370 0.510 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.005 ;
        RECT 1.205 -0.300 1.505 1.055 ;
        RECT 2.245 -0.300 2.545 1.055 ;
        RECT 3.285 -0.300 3.585 1.055 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.725 2.075 3.070 2.315 ;
        RECT 1.725 0.785 2.025 1.405 ;
        RECT 1.725 1.980 2.025 2.895 ;
        RECT 1.725 1.235 3.065 1.405 ;
        RECT 2.460 1.235 3.065 2.315 ;
        RECT 2.765 0.785 3.065 2.895 ;
        RECT 1.725 1.980 3.065 2.315 ;
        RECT 2.765 2.075 3.070 2.895 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.225 0.405 3.990 ;
        RECT 1.205 2.295 1.505 3.990 ;
        RECT 2.245 2.635 2.545 3.990 ;
        RECT 3.285 2.295 3.585 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 1.060 0.860 2.620 ;
        RECT 0.690 1.585 2.185 1.755 ;
  END 
END BUFHD4XHT

MACRO BUFHD3XHT
  CLASS  CORE ;
  FOREIGN BUFHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.730 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.770 -0.300 1.070 1.055 ;
        RECT 1.810 -0.300 2.110 1.055 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.355 0.720 1.525 1.450 ;
        RECT 1.295 1.980 1.590 2.895 ;
        RECT 1.290 2.230 1.590 2.895 ;
        RECT 1.355 1.235 2.630 1.450 ;
        RECT 2.295 1.235 2.630 2.360 ;
        RECT 1.295 1.980 2.630 2.360 ;
        RECT 2.320 0.785 2.630 2.360 ;
        RECT 1.290 2.230 2.630 2.360 ;
        RECT 2.330 0.785 2.630 2.895 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.770 2.635 1.070 3.990 ;
        RECT 1.810 2.635 2.110 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.315 0.720 0.485 1.405 ;
        RECT 0.315 2.195 0.485 3.175 ;
        RECT 0.315 1.235 1.110 1.405 ;
        RECT 0.940 1.235 1.110 2.365 ;
        RECT 0.315 2.195 1.110 2.365 ;
        RECT 0.940 1.630 2.095 1.800 ;
  END 
END BUFHD3XHT

MACRO BUFHD1XHT
  CLASS  CORE ;
  FOREIGN BUFHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.310 2.015 ;
        RECT 0.100 1.585 0.675 1.755 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.715 -0.300 1.015 1.055 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.300 0.720 1.470 2.960 ;
        RECT 1.300 1.235 1.540 1.640 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.750 2.570 0.920 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 1.405 ;
        RECT 0.170 1.235 1.120 1.405 ;
        RECT 0.950 1.235 1.120 2.365 ;
        RECT 0.105 2.195 1.120 2.365 ;
  END 
END BUFHD1XHT

MACRO BUFHD16XHT
  CLASS  CORE ;
  FOREIGN BUFHD16XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.480 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.445 1.605 0.795 1.950 ;
        RECT 0.445 1.605 1.905 1.775 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 -0.300 0.925 1.055 ;
        RECT 1.665 -0.300 1.965 1.055 ;
        RECT 2.705 -0.300 3.005 1.055 ;
        RECT 3.745 -0.300 4.045 0.715 ;
        RECT 4.785 -0.300 5.085 0.715 ;
        RECT 5.825 -0.300 6.125 0.715 ;
        RECT 6.865 -0.300 7.165 0.715 ;
        RECT 7.905 -0.300 8.205 0.715 ;
        RECT 8.945 -0.300 9.245 0.715 ;
        RECT 9.985 -0.300 10.285 0.715 ;
        RECT 11.025 -0.300 11.325 1.055 ;
        RECT 0.000 -0.300 11.480 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.225 0.785 3.525 1.360 ;
        RECT 3.225 1.995 3.525 2.895 ;
        RECT 4.265 0.785 4.565 1.360 ;
        RECT 4.265 1.990 4.565 2.895 ;
        RECT 5.305 0.785 5.605 1.360 ;
        RECT 5.305 1.995 5.605 2.895 ;
        RECT 6.410 0.720 6.580 1.360 ;
        RECT 6.345 1.990 6.645 2.895 ;
        RECT 7.385 0.785 7.685 1.360 ;
        RECT 7.385 1.995 7.685 2.895 ;
        RECT 8.490 0.720 8.660 1.360 ;
        RECT 8.425 1.990 8.725 2.895 ;
        RECT 3.225 0.915 10.805 1.360 ;
        RECT 9.465 0.785 9.765 2.895 ;
        RECT 9.150 0.915 10.805 2.435 ;
        RECT 3.220 1.995 10.805 2.435 ;
        RECT 10.505 0.745 10.805 2.895 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.635 0.925 3.990 ;
        RECT 1.665 2.635 1.965 3.990 ;
        RECT 2.705 2.295 3.005 3.990 ;
        RECT 3.745 2.635 4.045 3.990 ;
        RECT 4.785 2.635 5.085 3.990 ;
        RECT 5.825 2.635 6.125 3.990 ;
        RECT 6.865 2.635 7.165 3.990 ;
        RECT 7.905 2.635 8.205 3.990 ;
        RECT 8.945 2.635 9.245 3.990 ;
        RECT 9.985 2.635 10.285 3.990 ;
        RECT 11.025 2.295 11.325 3.990 ;
        RECT 0.000 3.390 11.480 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 0.720 0.340 1.405 ;
        RECT 0.170 2.170 0.340 3.150 ;
        RECT 1.210 0.720 1.380 1.405 ;
        RECT 1.210 2.170 1.380 3.150 ;
        RECT 0.170 1.235 2.420 1.405 ;
        RECT 0.170 2.170 2.420 2.340 ;
        RECT 2.250 0.720 2.420 2.960 ;
        RECT 2.250 1.585 8.785 1.755 ;
  END 
END BUFHD16XHT

MACRO BUFCLKHDUXHT
  CLASS  CORE ;
  FOREIGN BUFCLKHDUXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.615 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 0.845 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.270 1.060 1.440 2.280 ;
        RECT 1.270 1.060 1.470 1.605 ;
        RECT 1.270 1.265 1.540 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.545 0.955 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 1.090 1.295 ;
        RECT 0.920 1.125 1.090 2.365 ;
        RECT 0.105 2.195 1.090 2.365 ;
  END 
END BUFCLKHDUXHT

MACRO BUFCLKHDMXHT
  CLASS  CORE ;
  FOREIGN BUFCLKHDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.310 2.015 ;
        RECT 0.100 1.585 0.585 1.755 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.055 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.270 1.060 1.440 2.620 ;
        RECT 1.270 1.265 1.540 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.680 2.645 0.980 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 1.405 ;
        RECT 0.170 1.235 1.090 1.405 ;
        RECT 0.920 1.235 1.090 2.365 ;
        RECT 0.105 2.195 1.090 2.365 ;
  END 
END BUFCLKHDMXHT

MACRO BUFCLKHD8XHT
  CLASS  CORE ;
  FOREIGN BUFCLKHD8XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.650 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.245 -0.300 0.545 1.045 ;
        RECT 1.315 -0.300 1.615 1.045 ;
        RECT 2.355 -0.300 2.655 0.995 ;
        RECT 3.395 -0.300 3.695 0.995 ;
        RECT 4.435 -0.300 4.735 0.995 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.810 1.955 2.105 2.895 ;
        RECT 1.805 2.230 2.105 2.895 ;
        RECT 1.835 1.125 2.135 1.385 ;
        RECT 2.845 1.955 3.145 2.895 ;
        RECT 2.875 1.125 3.175 1.385 ;
        RECT 1.810 1.955 4.555 2.365 ;
        RECT 1.835 1.175 4.555 1.385 ;
        RECT 3.940 1.125 4.185 2.895 ;
        RECT 3.885 1.955 4.185 2.895 ;
        RECT 3.940 1.125 4.215 2.365 ;
        RECT 3.915 1.125 4.215 1.385 ;
        RECT 3.940 1.175 4.555 2.365 ;
        RECT 1.805 2.230 4.555 2.365 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.245 2.295 0.545 3.990 ;
        RECT 1.285 2.205 1.585 3.990 ;
        RECT 2.325 2.545 2.625 3.990 ;
        RECT 3.365 2.545 3.665 3.990 ;
        RECT 4.405 2.545 4.705 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.830 1.060 1.000 2.960 ;
        RECT 0.830 1.585 3.670 1.755 ;
  END 
END BUFCLKHD8XHT

MACRO AOI32HDMXHT
  CLASS  CORE ;
  FOREIGN AOI32HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.265 0.550 1.800 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.840 1.520 1.130 2.015 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 1.235 1.590 1.820 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.630 1.520 3.180 2.015 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.665 0.480 2.290 0.720 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.135 -0.300 0.435 1.025 ;
        RECT 2.710 -0.300 3.010 1.185 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.775 1.060 1.945 1.980 ;
        RECT 1.775 1.810 2.450 1.980 ;
        RECT 2.150 1.810 2.450 2.620 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.135 2.225 0.435 3.990 ;
        RECT 1.175 2.565 1.475 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.655 2.195 0.955 2.735 ;
        RECT 0.655 2.195 1.930 2.365 ;
        RECT 1.760 2.160 1.930 2.970 ;
        RECT 2.735 2.225 3.035 2.970 ;
        RECT 1.760 2.800 3.035 2.970 ;
  END 
END AOI32HDMXHT

MACRO BUFCLKHD3XHT
  CLASS  CORE ;
  FOREIGN BUFCLKHD3XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.625 0.700 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.770 -0.300 1.070 0.965 ;
        RECT 1.810 -0.300 2.110 0.965 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.355 1.030 1.525 1.405 ;
        RECT 1.295 1.980 1.590 2.895 ;
        RECT 1.290 2.230 1.590 2.895 ;
        RECT 1.355 1.225 2.630 1.405 ;
        RECT 1.295 1.980 2.630 2.315 ;
        RECT 1.955 1.225 2.630 2.315 ;
        RECT 1.290 2.230 2.630 2.315 ;
        RECT 2.330 1.115 2.630 2.895 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.770 2.635 1.070 3.990 ;
        RECT 1.810 2.635 2.110 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.285 1.040 0.455 1.445 ;
        RECT 0.285 2.195 0.455 2.835 ;
        RECT 0.285 1.265 1.085 1.445 ;
        RECT 0.915 1.265 1.085 2.365 ;
        RECT 0.285 2.195 1.085 2.365 ;
        RECT 0.915 1.585 1.755 1.755 ;
  END 
END BUFCLKHD3XHT

MACRO BUFCLKHD2XHT
  CLASS  CORE ;
  FOREIGN BUFCLKHD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.700 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.770 -0.300 1.070 1.035 ;
        RECT 1.870 -0.300 2.170 1.015 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.385 1.060 1.555 1.405 ;
        RECT 1.385 1.940 1.555 2.960 ;
        RECT 1.385 1.235 1.950 1.405 ;
        RECT 1.740 1.235 1.950 2.110 ;
        RECT 1.385 1.940 1.950 2.110 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.770 2.635 1.070 3.990 ;
        RECT 1.910 2.295 2.210 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.285 1.060 0.455 1.405 ;
        RECT 0.285 1.235 1.130 1.405 ;
        RECT 0.960 1.235 1.130 2.365 ;
        RECT 0.220 2.195 1.130 2.365 ;
        RECT 0.960 1.585 1.420 1.755 ;
  END 
END BUFCLKHD2XHT

MACRO BUFCLKHD1XHT
  CLASS  CORE ;
  FOREIGN BUFCLKHD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.675 0.585 2.015 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.105 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.240 1.060 1.410 2.960 ;
        RECT 1.240 1.265 1.430 2.960 ;
        RECT 1.240 1.265 1.540 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.635 0.955 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 1.495 ;
        RECT 0.170 1.325 1.060 1.495 ;
        RECT 0.890 1.325 1.060 2.365 ;
        RECT 0.100 2.195 1.060 2.365 ;
  END 
END BUFCLKHD1XHT

MACRO BUFCLKHD16XHT
  CLASS  CORE ;
  FOREIGN BUFCLKHD16XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.840 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.690 1.665 2.190 1.950 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.870 -0.300 1.170 1.045 ;
        RECT 1.910 -0.300 2.210 1.045 ;
        RECT 2.950 -0.300 3.250 1.045 ;
        RECT 3.990 -0.300 4.290 0.955 ;
        RECT 5.030 -0.300 5.330 0.955 ;
        RECT 6.070 -0.300 6.370 0.955 ;
        RECT 7.110 -0.300 7.410 0.955 ;
        RECT 8.150 -0.300 8.450 0.955 ;
        RECT 9.190 -0.300 9.490 1.035 ;
        RECT 0.000 -0.300 9.840 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.470 0.785 3.770 1.370 ;
        RECT 3.470 1.980 3.770 2.895 ;
        RECT 4.510 0.785 4.810 1.370 ;
        RECT 4.510 1.980 4.810 2.895 ;
        RECT 5.550 0.785 5.850 1.370 ;
        RECT 5.550 1.980 5.850 2.895 ;
        RECT 6.590 0.785 6.890 1.370 ;
        RECT 6.590 1.980 6.890 2.895 ;
        RECT 3.470 1.980 7.930 2.455 ;
        RECT 7.630 0.785 7.930 1.370 ;
        RECT 7.630 1.980 7.930 2.895 ;
        RECT 3.470 1.155 8.970 1.370 ;
        RECT 8.210 1.155 8.970 2.325 ;
        RECT 3.470 1.980 8.970 2.325 ;
        RECT 8.670 0.955 8.970 2.895 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.870 2.635 1.170 3.990 ;
        RECT 1.910 2.635 2.210 3.990 ;
        RECT 2.950 2.295 3.250 3.990 ;
        RECT 3.990 2.635 4.290 3.990 ;
        RECT 5.030 2.635 5.330 3.990 ;
        RECT 6.070 2.635 6.370 3.990 ;
        RECT 7.110 2.635 7.410 3.990 ;
        RECT 8.150 2.505 8.450 3.990 ;
        RECT 9.190 2.165 9.490 3.990 ;
        RECT 0.000 3.390 9.840 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.415 1.060 0.585 1.425 ;
        RECT 0.415 2.150 0.585 3.130 ;
        RECT 1.455 1.060 1.625 1.425 ;
        RECT 1.455 2.150 1.625 3.130 ;
        RECT 0.415 1.245 2.665 1.425 ;
        RECT 0.415 2.150 2.665 2.340 ;
        RECT 2.495 1.060 2.665 2.960 ;
        RECT 2.495 1.590 8.010 1.760 ;
  END 
END BUFCLKHD16XHT

MACRO BUFCLKHD14XHT
  CLASS  CORE ;
  FOREIGN BUFCLKHD14XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.200 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.690 1.595 1.755 1.950 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.310 -0.300 0.610 1.055 ;
        RECT 1.350 -0.300 1.650 1.055 ;
        RECT 2.390 -0.300 2.690 1.055 ;
        RECT 3.430 -0.300 3.730 1.055 ;
        RECT 4.470 -0.300 4.770 1.055 ;
        RECT 5.510 -0.300 5.810 1.055 ;
        RECT 6.550 -0.300 6.850 1.055 ;
        RECT 7.590 -0.300 7.890 1.055 ;
        RECT 0.000 -0.300 8.200 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.910 1.115 3.210 1.450 ;
        RECT 2.910 1.980 3.210 2.895 ;
        RECT 3.950 1.115 4.250 1.450 ;
        RECT 3.950 1.980 4.250 2.895 ;
        RECT 4.990 1.115 5.290 1.450 ;
        RECT 4.990 1.980 5.290 2.895 ;
        RECT 6.030 1.125 6.330 1.450 ;
        RECT 6.030 1.980 6.330 2.895 ;
        RECT 4.990 1.235 7.880 1.450 ;
        RECT 2.910 1.245 7.880 1.450 ;
        RECT 7.070 1.115 7.370 2.895 ;
        RECT 6.755 1.235 7.880 2.315 ;
        RECT 2.910 1.980 7.880 2.315 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.310 2.295 0.610 3.990 ;
        RECT 1.350 2.635 1.650 3.990 ;
        RECT 2.390 2.295 2.690 3.990 ;
        RECT 3.430 2.635 3.730 3.990 ;
        RECT 4.470 2.635 4.770 3.990 ;
        RECT 5.510 2.635 5.810 3.990 ;
        RECT 6.550 2.635 6.850 3.990 ;
        RECT 7.590 2.635 7.890 3.990 ;
        RECT 0.000 3.390 8.200 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.895 1.060 1.065 1.415 ;
        RECT 0.895 2.170 1.065 3.150 ;
        RECT 0.895 1.245 2.105 1.415 ;
        RECT 0.895 2.170 2.105 2.340 ;
        RECT 1.935 1.060 2.105 2.960 ;
        RECT 1.935 1.630 6.445 1.800 ;
  END 
END BUFCLKHD14XHT

MACRO BUFCLKHDLXHT
  CLASS  CORE ;
  FOREIGN BUFCLKHDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.640 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.310 2.015 ;
        RECT 0.100 1.585 0.585 1.755 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 -0.300 0.955 1.055 ;
        RECT 0.000 -0.300 1.640 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.270 1.060 1.440 2.620 ;
        RECT 1.270 1.265 1.540 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.655 2.545 0.955 3.990 ;
        RECT 0.000 3.390 1.640 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 1.060 0.340 1.405 ;
        RECT 0.170 1.235 1.090 1.405 ;
        RECT 0.920 1.235 1.090 2.365 ;
        RECT 0.105 2.195 1.090 2.365 ;
  END 
END BUFCLKHDLXHT

MACRO BUFCLKHD80XHT
  CLASS  CORE ;
  FOREIGN BUFCLKHD80XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 45.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.445 1.615 0.860 1.950 ;
        RECT 0.445 1.615 6.235 1.785 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.065 ;
        RECT 1.145 -0.300 1.445 1.065 ;
        RECT 2.185 -0.300 2.485 1.065 ;
        RECT 3.225 -0.300 3.525 1.065 ;
        RECT 4.265 -0.300 4.565 1.065 ;
        RECT 5.305 -0.300 5.605 1.055 ;
        RECT 6.345 -0.300 6.645 1.055 ;
        RECT 7.385 -0.300 7.685 1.055 ;
        RECT 8.425 -0.300 8.725 1.055 ;
        RECT 9.465 -0.300 9.765 1.055 ;
        RECT 10.535 -0.300 10.835 1.055 ;
        RECT 11.575 -0.300 11.875 0.715 ;
        RECT 12.615 -0.300 12.915 0.715 ;
        RECT 13.655 -0.300 13.955 0.715 ;
        RECT 14.695 -0.300 14.995 0.715 ;
        RECT 15.735 -0.300 16.035 0.715 ;
        RECT 16.775 -0.300 17.075 0.715 ;
        RECT 17.815 -0.300 18.115 0.715 ;
        RECT 18.855 -0.300 19.155 0.715 ;
        RECT 19.895 -0.300 20.195 0.715 ;
        RECT 20.935 -0.300 21.235 0.715 ;
        RECT 21.975 -0.300 22.275 0.715 ;
        RECT 23.015 -0.300 23.315 0.715 ;
        RECT 24.055 -0.300 24.355 0.715 ;
        RECT 25.095 -0.300 25.395 0.715 ;
        RECT 26.135 -0.300 26.435 0.715 ;
        RECT 27.175 -0.300 27.475 0.715 ;
        RECT 28.215 -0.300 28.515 0.715 ;
        RECT 29.255 -0.300 29.555 0.715 ;
        RECT 30.295 -0.300 30.595 0.715 ;
        RECT 31.335 -0.300 31.635 0.715 ;
        RECT 32.375 -0.300 32.675 0.715 ;
        RECT 33.415 -0.300 33.715 0.715 ;
        RECT 34.455 -0.300 34.755 0.715 ;
        RECT 35.495 -0.300 35.795 0.715 ;
        RECT 36.565 -0.300 36.865 0.715 ;
        RECT 0.000 -0.300 45.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 11.025 1.980 11.325 2.895 ;
        RECT 11.055 0.785 11.355 1.370 ;
        RECT 12.065 1.980 12.365 2.895 ;
        RECT 12.095 0.785 12.395 1.370 ;
        RECT 13.105 1.980 13.405 2.895 ;
        RECT 13.135 0.720 13.435 1.370 ;
        RECT 14.145 1.980 14.445 2.895 ;
        RECT 14.175 0.785 14.475 1.370 ;
        RECT 15.185 1.980 15.485 2.895 ;
        RECT 15.215 0.785 15.515 1.370 ;
        RECT 16.225 1.980 16.525 2.895 ;
        RECT 16.255 0.785 16.555 1.370 ;
        RECT 17.265 1.980 17.565 2.895 ;
        RECT 17.295 0.785 17.595 1.370 ;
        RECT 18.305 1.980 18.605 2.895 ;
        RECT 18.335 0.785 18.635 1.370 ;
        RECT 19.345 1.980 19.645 2.895 ;
        RECT 19.375 0.785 19.675 1.370 ;
        RECT 20.380 1.980 20.685 2.895 ;
        RECT 20.415 0.785 20.715 1.370 ;
        RECT 21.425 1.980 21.725 2.895 ;
        RECT 21.455 0.785 21.755 1.370 ;
        RECT 22.465 1.980 22.765 2.895 ;
        RECT 22.495 0.785 22.795 1.370 ;
        RECT 11.055 0.895 22.795 1.370 ;
        RECT 23.505 1.980 23.805 2.895 ;
        RECT 23.535 0.785 23.835 1.370 ;
        RECT 24.545 1.980 24.845 2.895 ;
        RECT 24.575 0.785 24.875 1.370 ;
        RECT 25.580 1.980 25.885 2.895 ;
        RECT 25.615 0.785 25.915 1.370 ;
        RECT 26.625 1.980 26.925 2.895 ;
        RECT 26.655 0.785 26.955 1.370 ;
        RECT 27.665 1.980 27.965 2.895 ;
        RECT 27.695 0.785 27.995 1.370 ;
        RECT 28.705 1.980 29.005 2.895 ;
        RECT 28.735 0.785 29.035 1.370 ;
        RECT 29.745 1.980 30.045 2.895 ;
        RECT 29.775 0.785 30.075 1.370 ;
        RECT 11.055 0.945 45.095 1.370 ;
        RECT 30.815 0.785 31.085 2.895 ;
        RECT 30.780 0.945 31.085 2.895 ;
        RECT 30.815 0.785 31.115 2.455 ;
        RECT 31.855 0.785 32.125 2.895 ;
        RECT 31.825 0.945 32.125 2.895 ;
        RECT 31.855 0.785 32.155 2.455 ;
        RECT 32.895 0.785 33.165 2.895 ;
        RECT 32.865 0.945 33.165 2.895 ;
        RECT 32.895 0.785 33.195 2.455 ;
        RECT 33.935 0.785 34.205 2.895 ;
        RECT 33.905 0.945 34.205 2.895 ;
        RECT 33.935 0.785 34.235 2.455 ;
        RECT 34.975 0.785 35.245 2.895 ;
        RECT 34.945 0.945 35.245 2.895 ;
        RECT 34.975 0.785 35.275 2.455 ;
        RECT 30.735 0.945 36.285 2.455 ;
        RECT 11.020 1.980 36.285 2.455 ;
        RECT 36.015 0.785 36.285 2.895 ;
        RECT 35.980 0.945 36.285 2.895 ;
        RECT 36.015 0.785 36.315 2.115 ;
        RECT 30.735 0.945 37.325 2.115 ;
        RECT 11.020 1.980 37.325 2.115 ;
        RECT 37.025 0.945 37.325 2.895 ;
        RECT 38.065 0.850 38.365 3.125 ;
        RECT 39.105 0.850 39.405 3.125 ;
        RECT 40.145 0.850 40.445 3.125 ;
        RECT 41.185 0.850 41.485 3.125 ;
        RECT 42.225 0.850 42.525 3.125 ;
        RECT 43.265 0.850 43.565 3.125 ;
        RECT 44.305 0.850 44.605 3.125 ;
        RECT 38.065 0.850 45.095 2.045 ;
        RECT 30.735 0.945 45.095 2.045 ;
        RECT 30.735 1.815 45.645 2.045 ;
        RECT 11.020 1.980 45.645 2.045 ;
        RECT 45.345 1.815 45.645 3.145 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 1.145 2.635 1.445 3.990 ;
        RECT 2.185 2.635 2.485 3.990 ;
        RECT 3.225 2.635 3.525 3.990 ;
        RECT 4.265 2.635 4.565 3.990 ;
        RECT 5.305 2.635 5.605 3.990 ;
        RECT 6.345 2.635 6.645 3.990 ;
        RECT 7.385 2.295 7.685 3.990 ;
        RECT 8.425 2.295 8.725 3.990 ;
        RECT 9.465 2.295 9.765 3.990 ;
        RECT 10.505 2.295 10.805 3.990 ;
        RECT 11.545 2.635 11.845 3.990 ;
        RECT 12.585 2.635 12.885 3.990 ;
        RECT 13.625 2.635 13.925 3.990 ;
        RECT 14.665 2.635 14.965 3.990 ;
        RECT 15.705 2.635 16.005 3.990 ;
        RECT 16.745 2.635 17.045 3.990 ;
        RECT 17.785 2.635 18.085 3.990 ;
        RECT 18.825 2.635 19.125 3.990 ;
        RECT 19.865 2.635 20.165 3.990 ;
        RECT 20.905 2.635 21.205 3.990 ;
        RECT 21.945 2.635 22.245 3.990 ;
        RECT 22.985 2.635 23.285 3.990 ;
        RECT 24.025 2.635 24.325 3.990 ;
        RECT 25.065 2.635 25.365 3.990 ;
        RECT 26.105 2.635 26.405 3.990 ;
        RECT 27.145 2.635 27.445 3.990 ;
        RECT 28.185 2.635 28.485 3.990 ;
        RECT 29.225 2.635 29.525 3.990 ;
        RECT 30.265 2.635 30.565 3.990 ;
        RECT 31.305 2.635 31.605 3.990 ;
        RECT 32.345 2.635 32.645 3.990 ;
        RECT 33.385 2.635 33.685 3.990 ;
        RECT 34.425 2.635 34.725 3.990 ;
        RECT 35.465 2.635 35.765 3.990 ;
        RECT 36.505 2.635 36.805 3.990 ;
        RECT 37.545 2.295 37.845 3.990 ;
        RECT 38.585 2.295 38.885 3.990 ;
        RECT 39.625 2.295 39.925 3.990 ;
        RECT 40.665 2.295 40.965 3.990 ;
        RECT 41.705 2.295 42.005 3.990 ;
        RECT 42.745 2.295 43.045 3.990 ;
        RECT 43.785 2.295 44.085 3.990 ;
        RECT 44.825 2.295 45.125 3.990 ;
        RECT 0.000 3.390 45.920 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.625 1.125 0.925 1.415 ;
        RECT 0.625 2.150 0.925 3.065 ;
        RECT 1.665 1.125 1.965 1.415 ;
        RECT 1.665 2.150 1.965 3.065 ;
        RECT 2.705 1.125 3.005 1.415 ;
        RECT 2.705 2.150 3.005 3.065 ;
        RECT 3.745 1.125 4.045 1.415 ;
        RECT 3.745 2.150 4.045 3.065 ;
        RECT 4.785 1.125 5.085 1.415 ;
        RECT 4.785 2.150 5.085 3.065 ;
        RECT 5.825 1.125 6.125 1.415 ;
        RECT 5.825 2.150 6.125 3.065 ;
        RECT 0.625 1.245 7.165 1.415 ;
        RECT 0.625 2.150 7.165 2.335 ;
        RECT 6.865 1.125 7.165 2.895 ;
        RECT 7.905 1.125 8.205 2.895 ;
        RECT 8.945 1.125 9.245 2.895 ;
        RECT 9.985 1.125 10.285 2.895 ;
        RECT 6.865 1.590 30.220 1.760 ;
  END 
END BUFCLKHD80XHT

MACRO BUFCLKHD7XHT
  CLASS  CORE ;
  FOREIGN BUFCLKHD7XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.425 1.645 1.175 1.950 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.175 -0.300 0.475 0.675 ;
        RECT 1.245 -0.300 1.545 0.945 ;
        RECT 2.335 -0.300 2.635 0.945 ;
        RECT 3.375 -0.300 3.675 0.945 ;
        RECT 4.415 -0.300 4.715 0.945 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.815 1.060 2.115 1.465 ;
        RECT 1.815 2.015 2.115 2.960 ;
        RECT 1.815 1.255 4.195 1.465 ;
        RECT 2.855 1.060 3.155 1.465 ;
        RECT 2.855 2.015 3.155 2.960 ;
        RECT 3.155 1.255 4.195 2.455 ;
        RECT 1.815 2.015 4.195 2.455 ;
        RECT 3.895 1.060 4.195 2.960 ;
        RECT 3.890 1.255 4.195 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.175 2.325 0.475 3.990 ;
        RECT 1.245 2.635 1.545 3.990 ;
        RECT 2.335 2.635 2.635 3.990 ;
        RECT 3.375 2.635 3.675 3.990 ;
        RECT 4.415 2.295 4.715 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.760 1.060 0.930 1.465 ;
        RECT 0.760 2.130 0.930 2.770 ;
        RECT 0.760 1.295 1.625 1.465 ;
        RECT 1.455 1.295 1.625 2.350 ;
        RECT 0.760 2.130 1.625 2.350 ;
        RECT 1.455 1.645 2.955 1.815 ;
  END 
END BUFCLKHD7XHT

MACRO BUFCLKHD5XHT
  CLASS  CORE ;
  FOREIGN BUFCLKHD5XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.590 0.310 2.025 ;
        RECT 0.100 1.590 1.030 1.760 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 0.855 ;
        RECT 1.175 -0.300 1.475 0.745 ;
        RECT 2.215 -0.300 2.515 0.745 ;
        RECT 3.255 -0.300 3.555 0.745 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.615 1.980 1.915 2.960 ;
        RECT 1.695 0.785 1.995 1.410 ;
        RECT 1.695 1.175 4.000 1.410 ;
        RECT 2.935 0.785 2.955 2.960 ;
        RECT 2.655 1.980 2.955 2.960 ;
        RECT 2.935 0.785 3.035 2.355 ;
        RECT 2.735 0.785 3.035 1.410 ;
        RECT 2.935 1.175 3.930 2.355 ;
        RECT 1.615 1.980 3.930 2.355 ;
        RECT 3.690 1.175 3.930 2.960 ;
        RECT 2.935 1.175 4.000 1.640 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.995 0.405 3.990 ;
        RECT 1.090 2.965 1.390 3.990 ;
        RECT 2.135 2.625 2.435 3.990 ;
        RECT 3.175 2.625 3.475 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 1.060 0.860 1.410 ;
        RECT 0.690 1.240 1.425 1.410 ;
        RECT 1.255 1.240 1.425 2.215 ;
        RECT 0.570 2.045 1.425 2.215 ;
        RECT 1.255 1.590 2.755 1.760 ;
  END 
END BUFCLKHD5XHT

MACRO BUFCLKHD40XHT
  CLASS  CORE ;
  FOREIGN BUFCLKHD40XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.190 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.440 1.665 0.825 1.950 ;
        RECT 0.440 1.665 3.460 1.835 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.105 ;
        RECT 1.145 -0.300 1.445 1.105 ;
        RECT 2.185 -0.300 2.485 1.105 ;
        RECT 3.225 -0.300 3.525 1.105 ;
        RECT 4.265 -0.300 4.565 1.105 ;
        RECT 5.305 -0.300 5.605 1.105 ;
        RECT 6.345 -0.300 6.645 0.715 ;
        RECT 7.385 -0.300 7.685 0.715 ;
        RECT 8.425 -0.300 8.725 0.715 ;
        RECT 9.465 -0.300 9.765 0.715 ;
        RECT 10.505 -0.300 10.805 0.715 ;
        RECT 11.545 -0.300 11.845 0.715 ;
        RECT 12.585 -0.300 12.885 0.715 ;
        RECT 13.625 -0.300 13.925 0.715 ;
        RECT 14.665 -0.300 14.965 0.715 ;
        RECT 15.705 -0.300 16.005 0.715 ;
        RECT 16.745 -0.300 17.045 0.715 ;
        RECT 17.785 -0.300 18.085 0.715 ;
        RECT 18.825 -0.300 19.125 0.715 ;
        RECT 0.000 -0.300 24.190 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.825 0.785 6.125 1.370 ;
        RECT 5.825 1.980 6.125 2.895 ;
        RECT 6.865 0.785 7.165 1.370 ;
        RECT 6.865 1.980 7.165 2.895 ;
        RECT 7.905 0.785 8.205 1.370 ;
        RECT 7.905 1.980 8.205 2.895 ;
        RECT 8.945 0.785 9.245 1.370 ;
        RECT 8.945 1.980 9.245 2.895 ;
        RECT 9.985 0.785 10.285 1.370 ;
        RECT 9.985 1.980 10.285 2.895 ;
        RECT 11.025 0.785 11.325 1.370 ;
        RECT 11.025 1.980 11.325 2.895 ;
        RECT 12.065 0.785 12.365 1.370 ;
        RECT 12.065 1.980 12.365 2.895 ;
        RECT 13.105 0.785 13.405 1.370 ;
        RECT 13.105 1.980 13.405 2.895 ;
        RECT 14.145 0.785 14.445 1.370 ;
        RECT 14.145 1.980 14.445 2.895 ;
        RECT 15.185 0.785 15.485 1.370 ;
        RECT 15.180 1.980 15.485 2.895 ;
        RECT 5.825 0.895 16.525 1.370 ;
        RECT 5.825 0.965 22.765 1.370 ;
        RECT 16.195 0.895 16.525 2.450 ;
        RECT 5.825 1.980 16.525 2.450 ;
        RECT 16.225 0.785 16.525 2.895 ;
        RECT 17.265 0.785 17.565 2.895 ;
        RECT 18.305 0.545 18.605 2.895 ;
        RECT 19.345 0.965 19.645 2.895 ;
        RECT 16.195 0.965 22.765 2.385 ;
        RECT 20.380 0.965 20.685 2.685 ;
        RECT 20.385 0.895 20.685 3.105 ;
        RECT 21.425 0.895 21.725 3.105 ;
        RECT 20.385 0.895 22.765 2.385 ;
        RECT 5.825 1.980 22.765 2.385 ;
        RECT 22.465 0.895 22.765 3.105 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 1.145 2.635 1.445 3.990 ;
        RECT 2.185 2.635 2.485 3.990 ;
        RECT 3.225 2.635 3.525 3.990 ;
        RECT 4.265 2.295 4.565 3.990 ;
        RECT 5.305 2.295 5.605 3.990 ;
        RECT 6.345 2.635 6.645 3.990 ;
        RECT 7.385 2.635 7.685 3.990 ;
        RECT 8.425 2.635 8.725 3.990 ;
        RECT 9.465 2.635 9.765 3.990 ;
        RECT 10.505 2.635 10.805 3.990 ;
        RECT 11.545 2.635 11.845 3.990 ;
        RECT 12.585 2.635 12.885 3.990 ;
        RECT 13.625 2.635 13.925 3.990 ;
        RECT 14.665 2.635 14.965 3.990 ;
        RECT 15.705 2.635 16.005 3.990 ;
        RECT 16.745 2.635 17.045 3.990 ;
        RECT 17.785 2.635 18.085 3.990 ;
        RECT 18.825 2.635 19.125 3.990 ;
        RECT 19.865 2.635 20.165 3.990 ;
        RECT 20.905 2.635 21.205 3.990 ;
        RECT 21.945 2.635 22.245 3.990 ;
        RECT 22.985 0.935 23.285 3.990 ;
        RECT 0.000 3.390 24.190 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.625 1.125 0.925 1.465 ;
        RECT 0.625 2.150 0.925 3.065 ;
        RECT 1.665 1.125 1.965 1.465 ;
        RECT 1.665 2.150 1.965 3.065 ;
        RECT 2.705 1.125 3.005 1.465 ;
        RECT 2.705 2.150 3.005 3.065 ;
        RECT 0.625 1.295 4.045 1.465 ;
        RECT 0.625 2.150 4.045 2.340 ;
        RECT 3.745 1.125 4.045 2.895 ;
        RECT 4.785 1.125 5.085 2.895 ;
        RECT 3.745 1.590 15.895 1.760 ;
  END 
END BUFCLKHD40XHT

MACRO BUFCLKHD30XHT
  CLASS  CORE ;
  FOREIGN BUFCLKHD30XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.450 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.445 1.640 0.805 1.950 ;
        RECT 0.445 1.640 2.450 1.810 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.105 ;
        RECT 1.145 -0.300 1.445 1.105 ;
        RECT 2.185 -0.300 2.485 1.105 ;
        RECT 3.225 -0.300 3.525 1.105 ;
        RECT 4.265 -0.300 4.565 1.105 ;
        RECT 5.305 -0.300 5.605 0.715 ;
        RECT 6.345 -0.300 6.645 0.715 ;
        RECT 7.385 -0.300 7.685 0.715 ;
        RECT 8.425 -0.300 8.725 0.715 ;
        RECT 9.465 -0.300 9.765 0.715 ;
        RECT 10.505 -0.300 10.805 0.715 ;
        RECT 11.545 -0.300 11.845 0.715 ;
        RECT 12.585 -0.300 12.885 0.715 ;
        RECT 13.625 -0.300 13.925 0.715 ;
        RECT 0.000 -0.300 18.450 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.785 0.785 5.085 1.365 ;
        RECT 4.785 1.980 5.085 2.895 ;
        RECT 5.825 0.785 6.125 1.365 ;
        RECT 5.825 1.980 6.125 2.895 ;
        RECT 6.865 0.785 7.165 1.365 ;
        RECT 6.865 1.980 7.165 2.895 ;
        RECT 7.905 0.785 8.205 1.365 ;
        RECT 7.905 1.980 8.205 2.895 ;
        RECT 8.945 0.785 9.245 1.365 ;
        RECT 8.945 1.980 9.245 2.895 ;
        RECT 9.985 0.785 10.285 1.365 ;
        RECT 9.985 1.980 10.285 2.895 ;
        RECT 11.025 0.785 11.325 1.365 ;
        RECT 11.025 1.980 11.325 2.895 ;
        RECT 12.065 0.785 12.365 1.365 ;
        RECT 12.065 1.980 12.365 2.895 ;
        RECT 4.785 0.895 13.405 1.365 ;
        RECT 4.785 1.980 13.405 2.455 ;
        RECT 13.105 0.785 13.405 1.365 ;
        RECT 4.785 0.965 17.610 1.365 ;
        RECT 13.335 0.785 13.405 2.895 ;
        RECT 13.105 1.980 13.405 2.895 ;
        RECT 13.335 0.965 17.610 2.385 ;
        RECT 14.145 0.605 14.445 2.895 ;
        RECT 14.140 0.965 14.445 2.895 ;
        RECT 15.215 0.750 15.515 3.125 ;
        RECT 16.255 0.750 16.555 3.125 ;
        RECT 14.145 0.750 17.610 2.385 ;
        RECT 4.785 1.980 17.610 2.385 ;
        RECT 17.295 0.750 17.595 3.125 ;
        RECT 17.295 0.750 17.610 2.455 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.215 0.405 3.990 ;
        RECT 1.145 2.555 1.445 3.990 ;
        RECT 2.185 2.555 2.485 3.990 ;
        RECT 3.225 2.225 3.525 3.990 ;
        RECT 4.265 2.225 4.565 3.990 ;
        RECT 5.305 2.635 5.605 3.990 ;
        RECT 6.345 2.635 6.645 3.990 ;
        RECT 7.385 2.635 7.685 3.990 ;
        RECT 8.425 2.635 8.725 3.990 ;
        RECT 9.465 2.635 9.765 3.990 ;
        RECT 10.505 2.635 10.805 3.990 ;
        RECT 11.545 2.635 11.845 3.990 ;
        RECT 12.585 2.635 12.885 3.990 ;
        RECT 13.625 2.635 13.925 3.990 ;
        RECT 14.665 2.635 14.965 3.990 ;
        RECT 15.735 2.635 16.035 3.990 ;
        RECT 16.775 2.635 17.075 3.990 ;
        RECT 17.845 2.295 18.145 3.990 ;
        RECT 0.000 3.390 18.450 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 1.030 0.860 1.455 ;
        RECT 0.690 2.130 0.860 3.110 ;
        RECT 1.730 1.030 1.900 1.455 ;
        RECT 1.730 2.130 1.900 3.110 ;
        RECT 0.690 1.285 2.940 1.455 ;
        RECT 0.690 2.130 2.940 2.300 ;
        RECT 2.770 1.030 2.940 2.960 ;
        RECT 3.810 1.030 3.980 2.960 ;
        RECT 2.770 1.585 13.125 1.755 ;
  END 
END BUFCLKHD30XHT

MACRO BUFCLKHD20XHT
  CLASS  CORE ;
  FOREIGN BUFCLKHD20XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.940 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.635 1.645 2.040 1.950 ;
        RECT 0.635 1.645 2.980 1.815 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.335 -0.300 1.635 0.895 ;
        RECT 2.375 -0.300 2.675 0.895 ;
        RECT 3.415 -0.300 3.715 0.895 ;
        RECT 4.455 -0.300 4.755 0.715 ;
        RECT 5.495 -0.300 5.795 0.715 ;
        RECT 6.535 -0.300 6.835 0.715 ;
        RECT 7.575 -0.300 7.875 0.715 ;
        RECT 8.615 -0.300 8.915 0.715 ;
        RECT 9.655 -0.300 9.955 0.720 ;
        RECT 10.700 -0.300 11.000 0.715 ;
        RECT 0.000 -0.300 13.940 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.935 0.985 13.105 1.025 ;
        RECT 3.935 0.785 4.235 1.370 ;
        RECT 4.455 1.980 4.755 2.895 ;
        RECT 4.975 0.785 5.275 1.370 ;
        RECT 5.495 1.980 5.795 2.895 ;
        RECT 6.015 0.785 6.315 1.370 ;
        RECT 6.535 1.980 6.835 2.895 ;
        RECT 7.055 0.785 7.355 1.370 ;
        RECT 7.575 1.980 7.875 2.895 ;
        RECT 8.095 0.785 8.395 1.370 ;
        RECT 8.615 1.980 8.915 2.895 ;
        RECT 9.135 0.785 9.435 1.370 ;
        RECT 9.655 1.980 9.955 2.895 ;
        RECT 10.175 0.765 10.475 1.370 ;
        RECT 9.135 0.920 10.475 1.370 ;
        RECT 9.135 0.965 12.065 1.370 ;
        RECT 3.935 0.985 12.065 1.370 ;
        RECT 10.620 0.965 10.995 2.450 ;
        RECT 4.455 1.980 10.995 2.450 ;
        RECT 10.695 0.965 10.995 2.895 ;
        RECT 10.620 0.965 12.065 2.385 ;
        RECT 11.225 0.570 12.065 2.385 ;
        RECT 4.455 1.980 12.065 2.385 ;
        RECT 11.765 0.570 12.065 3.025 ;
        RECT 12.805 0.570 13.100 3.025 ;
        RECT 11.225 0.570 13.100 1.025 ;
        RECT 12.805 0.855 13.105 3.025 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.815 2.575 1.115 3.990 ;
        RECT 1.855 2.575 2.155 3.990 ;
        RECT 2.895 2.575 3.195 3.990 ;
        RECT 3.935 2.235 4.235 3.990 ;
        RECT 4.975 2.635 5.275 3.990 ;
        RECT 6.015 2.635 6.315 3.990 ;
        RECT 7.055 2.635 7.355 3.990 ;
        RECT 8.095 2.635 8.395 3.990 ;
        RECT 9.135 2.635 9.435 3.990 ;
        RECT 10.175 2.635 10.475 3.990 ;
        RECT 11.215 2.635 11.515 3.990 ;
        RECT 12.285 1.275 12.585 3.990 ;
        RECT 13.355 2.295 13.655 3.990 ;
        RECT 0.000 3.390 13.940 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.295 2.150 0.595 3.065 ;
        RECT 0.815 1.115 1.115 1.445 ;
        RECT 1.335 2.150 1.635 3.065 ;
        RECT 1.855 1.115 2.155 1.445 ;
        RECT 2.375 2.150 2.675 3.065 ;
        RECT 2.895 1.115 3.195 1.445 ;
        RECT 0.815 1.160 3.715 1.445 ;
        RECT 0.295 2.150 3.715 2.365 ;
        RECT 3.415 1.160 3.715 2.895 ;
        RECT 3.415 1.590 10.420 1.760 ;
  END 
END BUFCLKHD20XHT

MACRO AOI22B2HD1XHT
  CLASS  CORE ;
  FOREIGN AOI22B2HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.540 0.470 2.015 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.360 1.265 3.590 1.820 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.650 1.520 3.180 2.015 ;
    END
  END D
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.810 2.685 1.215 3.180 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.295 ;
        RECT 1.255 -0.300 1.895 1.295 ;
        RECT 3.260 -0.300 3.560 1.055 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.765 1.935 1.935 2.960 ;
        RECT 2.150 0.855 2.455 1.190 ;
        RECT 2.285 0.720 2.455 2.105 ;
        RECT 1.765 1.935 2.455 2.105 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.315 0.405 3.990 ;
        RECT 2.740 2.635 3.040 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.705 1.060 0.875 1.755 ;
        RECT 1.115 1.585 1.285 2.280 ;
        RECT 0.705 1.585 2.105 1.755 ;
        RECT 2.220 2.285 2.520 3.145 ;
        RECT 2.220 2.285 3.560 2.455 ;
        RECT 3.260 2.285 3.560 3.145 ;
  END 
END AOI22B2HD1XHT

MACRO AOI222HDLXHT
  CLASS  CORE ;
  FOREIGN AOI222HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.520 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 1.585 1.330 1.955 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.035 1.595 2.575 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.540 0.510 2.065 0.925 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.765 1.585 3.245 1.950 ;
    END
  END E
  PIN F
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.775 1.530 4.010 2.215 ;
    END
  END F
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.295 ;
        RECT 2.485 -0.300 2.785 0.940 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.425 0.920 3.475 2.640 ;
        RECT 3.175 2.130 3.475 2.640 ;
        RECT 3.425 0.920 3.595 2.305 ;
        RECT 3.175 2.130 3.595 2.305 ;
        RECT 3.315 0.920 3.675 1.295 ;
        RECT 1.140 1.125 3.900 1.295 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.355 0.405 3.990 ;
        RECT 1.175 2.830 1.475 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 2.195 0.860 2.835 ;
        RECT 0.690 2.480 2.435 2.650 ;
        RECT 1.615 2.130 2.890 2.300 ;
        RECT 2.720 2.130 2.890 2.990 ;
        RECT 3.760 2.630 3.930 2.990 ;
        RECT 2.720 2.820 3.930 2.990 ;
  END 
END AOI222HDLXHT

MACRO AOI222HD2XHT
  CLASS  CORE ;
  FOREIGN AOI222HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.150 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.520 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.830 1.590 1.305 1.960 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.065 1.595 2.625 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.630 0.510 2.075 0.925 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.015 0.510 3.655 0.940 ;
    END
  END E
  PIN F
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.630 1.530 4.000 2.015 ;
    END
  END F
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.295 ;
        RECT 2.535 -0.300 2.835 0.945 ;
        RECT 4.770 -0.300 4.940 1.120 ;
        RECT 5.745 -0.300 6.045 1.055 ;
        RECT 0.000 -0.300 6.150 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.015 2.045 5.460 2.425 ;
        RECT 5.290 0.720 5.545 1.360 ;
        RECT 5.375 0.720 5.460 2.960 ;
        RECT 5.290 2.045 5.460 2.960 ;
        RECT 5.375 0.720 5.545 2.215 ;
        RECT 5.015 2.045 5.545 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.355 0.405 3.990 ;
        RECT 1.175 2.830 1.475 3.990 ;
        RECT 4.705 2.975 5.005 3.990 ;
        RECT 5.745 2.295 6.045 3.990 ;
        RECT 0.000 3.390 6.150 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 2.195 0.860 2.835 ;
        RECT 0.690 2.480 2.470 2.650 ;
        RECT 1.635 2.130 2.925 2.300 ;
        RECT 2.755 2.130 2.925 2.970 ;
        RECT 3.795 2.290 3.965 2.970 ;
        RECT 2.755 2.800 3.965 2.970 ;
        RECT 3.275 1.125 3.445 2.620 ;
        RECT 3.835 0.615 4.005 1.295 ;
        RECT 1.190 1.125 4.005 1.295 ;
        RECT 3.835 0.615 4.590 0.785 ;
        RECT 4.220 1.060 4.505 1.360 ;
        RECT 4.310 1.060 4.480 2.280 ;
        RECT 4.310 1.060 4.505 1.820 ;
        RECT 4.310 1.520 5.175 1.820 ;
  END 
END AOI222HD2XHT

MACRO AOI222HD1XHT
  CLASS  CORE ;
  FOREIGN AOI222HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.740 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.540 0.520 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.735 1.590 1.195 1.955 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.085 1.595 2.685 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.640 0.510 2.030 0.925 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.075 0.510 3.655 0.940 ;
    END
  END E
  PIN F
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.665 1.530 4.005 2.020 ;
    END
  END F
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.295 ;
        RECT 2.555 -0.300 2.855 0.915 ;
        RECT 4.870 -0.300 5.040 1.120 ;
        RECT 0.000 -0.300 5.740 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 5.395 0.720 5.640 1.360 ;
        RECT 5.470 0.720 5.640 2.960 ;
        RECT 5.395 1.980 5.640 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.355 0.405 3.990 ;
        RECT 1.175 2.830 1.475 3.990 ;
        RECT 4.810 2.165 5.110 3.990 ;
        RECT 0.000 3.390 5.740 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 2.195 0.860 2.835 ;
        RECT 0.690 2.480 2.505 2.650 ;
        RECT 1.685 2.130 2.960 2.300 ;
        RECT 2.790 2.130 2.960 2.970 ;
        RECT 3.830 2.290 4.000 2.970 ;
        RECT 2.790 2.800 4.000 2.970 ;
        RECT 3.310 1.125 3.480 2.620 ;
        RECT 3.845 0.755 4.015 1.295 ;
        RECT 1.180 1.125 4.015 1.295 ;
        RECT 3.845 0.755 4.690 0.925 ;
        RECT 4.225 1.125 4.525 1.295 ;
        RECT 4.340 1.125 4.510 2.280 ;
        RECT 4.340 1.125 4.525 1.755 ;
        RECT 4.340 1.585 5.290 1.755 ;
  END 
END AOI222HD1XHT

MACRO AOI221HDMXHT
  CLASS  CORE ;
  FOREIGN AOI221HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.520 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 1.590 1.195 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.355 1.595 2.915 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.650 1.600 2.135 1.950 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.045 0.510 3.655 0.875 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.205 ;
        RECT 2.565 -0.300 2.865 0.945 ;
        RECT 4.290 -0.300 4.590 1.145 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.935 0.810 5.230 1.360 ;
        RECT 5.060 0.810 5.230 2.215 ;
        RECT 4.840 2.045 5.230 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 1.145 2.975 1.445 3.990 ;
        RECT 4.355 2.310 4.525 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 2.565 0.860 3.205 ;
        RECT 0.690 2.565 2.410 2.735 ;
        RECT 2.240 2.565 2.410 3.205 ;
        RECT 1.655 2.215 2.930 2.385 ;
        RECT 2.760 2.215 2.930 3.195 ;
        RECT 3.280 1.125 3.450 2.960 ;
        RECT 1.110 1.125 3.515 1.295 ;
        RECT 3.280 2.535 4.155 2.705 ;
        RECT 3.985 2.470 4.155 2.770 ;
        RECT 3.785 1.060 3.970 2.280 ;
        RECT 3.785 1.585 4.820 1.755 ;
  END 
END AOI221HDMXHT

MACRO AOI221HDLXHT
  CLASS  CORE ;
  FOREIGN AOI221HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.520 2.020 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 1.615 1.195 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.955 0.510 2.485 0.900 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.650 1.640 2.135 1.950 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.495 1.595 2.855 1.955 ;
        RECT 2.495 1.595 3.175 1.765 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.205 ;
        RECT 2.665 -0.300 2.965 0.990 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.145 1.125 1.785 1.340 ;
        RECT 3.270 1.125 3.590 1.340 ;
        RECT 1.145 1.170 3.590 1.340 ;
        RECT 3.390 1.125 3.590 2.960 ;
        RECT 3.230 2.045 3.590 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 1.145 2.975 1.445 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 2.565 0.860 3.205 ;
        RECT 0.690 2.565 2.410 2.735 ;
        RECT 2.240 2.565 2.410 3.205 ;
        RECT 1.655 2.215 2.930 2.385 ;
        RECT 2.760 2.215 2.930 3.195 ;
  END 
END AOI221HDLXHT

MACRO BUFHD12XHT
  CLASS  CORE ;
  FOREIGN BUFHD12XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.020 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.445 1.585 0.790 1.950 ;
        RECT 0.445 1.585 1.485 1.755 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.065 ;
        RECT 1.145 -0.300 1.445 1.055 ;
        RECT 2.185 -0.300 2.485 1.055 ;
        RECT 3.225 -0.300 3.525 0.715 ;
        RECT 4.265 -0.300 4.565 0.715 ;
        RECT 5.305 -0.300 5.605 0.725 ;
        RECT 6.345 -0.300 6.645 0.715 ;
        RECT 7.385 -0.300 7.685 0.725 ;
        RECT 8.425 -0.300 8.725 1.055 ;
        RECT 0.000 -0.300 9.020 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.700 2.075 8.210 2.405 ;
        RECT 2.705 0.785 3.005 1.365 ;
        RECT 2.705 1.980 3.005 2.895 ;
        RECT 3.745 0.785 4.045 1.365 ;
        RECT 3.745 1.980 4.045 2.895 ;
        RECT 4.785 0.785 5.085 1.365 ;
        RECT 4.785 1.980 5.085 2.895 ;
        RECT 5.825 0.785 6.125 1.365 ;
        RECT 5.825 1.980 6.125 2.895 ;
        RECT 2.705 0.940 8.205 1.365 ;
        RECT 6.865 0.785 7.165 2.895 ;
        RECT 6.835 0.940 8.205 2.405 ;
        RECT 7.905 0.785 8.205 2.895 ;
        RECT 2.700 1.980 8.205 2.405 ;
        RECT 7.905 2.075 8.210 2.895 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 1.145 2.635 1.445 3.990 ;
        RECT 2.185 2.295 2.485 3.990 ;
        RECT 3.225 2.635 3.525 3.990 ;
        RECT 4.265 2.635 4.565 3.990 ;
        RECT 5.305 2.635 5.605 3.990 ;
        RECT 6.345 2.635 6.645 3.990 ;
        RECT 7.385 2.635 7.685 3.990 ;
        RECT 8.425 2.295 8.725 3.990 ;
        RECT 0.000 3.390 9.020 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 0.720 0.860 1.405 ;
        RECT 0.690 2.130 0.860 3.110 ;
        RECT 0.690 1.235 1.900 1.405 ;
        RECT 0.690 2.130 1.900 2.300 ;
        RECT 1.730 0.720 1.900 2.960 ;
        RECT 1.730 1.585 6.565 1.755 ;
  END 
END BUFHD12XHT

MACRO AOI21B2HDLXHT
  CLASS  CORE ;
  FOREIGN AOI21B2HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.495 2.860 2.035 3.180 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.310 2.015 ;
        RECT 0.100 1.520 0.485 1.820 ;
    END
  END C
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.265 2.360 1.820 ;
        RECT 1.925 1.520 2.360 1.820 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.295 ;
        RECT 1.175 -0.300 1.475 0.745 ;
        RECT 2.055 -0.300 2.355 0.745 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 2.085 0.835 2.425 ;
        RECT 0.665 1.060 0.835 2.425 ;
        RECT 0.105 2.255 0.835 2.425 ;
        RECT 0.665 1.060 0.860 1.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.125 2.250 1.295 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.015 1.520 1.645 1.820 ;
        RECT 1.475 1.125 1.645 2.215 ;
        RECT 1.475 1.125 1.910 1.295 ;
        RECT 1.475 2.045 2.340 2.215 ;
  END 
END AOI21B2HDLXHT

MACRO AOI21B2HD1XHT
  CLASS  CORE ;
  FOREIGN AOI21B2HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.495 2.880 2.035 3.180 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.310 2.015 ;
        RECT 0.100 1.520 0.485 1.820 ;
    END
  END C
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.265 2.360 1.820 ;
        RECT 1.865 1.520 2.360 1.820 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.295 ;
        RECT 1.180 -0.300 1.480 0.705 ;
        RECT 2.050 -0.300 2.350 0.720 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.170 2.230 0.340 3.210 ;
        RECT 0.510 2.085 0.835 2.425 ;
        RECT 0.665 0.720 0.835 2.425 ;
        RECT 0.170 2.230 0.835 2.425 ;
        RECT 0.665 0.720 0.860 1.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.125 2.230 1.295 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.015 1.520 1.645 1.820 ;
        RECT 1.475 1.125 1.645 2.215 ;
        RECT 1.475 1.125 1.915 1.295 ;
        RECT 1.475 2.045 2.340 2.215 ;
  END 
END AOI21B2HD1XHT

MACRO AOI211HDMXHT
  CLASS  CORE ;
  FOREIGN AOI211HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.520 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.825 1.550 1.020 2.360 ;
        RECT 0.825 2.125 1.195 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.135 0.500 1.605 0.890 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.160 0.510 2.835 0.875 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.205 ;
        RECT 1.795 -0.300 1.965 1.295 ;
        RECT 1.560 1.125 1.965 1.295 ;
        RECT 3.170 -0.300 3.470 1.145 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.750 1.060 4.000 1.360 ;
        RECT 3.790 1.060 4.000 2.280 ;
        RECT 3.750 1.980 4.000 2.280 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.975 0.925 3.990 ;
        RECT 3.235 2.310 3.405 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 2.230 0.340 3.210 ;
        RECT 0.170 2.570 1.380 2.740 ;
        RECT 1.210 2.570 1.380 3.210 ;
        RECT 0.995 1.125 1.375 1.295 ;
        RECT 1.205 1.125 1.375 1.645 ;
        RECT 2.100 1.475 2.270 2.960 ;
        RECT 2.175 1.060 2.345 1.645 ;
        RECT 1.205 1.475 2.345 1.645 ;
        RECT 2.100 2.535 3.020 2.705 ;
        RECT 2.850 2.470 3.020 2.770 ;
        RECT 2.670 1.060 2.840 2.280 ;
        RECT 2.670 1.060 2.855 1.820 ;
        RECT 2.670 1.520 3.585 1.820 ;
  END 
END AOI211HDMXHT

MACRO BUFCLKHD10XHT
  CLASS  CORE ;
  FOREIGN BUFCLKHD10XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.510 1.520 1.100 2.020 ;
    END
  END A
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.695 -0.300 0.995 1.065 ;
        RECT 1.735 -0.300 2.035 1.065 ;
        RECT 2.780 -0.300 3.080 0.935 ;
        RECT 3.845 -0.300 4.485 0.935 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.255 1.980 2.555 2.895 ;
        RECT 2.260 0.785 2.560 1.385 ;
        RECT 3.295 1.980 3.595 2.895 ;
        RECT 3.300 0.785 3.600 1.385 ;
        RECT 2.255 1.980 4.635 2.355 ;
        RECT 2.260 1.115 5.005 1.385 ;
        RECT 4.390 1.115 4.635 2.895 ;
        RECT 4.335 1.980 4.635 2.895 ;
        RECT 4.390 1.115 5.005 2.225 ;
        RECT 4.705 0.785 5.005 2.225 ;
        RECT 2.255 1.980 5.005 2.225 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.695 2.635 0.995 3.990 ;
        RECT 1.735 2.195 2.035 3.990 ;
        RECT 2.775 2.535 3.075 3.990 ;
        RECT 3.815 2.535 4.115 3.990 ;
        RECT 4.855 2.405 5.155 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.160 1.060 0.330 3.130 ;
        RECT 0.160 1.060 0.410 1.360 ;
        RECT 0.160 2.215 0.475 3.130 ;
        RECT 0.160 2.215 1.450 2.420 ;
        RECT 1.280 1.060 1.450 2.960 ;
        RECT 1.280 1.585 4.115 1.755 ;
  END 
END BUFCLKHD10XHT

MACRO AOI33HDMXHT
  CLASS  CORE ;
  FOREIGN AOI33HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.285 1.330 0.785 1.755 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.805 0.605 1.130 0.775 ;
        RECT 0.920 0.605 1.130 1.195 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.305 1.265 1.540 1.820 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.125 2.480 3.590 3.000 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.395 0.510 2.840 0.880 ;
    END
  END E
  PIN F
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.540 1.950 2.015 ;
        RECT 1.740 1.540 2.070 1.840 ;
    END
  END F
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.145 ;
        RECT 3.225 -0.300 3.525 1.145 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.720 1.125 2.420 1.295 ;
        RECT 2.250 1.125 2.420 2.445 ;
        RECT 2.150 2.085 2.420 2.445 ;
        RECT 2.250 1.880 3.460 2.050 ;
        RECT 3.290 1.880 3.460 2.280 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.055 0.405 3.990 ;
        RECT 1.115 2.945 1.415 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 1.990 0.860 2.630 ;
        RECT 0.690 2.330 1.900 2.500 ;
        RECT 1.730 2.330 1.900 2.800 ;
        RECT 2.770 2.330 2.940 2.800 ;
        RECT 1.730 2.630 2.940 2.800 ;
  END 
END AOI33HDMXHT

MACRO AOI33HDLXHT
  CLASS  CORE ;
  FOREIGN AOI33HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.540 0.520 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.870 0.855 1.130 1.840 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 1.265 1.560 1.820 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.125 2.495 3.590 2.890 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.395 0.510 2.840 0.925 ;
    END
  END E
  PIN F
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.545 1.970 2.015 ;
        RECT 1.740 1.545 2.070 1.845 ;
    END
  END F
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.295 ;
        RECT 3.225 -0.300 3.525 1.295 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.745 1.060 1.915 1.360 ;
        RECT 1.745 1.170 2.420 1.360 ;
        RECT 2.250 1.170 2.420 2.445 ;
        RECT 2.150 2.085 2.420 2.445 ;
        RECT 2.250 1.730 3.460 1.900 ;
        RECT 3.290 1.730 3.460 2.300 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.195 0.405 3.990 ;
        RECT 1.115 2.745 1.415 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.625 2.195 1.965 2.365 ;
        RECT 1.795 2.195 1.965 2.805 ;
        RECT 2.770 2.130 2.940 2.805 ;
        RECT 1.795 2.635 2.940 2.805 ;
  END 
END AOI33HDLXHT

MACRO AOI33HD2XHT
  CLASS  CORE ;
  FOREIGN AOI33HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.740 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.540 0.520 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.870 1.260 1.130 1.820 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.125 0.510 1.645 0.875 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.055 2.560 3.675 2.940 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.065 0.755 2.590 1.130 ;
    END
  END E
  PIN F
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.675 2.830 2.315 3.180 ;
    END
  END F
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.295 ;
        RECT 3.070 -0.300 3.370 1.295 ;
        RECT 4.360 -0.300 4.530 1.120 ;
        RECT 5.400 -0.300 5.570 1.120 ;
        RECT 0.000 -0.300 5.740 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.880 1.175 5.220 1.360 ;
        RECT 4.605 2.045 5.050 2.425 ;
        RECT 4.880 0.720 5.050 1.360 ;
        RECT 4.880 2.045 5.050 2.960 ;
        RECT 5.050 1.175 5.220 2.215 ;
        RECT 4.605 2.045 5.220 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.195 0.405 3.990 ;
        RECT 1.060 2.745 1.360 3.990 ;
        RECT 4.295 2.635 4.595 3.990 ;
        RECT 5.400 2.230 5.570 3.990 ;
        RECT 0.000 3.390 5.740 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.625 2.195 1.975 2.365 ;
        RECT 1.805 2.195 1.975 2.650 ;
        RECT 2.675 2.195 2.845 2.650 ;
        RECT 1.805 2.480 2.845 2.650 ;
        RECT 2.675 2.195 3.015 2.365 ;
        RECT 1.530 1.060 1.700 1.710 ;
        RECT 2.260 1.540 2.430 2.300 ;
        RECT 1.530 1.540 3.825 1.710 ;
        RECT 3.300 1.540 3.470 2.300 ;
        RECT 3.300 1.540 3.825 1.840 ;
        RECT 3.745 1.125 4.180 1.295 ;
        RECT 4.010 1.125 4.180 2.215 ;
        RECT 3.745 2.045 4.180 2.215 ;
        RECT 4.010 1.540 4.870 1.840 ;
  END 
END AOI33HD2XHT

MACRO AOI33HD1XHT
  CLASS  CORE ;
  FOREIGN AOI33HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.265 0.520 1.820 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.810 1.520 1.130 2.015 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 0.860 1.560 1.200 ;
        RECT 1.390 0.860 1.560 1.820 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.110 1.265 3.590 1.820 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.500 0.510 2.835 0.720 ;
        RECT 2.600 0.510 2.835 1.820 ;
    END
  END E
  PIN F
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.520 2.070 2.015 ;
    END
  END F
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.085 ;
        RECT 3.225 -0.300 3.525 1.085 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.745 0.695 1.915 1.335 ;
        RECT 1.745 1.165 2.420 1.335 ;
        RECT 2.250 1.165 2.420 2.770 ;
        RECT 2.250 2.110 2.425 2.770 ;
        RECT 2.085 2.560 2.425 2.770 ;
        RECT 2.250 2.110 3.460 2.280 ;
        RECT 3.290 2.110 3.460 3.090 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 1.145 2.635 1.445 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 2.210 0.860 3.190 ;
        RECT 0.690 2.210 1.900 2.380 ;
        RECT 1.730 2.210 1.900 3.190 ;
        RECT 2.770 2.485 2.940 3.125 ;
        RECT 1.730 2.955 2.940 3.125 ;
  END 
END AOI33HD1XHT

MACRO AOI32HDLXHT
  CLASS  CORE ;
  FOREIGN AOI32HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.515 0.520 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.740 2.560 0.910 3.045 ;
        RECT 0.740 2.560 1.195 2.770 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.160 1.585 1.540 2.020 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.365 1.520 2.770 1.820 ;
        RECT 2.560 1.520 2.770 2.080 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.680 0.505 2.200 0.845 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.175 ;
        RECT 2.465 -0.300 2.765 1.295 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.495 1.125 2.185 1.295 ;
        RECT 2.015 1.125 2.185 2.420 ;
        RECT 2.015 2.090 2.360 2.420 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.895 0.405 3.990 ;
        RECT 1.090 2.950 1.390 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.535 2.200 1.820 2.370 ;
        RECT 1.650 2.200 1.820 3.100 ;
        RECT 1.650 2.930 2.765 3.100 ;
  END 
END AOI32HDLXHT

MACRO AOI32HD2XHT
  CLASS  CORE ;
  FOREIGN AOI32HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.920 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.430 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.840 1.265 1.130 1.820 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.125 0.510 1.645 0.860 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.960 0.510 2.425 0.940 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.550 2.810 2.020 3.180 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.175 ;
        RECT 2.605 -0.300 2.775 1.295 ;
        RECT 2.405 1.125 2.775 1.295 ;
        RECT 3.540 -0.300 3.710 1.120 ;
        RECT 4.580 -0.300 4.750 1.125 ;
        RECT 0.000 -0.300 4.920 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.995 1.130 4.400 1.295 ;
        RECT 3.790 2.050 4.230 2.425 ;
        RECT 4.060 2.050 4.230 2.965 ;
        RECT 4.230 0.720 4.295 2.220 ;
        RECT 3.995 0.720 4.295 1.295 ;
        RECT 4.230 1.130 4.400 2.220 ;
        RECT 3.790 2.050 4.400 2.220 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.895 0.405 3.990 ;
        RECT 0.965 2.895 1.265 3.990 ;
        RECT 3.475 2.975 3.775 3.990 ;
        RECT 4.580 2.230 4.750 3.990 ;
        RECT 0.000 3.390 4.920 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.535 2.195 1.815 2.365 ;
        RECT 1.645 2.195 1.815 2.630 ;
        RECT 1.645 2.460 2.700 2.630 ;
        RECT 2.530 2.460 2.700 3.130 ;
        RECT 1.510 1.060 1.680 1.840 ;
        RECT 2.100 1.670 2.270 2.280 ;
        RECT 2.825 1.540 2.995 1.840 ;
        RECT 1.510 1.670 2.995 1.840 ;
        RECT 2.990 1.060 3.345 1.360 ;
        RECT 3.175 1.060 3.345 2.215 ;
        RECT 2.975 2.045 3.345 2.215 ;
        RECT 3.175 1.520 4.035 1.820 ;
  END 
END AOI32HD2XHT

MACRO AOI32HD1XHT
  CLASS  CORE ;
  FOREIGN AOI32HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.265 0.550 1.820 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.775 1.465 1.130 2.015 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 0.860 1.550 1.195 ;
        RECT 1.380 0.860 1.550 1.820 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.735 1.265 3.180 1.820 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 1.585 1.950 2.015 ;
        RECT 1.740 1.585 2.205 1.755 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.135 -0.300 0.435 1.085 ;
        RECT 2.710 -0.300 3.010 0.985 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.745 0.720 1.945 1.405 ;
        RECT 1.745 1.235 2.555 1.405 ;
        RECT 2.385 1.235 2.555 2.755 ;
        RECT 2.150 2.035 2.555 2.755 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.135 2.295 0.435 3.990 ;
        RECT 1.175 2.635 1.475 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.720 2.210 0.890 3.190 ;
        RECT 0.720 2.210 1.930 2.380 ;
        RECT 1.760 2.210 1.930 3.190 ;
        RECT 2.800 2.145 2.970 3.125 ;
        RECT 1.760 2.955 2.970 3.125 ;
  END 
END AOI32HD1XHT

MACRO AOI31HDMXHT
  CLASS  CORE ;
  FOREIGN AOI31HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.590 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.895 1.235 1.205 1.820 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.555 1.570 1.950 2.015 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.585 2.415 2.060 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.210 -0.300 0.510 1.265 ;
        RECT 2.420 -0.300 2.720 0.925 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.895 0.720 2.065 1.360 ;
        RECT 1.895 1.190 2.770 1.360 ;
        RECT 2.595 1.190 2.770 2.940 ;
        RECT 2.485 2.300 2.770 2.940 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.210 2.365 0.510 3.990 ;
        RECT 1.310 2.705 1.610 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.815 2.245 0.985 2.885 ;
        RECT 0.815 2.245 2.115 2.415 ;
        RECT 1.945 2.245 2.115 2.885 ;
  END 
END AOI31HDMXHT

MACRO AOI31HDLXHT
  CLASS  CORE ;
  FOREIGN AOI31HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.310 2.015 ;
        RECT 0.100 1.520 0.530 1.820 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.775 1.225 1.130 1.755 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.950 0.505 1.670 0.720 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.615 2.895 2.175 3.180 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.045 ;
        RECT 2.020 -0.300 2.320 1.295 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.525 1.060 1.700 1.750 ;
        RECT 1.525 1.580 2.360 1.750 ;
        RECT 2.120 1.580 2.360 2.620 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 3.075 0.405 3.990 ;
        RECT 0.985 3.075 1.285 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.610 2.020 0.780 2.660 ;
        RECT 0.610 2.020 1.770 2.190 ;
        RECT 1.600 2.020 1.770 2.660 ;
  END 
END AOI31HDLXHT

MACRO AOI31HD2XHT
  CLASS  CORE ;
  FOREIGN AOI31HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.510 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.310 2.015 ;
        RECT 0.100 1.585 0.595 1.755 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 0.920 1.035 1.815 ;
        RECT 0.855 0.920 1.200 1.130 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.120 0.485 1.760 0.720 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.560 2.925 2.145 3.180 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.045 ;
        RECT 1.990 -0.300 2.290 1.295 ;
        RECT 3.130 -0.300 3.300 1.120 ;
        RECT 4.105 -0.300 4.405 1.055 ;
        RECT 0.000 -0.300 4.510 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.380 2.045 3.890 2.425 ;
        RECT 3.650 0.720 3.890 1.360 ;
        RECT 3.720 0.720 3.890 2.960 ;
        RECT 3.650 2.045 3.890 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 3.075 0.405 3.990 ;
        RECT 0.985 3.075 1.285 3.990 ;
        RECT 3.065 2.975 3.365 3.990 ;
        RECT 4.105 2.295 4.405 3.990 ;
        RECT 0.000 3.390 4.510 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.545 2.185 0.845 2.695 ;
        RECT 0.545 2.185 1.835 2.355 ;
        RECT 1.535 2.185 1.835 2.695 ;
        RECT 1.535 1.060 1.705 1.705 ;
        RECT 1.535 1.535 2.600 1.705 ;
        RECT 2.120 1.535 2.290 2.620 ;
        RECT 2.120 1.535 2.600 1.835 ;
        RECT 2.515 1.125 2.950 1.295 ;
        RECT 2.780 1.125 2.950 2.215 ;
        RECT 2.565 2.045 2.950 2.215 ;
        RECT 2.780 1.520 3.540 1.820 ;
  END 
END AOI31HD2XHT

MACRO AOI31HD1XHT
  CLASS  CORE ;
  FOREIGN AOI31HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.265 0.645 1.800 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.920 0.850 1.165 1.800 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.555 1.585 1.950 2.015 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.130 1.585 2.415 2.050 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.210 -0.300 0.510 1.055 ;
        RECT 2.420 -0.300 2.720 1.055 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.895 0.720 2.065 1.405 ;
        RECT 1.895 1.235 2.770 1.405 ;
        RECT 2.595 1.235 2.770 3.210 ;
        RECT 2.470 2.225 2.770 3.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.210 2.295 0.510 3.990 ;
        RECT 1.320 2.635 1.620 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.815 2.230 0.985 3.210 ;
        RECT 0.815 2.230 2.115 2.400 ;
        RECT 1.945 2.230 2.115 3.210 ;
  END 
END AOI31HD1XHT

MACRO AOI22HDUXHT
  CLASS  CORE ;
  FOREIGN AOI22HDUXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.540 0.620 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.755 0.510 1.450 0.825 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.105 2.815 1.730 3.180 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.130 1.435 2.360 2.070 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.275 ;
        RECT 2.055 -0.300 2.355 1.100 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.150 1.040 1.320 1.435 ;
        RECT 1.150 1.265 1.950 1.435 ;
        RECT 1.740 1.265 1.950 2.285 ;
        RECT 1.625 2.115 1.950 2.285 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.535 2.745 0.835 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.195 1.430 2.365 ;
        RECT 1.260 2.195 1.430 2.635 ;
        RECT 1.260 2.465 2.290 2.635 ;
        RECT 2.120 2.465 2.290 2.980 ;
  END 
END AOI22HDUXHT

MACRO AOI22HDMXHT
  CLASS  CORE ;
  FOREIGN AOI22HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.520 2.020 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.795 0.510 1.265 0.840 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.205 2.890 1.685 3.180 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.040 1.265 2.360 1.820 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.085 ;
        RECT 2.000 -0.300 2.300 1.085 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.025 1.065 1.325 1.235 ;
        RECT 1.155 1.065 1.325 1.540 ;
        RECT 1.155 1.370 1.860 1.540 ;
        RECT 1.675 1.370 1.860 2.360 ;
        RECT 1.675 2.150 2.035 2.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.575 2.945 0.875 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.235 1.405 2.405 ;
        RECT 1.235 2.235 1.405 2.710 ;
        RECT 1.235 2.540 2.290 2.710 ;
        RECT 2.120 2.540 2.290 3.180 ;
  END 
END AOI22HDMXHT

MACRO AOI22HDLXHT
  CLASS  CORE ;
  FOREIGN AOI22HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.540 0.550 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.795 0.510 1.225 0.875 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.205 2.745 1.605 3.180 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.130 1.435 2.360 2.040 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.295 ;
        RECT 2.000 -0.300 2.300 1.085 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.090 1.060 1.260 1.435 ;
        RECT 1.090 1.265 1.950 1.435 ;
        RECT 1.740 1.265 1.950 2.215 ;
        RECT 1.625 2.045 1.950 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.555 2.745 0.855 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.195 1.430 2.365 ;
        RECT 1.260 2.195 1.430 2.565 ;
        RECT 1.260 2.395 2.290 2.565 ;
        RECT 2.120 2.395 2.290 2.980 ;
  END 
END AOI22HDLXHT

MACRO AOI22HD2XHT
  CLASS  CORE ;
  FOREIGN AOI22HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.510 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.540 0.525 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.795 0.510 1.225 0.860 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.205 2.810 1.675 3.195 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.615 0.510 2.015 0.925 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.295 ;
        RECT 2.195 -0.300 2.400 1.295 ;
        RECT 2.005 1.125 2.400 1.295 ;
        RECT 3.130 -0.300 3.300 1.120 ;
        RECT 4.105 -0.300 4.405 1.055 ;
        RECT 0.000 -0.300 4.510 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.380 1.980 3.890 2.435 ;
        RECT 3.650 0.720 3.890 1.360 ;
        RECT 3.720 0.720 3.890 2.960 ;
        RECT 3.650 1.980 3.890 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.555 2.745 0.855 3.990 ;
        RECT 3.065 2.975 3.365 3.990 ;
        RECT 4.105 2.295 4.405 3.990 ;
        RECT 0.000 3.390 4.510 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.195 1.405 2.365 ;
        RECT 1.235 2.195 1.405 2.630 ;
        RECT 1.235 2.460 2.290 2.630 ;
        RECT 2.120 2.460 2.290 2.980 ;
        RECT 1.090 1.060 1.260 1.750 ;
        RECT 1.690 1.580 1.860 2.280 ;
        RECT 1.690 1.580 1.980 1.755 ;
        RECT 1.090 1.580 1.980 1.750 ;
        RECT 1.690 1.585 2.585 1.755 ;
        RECT 2.580 1.060 2.935 1.360 ;
        RECT 2.765 1.060 2.935 2.215 ;
        RECT 2.565 2.045 2.935 2.215 ;
        RECT 2.765 1.585 3.525 1.755 ;
  END 
END AOI22HD2XHT

MACRO AOI22HD1XHT
  CLASS  CORE ;
  FOREIGN AOI22HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.265 0.655 1.820 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.835 1.585 1.240 2.015 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.500 1.585 1.950 2.015 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.480 1.265 2.770 1.830 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.240 -0.300 0.540 1.055 ;
        RECT 2.300 -0.300 2.600 1.055 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 0.720 1.560 1.405 ;
        RECT 1.805 2.200 2.105 2.775 ;
        RECT 1.330 1.235 2.300 1.405 ;
        RECT 2.130 1.235 2.300 2.370 ;
        RECT 1.805 2.200 2.300 2.370 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.760 2.635 1.060 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.305 2.210 0.475 3.190 ;
        RECT 0.305 2.210 1.580 2.380 ;
        RECT 1.280 2.210 1.580 3.125 ;
        RECT 2.480 2.145 2.650 3.125 ;
        RECT 1.280 2.955 2.650 3.125 ;
  END 
END AOI22HD1XHT

MACRO AOI22B2HDMXHT
  CLASS  CORE ;
  FOREIGN AOI22B2HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.445 2.430 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.950 1.450 3.180 2.015 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.270 1.265 2.770 1.820 ;
    END
  END D
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.790 2.620 1.200 3.180 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.295 ;
        RECT 1.235 -0.300 1.535 1.295 ;
        RECT 2.870 -0.300 3.170 1.005 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.390 1.895 1.560 2.840 ;
        RECT 1.740 0.850 2.080 1.195 ;
        RECT 1.910 0.850 2.080 2.065 ;
        RECT 1.390 1.895 2.080 2.065 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.865 0.405 3.990 ;
        RECT 2.320 3.155 2.620 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.720 1.060 0.890 1.715 ;
        RECT 0.970 1.545 1.140 2.280 ;
        RECT 0.720 1.545 1.720 1.715 ;
        RECT 1.845 2.265 2.145 2.775 ;
        RECT 1.845 2.265 3.170 2.435 ;
        RECT 2.870 2.265 3.170 2.775 ;
  END 
END AOI22B2HDMXHT

MACRO AOI22B2HDLXHT
  CLASS  CORE ;
  FOREIGN AOI22B2HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.445 2.425 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.950 1.435 3.180 2.065 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.270 1.520 2.770 2.015 ;
    END
  END D
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.790 2.620 1.195 3.180 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.295 ;
        RECT 1.240 -0.300 1.540 1.295 ;
        RECT 2.870 -0.300 3.170 1.205 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.395 1.895 1.565 2.770 ;
        RECT 1.740 0.850 2.085 1.205 ;
        RECT 1.915 0.850 2.085 2.065 ;
        RECT 1.395 1.895 2.085 2.065 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.865 0.405 3.990 ;
        RECT 2.320 3.085 2.620 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.720 1.060 0.890 1.715 ;
        RECT 0.970 1.545 1.140 2.280 ;
        RECT 0.720 1.545 1.720 1.715 ;
        RECT 1.840 2.375 3.170 2.545 ;
  END 
END AOI22B2HDLXHT

MACRO AOI221HD2XHT
  CLASS  CORE ;
  FOREIGN AOI221HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.740 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.520 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.860 1.615 1.195 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.315 1.595 2.915 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.650 1.535 2.070 1.950 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.045 0.510 3.655 0.925 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.205 ;
        RECT 2.565 -0.300 2.865 0.945 ;
        RECT 4.290 -0.300 4.590 1.055 ;
        RECT 5.330 -0.300 5.630 1.055 ;
        RECT 0.000 -0.300 5.740 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.875 0.720 5.045 1.370 ;
        RECT 4.875 1.210 5.230 1.370 ;
        RECT 4.985 0.720 5.045 2.960 ;
        RECT 4.875 1.980 5.045 2.960 ;
        RECT 4.985 1.210 5.155 2.200 ;
        RECT 4.875 1.980 5.155 2.200 ;
        RECT 4.985 1.210 5.230 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 1.145 2.975 1.445 3.990 ;
        RECT 4.355 2.230 4.525 3.990 ;
        RECT 5.335 2.295 5.635 3.990 ;
        RECT 0.000 3.390 5.740 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 2.565 0.860 3.205 ;
        RECT 0.690 2.565 2.410 2.735 ;
        RECT 2.240 2.565 2.410 3.205 ;
        RECT 1.655 2.215 2.935 2.385 ;
        RECT 2.760 2.215 2.935 3.195 ;
        RECT 1.095 1.125 3.460 1.295 ;
        RECT 3.280 1.125 3.460 2.960 ;
        RECT 3.280 2.735 4.140 2.905 ;
        RECT 3.970 2.670 4.140 2.970 ;
        RECT 3.790 1.060 3.960 2.280 ;
        RECT 3.790 1.060 3.975 1.755 ;
        RECT 3.790 1.585 4.805 1.755 ;
  END 
END AOI221HD2XHT

MACRO AOI221HD1XHT
  CLASS  CORE ;
  FOREIGN AOI221HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.330 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.520 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 1.550 1.195 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.405 1.595 2.985 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.630 1.640 2.185 1.950 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 3.085 0.510 3.655 0.925 ;
    END
  END E
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.205 ;
        RECT 2.605 -0.300 2.905 0.945 ;
        RECT 4.370 -0.300 4.670 1.055 ;
        RECT 0.000 -0.300 5.330 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 4.955 0.720 5.230 1.360 ;
        RECT 5.050 0.720 5.230 2.960 ;
        RECT 4.955 1.980 5.230 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.295 0.405 3.990 ;
        RECT 1.145 2.975 1.445 3.990 ;
        RECT 4.435 2.230 4.605 3.990 ;
        RECT 0.000 3.390 5.330 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.690 2.565 0.860 3.205 ;
        RECT 0.690 2.565 2.460 2.735 ;
        RECT 2.290 2.565 2.460 3.205 ;
        RECT 1.705 2.215 2.980 2.385 ;
        RECT 2.810 2.215 2.980 3.195 ;
        RECT 1.135 1.125 3.500 1.295 ;
        RECT 3.330 1.125 3.500 2.960 ;
        RECT 3.330 2.535 4.205 2.705 ;
        RECT 4.035 2.470 4.205 2.770 ;
        RECT 3.840 1.060 4.010 2.280 ;
        RECT 3.840 1.060 4.025 1.755 ;
        RECT 3.840 1.585 4.850 1.755 ;
  END 
END AOI221HD1XHT

MACRO AOI21HDUXHT
  CLASS  CORE ;
  FOREIGN AOI21HDUXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.550 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.670 0.510 1.330 0.860 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.205 2.685 1.605 3.180 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.270 ;
        RECT 1.640 -0.300 1.940 1.295 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.125 1.060 1.295 1.750 ;
        RECT 1.125 1.580 1.950 1.750 ;
        RECT 1.710 1.580 1.950 2.460 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.575 2.880 0.875 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.195 1.425 2.365 ;
  END 
END AOI21HDUXHT

MACRO AOI21HDMXHT
  CLASS  CORE ;
  FOREIGN AOI21HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.265 0.550 1.820 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.795 1.625 1.295 1.950 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.240 2.970 1.840 3.180 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.005 ;
        RECT 1.580 -0.300 1.880 1.005 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.090 1.060 1.260 1.380 ;
        RECT 1.090 1.210 1.950 1.380 ;
        RECT 1.710 1.210 1.950 2.620 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.575 3.155 0.875 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 2.130 0.340 2.770 ;
        RECT 0.170 2.130 1.360 2.300 ;
        RECT 1.190 2.130 1.360 2.770 ;
  END 
END AOI21HDMXHT

MACRO AOI21HDLXHT
  CLASS  CORE ;
  FOREIGN AOI21HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.550 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.795 0.510 1.225 0.835 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.205 2.685 1.605 3.180 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.205 ;
        RECT 1.580 -0.300 1.880 1.295 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.090 1.060 1.260 1.750 ;
        RECT 1.090 1.580 1.950 1.750 ;
        RECT 1.710 1.580 1.950 2.430 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.575 2.880 0.875 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.195 1.425 2.365 ;
  END 
END AOI21HDLXHT

MACRO AOI21HD2XHT
  CLASS  CORE ;
  FOREIGN AOI21HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.550 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.795 0.510 1.225 0.835 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.205 2.685 1.605 3.180 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.205 ;
        RECT 1.580 -0.300 1.880 1.295 ;
        RECT 2.655 -0.300 2.955 1.055 ;
        RECT 3.695 -0.300 3.995 1.055 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.970 2.000 3.480 2.460 ;
        RECT 3.240 0.720 3.480 1.360 ;
        RECT 3.310 0.720 3.480 2.980 ;
        RECT 3.240 2.000 3.480 2.980 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.575 2.880 0.875 3.990 ;
        RECT 2.655 2.975 2.955 3.990 ;
        RECT 3.695 2.295 3.995 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 2.195 1.425 2.365 ;
        RECT 1.090 1.060 1.260 1.690 ;
        RECT 1.090 1.520 2.040 1.690 ;
        RECT 1.710 1.520 1.880 2.280 ;
        RECT 1.710 1.520 2.040 1.820 ;
        RECT 2.170 1.040 2.390 1.340 ;
        RECT 2.220 1.040 2.390 2.280 ;
        RECT 2.220 1.520 3.070 1.820 ;
  END 
END AOI21HD2XHT

MACRO AOI21HD1XHT
  CLASS  CORE ;
  FOREIGN AOI21HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.265 0.645 1.820 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.890 1.540 1.265 2.020 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.560 1.585 1.950 1.755 ;
        RECT 1.740 1.585 1.950 2.425 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.205 -0.300 0.505 1.055 ;
        RECT 1.920 -0.300 2.220 1.055 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.410 0.480 1.580 1.405 ;
        RECT 1.410 1.235 2.360 1.405 ;
        RECT 2.150 1.235 2.360 3.145 ;
        RECT 1.915 2.635 2.360 3.145 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.765 2.635 1.065 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.270 2.230 0.440 3.210 ;
        RECT 0.270 2.230 1.560 2.400 ;
        RECT 1.390 2.230 1.560 3.210 ;
  END 
END AOI21HD1XHT

MACRO AOI21B2HDMXHT
  CLASS  CORE ;
  FOREIGN AOI21B2HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.495 2.880 2.015 3.180 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.310 2.015 ;
        RECT 0.100 1.520 0.485 1.820 ;
    END
  END C
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.150 1.240 2.360 1.820 ;
        RECT 1.865 1.520 2.360 1.820 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.145 ;
        RECT 1.175 -0.300 1.475 0.745 ;
        RECT 2.055 -0.300 2.355 0.745 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.170 2.200 0.340 2.840 ;
        RECT 0.510 2.085 0.835 2.425 ;
        RECT 0.665 1.060 0.835 2.425 ;
        RECT 0.170 2.200 0.835 2.425 ;
        RECT 0.665 1.060 0.860 1.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.125 2.200 1.295 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 1.015 1.520 1.645 1.820 ;
        RECT 1.475 1.125 1.645 2.215 ;
        RECT 1.475 1.125 1.910 1.295 ;
        RECT 1.475 2.045 2.340 2.215 ;
  END 
END AOI21B2HDMXHT

MACRO AOI21B2HD2XHT
  CLASS  CORE ;
  FOREIGN AOI21B2HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN AN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.390 2.560 2.940 2.960 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 1.325 1.475 1.540 ;
    END
  END C
  PIN BN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.905 1.615 3.300 1.950 ;
    END
  END BN
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 0.760 ;
        RECT 1.145 -0.300 1.445 0.760 ;
        RECT 2.210 -0.300 2.510 1.080 ;
        RECT 3.250 -0.300 3.550 1.080 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 0.940 0.310 2.240 ;
        RECT 0.625 0.590 0.925 1.110 ;
        RECT 0.100 2.070 1.230 2.240 ;
        RECT 1.060 2.070 1.230 3.050 ;
        RECT 1.665 0.590 1.965 1.110 ;
        RECT 0.100 0.940 1.965 1.110 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.635 0.405 3.990 ;
        RECT 1.890 2.295 2.190 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.495 1.295 0.665 1.890 ;
        RECT 1.710 1.675 2.010 1.890 ;
        RECT 0.495 1.720 2.655 1.890 ;
        RECT 2.485 1.265 2.655 2.300 ;
        RECT 2.795 0.865 2.965 1.435 ;
        RECT 2.485 1.265 2.965 1.435 ;
        RECT 2.485 2.130 3.490 2.300 ;
  END 
END AOI21B2HD2XHT

MACRO AOI211HDLXHT
  CLASS  CORE ;
  FOREIGN AOI211HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.520 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.850 1.550 1.040 2.360 ;
        RECT 0.850 2.150 1.195 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.235 1.635 1.645 1.955 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.675 0.510 2.190 0.925 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.205 ;
        RECT 1.325 -0.300 1.495 0.760 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.995 1.125 2.360 1.295 ;
        RECT 2.100 1.125 2.360 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.975 0.925 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 2.230 0.340 3.210 ;
        RECT 0.170 2.570 1.380 2.740 ;
        RECT 1.210 2.570 1.380 3.210 ;
  END 
END AOI211HDLXHT

MACRO AOI211HD2XHT
  CLASS  CORE ;
  FOREIGN AOI211HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.510 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.520 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.870 1.550 1.040 2.360 ;
        RECT 0.870 2.150 1.605 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 0.510 1.400 0.890 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.930 0.500 2.425 0.875 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.205 ;
        RECT 1.580 -0.300 1.750 1.360 ;
        RECT 3.065 -0.300 3.365 1.155 ;
        RECT 4.105 -0.300 4.405 1.055 ;
        RECT 0.000 -0.300 4.510 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.650 0.720 3.820 2.960 ;
        RECT 3.650 1.265 4.000 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.975 0.925 3.990 ;
        RECT 3.065 2.975 3.365 3.990 ;
        RECT 4.105 2.295 4.405 3.990 ;
        RECT 0.000 3.390 4.510 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 2.230 0.340 3.210 ;
        RECT 0.170 2.570 1.380 2.740 ;
        RECT 1.210 2.570 1.380 3.210 ;
        RECT 0.995 1.125 1.400 1.295 ;
        RECT 1.230 1.125 1.400 1.710 ;
        RECT 1.230 1.540 2.430 1.710 ;
        RECT 2.100 1.060 2.270 2.960 ;
        RECT 2.100 1.520 2.430 1.820 ;
        RECT 2.610 1.060 2.780 2.280 ;
        RECT 2.610 1.520 3.470 1.820 ;
  END 
END AOI211HD2XHT

MACRO AOI211HD1XHT
  CLASS  CORE ;
  FOREIGN AOI211HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.100 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.520 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.830 1.550 1.000 2.360 ;
        RECT 0.830 2.150 1.195 2.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.135 0.510 1.605 0.925 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 2.160 0.510 2.840 0.875 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 -0.300 0.405 1.205 ;
        RECT 1.795 -0.300 1.965 1.295 ;
        RECT 1.545 1.125 1.965 1.295 ;
        RECT 3.170 -0.300 3.470 1.055 ;
        RECT 0.000 -0.300 4.100 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 3.755 0.720 4.000 1.360 ;
        RECT 3.790 0.720 4.000 2.960 ;
        RECT 3.755 1.980 4.000 2.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.625 2.975 0.925 3.990 ;
        RECT 3.235 2.230 3.405 3.990 ;
        RECT 0.000 3.390 4.100 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 2.200 0.340 3.180 ;
        RECT 0.170 2.560 1.380 2.730 ;
        RECT 1.210 2.560 1.380 3.200 ;
        RECT 0.995 1.125 1.360 1.295 ;
        RECT 1.190 1.125 1.360 1.830 ;
        RECT 2.100 1.660 2.270 2.960 ;
        RECT 2.175 1.060 2.345 1.830 ;
        RECT 1.190 1.660 2.345 1.830 ;
        RECT 2.100 2.535 3.020 2.705 ;
        RECT 2.850 2.470 3.020 2.770 ;
        RECT 2.670 1.060 2.840 2.280 ;
        RECT 2.670 1.060 2.855 1.755 ;
        RECT 2.670 1.585 3.610 1.755 ;
  END 
END AOI211HD1XHT

MACRO ANTFIXHDHT
  CLASS  CORE ;
  FOREIGN ANTFIXHDHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.230 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 -0.300 1.230 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.370 0.750 0.855 1.265 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 3.390 1.230 3.990 ;
    END
  END VDD
END ANTFIXHDHT

MACRO AND4HDMXHT
  CLASS  CORE ;
  FOREIGN AND4HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 2.395 2.190 2.865 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 0.660 1.650 1.225 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.445 0.510 0.785 0.895 ;
        RECT 0.445 0.725 1.135 0.895 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.540 0.540 2.015 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.305 -0.300 2.605 1.265 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.900 1.060 3.070 2.280 ;
        RECT 2.900 1.265 3.180 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.195 0.405 3.990 ;
        RECT 1.205 2.395 1.505 3.990 ;
        RECT 2.370 1.980 2.540 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.135 1.125 0.890 1.295 ;
        RECT 0.720 1.125 0.890 2.280 ;
        RECT 0.720 2.045 2.065 2.215 ;
        RECT 0.720 1.555 2.720 1.725 ;
        RECT 2.550 1.490 2.720 1.790 ;
  END 
END AND4HDMXHT

MACRO AND4HDLXHT
  CLASS  CORE ;
  FOREIGN AND4HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.740 2.405 2.170 2.850 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.330 0.660 1.650 1.210 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.445 0.510 1.135 0.720 ;
        RECT 0.835 0.510 1.135 0.895 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.540 0.490 2.015 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.305 -0.300 2.605 1.295 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.900 1.060 3.070 2.290 ;
        RECT 2.900 1.265 3.180 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.195 0.405 3.990 ;
        RECT 1.205 2.405 1.505 3.990 ;
        RECT 2.370 1.990 2.540 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 0.890 1.295 ;
        RECT 0.720 1.125 0.890 2.290 ;
        RECT 0.720 2.055 2.065 2.225 ;
        RECT 0.720 1.560 2.720 1.730 ;
        RECT 2.550 1.495 2.720 1.795 ;
  END 
END AND4HDLXHT

MACRO AND4HD2XHT
  CLASS  CORE ;
  FOREIGN AND4HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.675 1.585 2.110 1.950 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.265 2.795 1.750 3.180 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.830 1.330 1.195 1.755 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.310 2.015 ;
        RECT 0.100 1.585 0.610 1.800 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.180 -0.300 2.480 1.055 ;
        RECT 3.240 -0.300 3.540 1.055 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.775 0.720 2.945 2.960 ;
        RECT 2.775 1.330 3.245 1.540 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.130 2.425 0.430 3.990 ;
        RECT 0.915 2.910 1.085 3.990 ;
        RECT 2.180 2.635 2.480 3.990 ;
        RECT 3.240 2.295 3.540 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.130 0.785 0.430 1.295 ;
        RECT 0.130 0.935 1.575 1.105 ;
        RECT 1.405 0.935 1.575 1.405 ;
        RECT 1.405 1.235 2.595 1.405 ;
        RECT 0.650 2.130 2.575 2.300 ;
        RECT 2.425 1.235 2.595 2.295 ;
  END 
END AND4HD2XHT

MACRO AND4HD1XHT
  CLASS  CORE ;
  FOREIGN AND4HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.975 1.585 2.275 1.950 ;
        RECT 1.260 1.740 2.275 1.950 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.615 2.485 2.030 2.840 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.800 0.510 1.295 0.900 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.605 0.310 2.015 ;
        RECT 0.100 1.605 0.775 1.775 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.345 -0.300 2.645 1.055 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.940 0.720 3.110 2.960 ;
        RECT 2.940 1.265 3.180 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.265 2.195 0.565 3.990 ;
        RECT 1.265 2.640 1.435 3.990 ;
        RECT 2.345 2.635 2.645 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.295 1.125 0.595 1.405 ;
        RECT 0.295 1.235 2.760 1.405 ;
        RECT 0.815 2.135 2.695 2.305 ;
        RECT 2.590 1.235 2.760 2.295 ;
  END 
END AND4HD1XHT

MACRO AND3HDMXHT
  CLASS  CORE ;
  FOREIGN AND3HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.255 2.435 1.630 2.810 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.815 0.510 1.220 0.925 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.330 2.015 ;
        RECT 0.100 1.585 0.620 1.755 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.505 -0.300 1.805 0.745 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.055 1.125 2.360 1.295 ;
        RECT 2.150 1.125 2.360 2.215 ;
        RECT 2.055 2.045 2.360 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.645 2.595 0.945 3.990 ;
        RECT 1.810 2.860 1.980 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 2.205 0.340 2.830 ;
        RECT 0.690 2.045 0.860 2.375 ;
        RECT 0.170 2.205 0.860 2.375 ;
        RECT 0.140 1.125 1.500 1.295 ;
        RECT 0.690 2.045 1.500 2.215 ;
        RECT 1.330 1.120 1.500 2.215 ;
        RECT 1.330 1.520 1.970 1.820 ;
  END 
END AND3HDMXHT

MACRO AND3HDLXHT
  CLASS  CORE ;
  FOREIGN AND3HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.255 2.435 1.630 2.800 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.860 0.510 1.245 0.925 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.330 2.015 ;
        RECT 0.100 1.585 0.635 1.755 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.625 -0.300 1.925 0.745 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.055 1.125 2.360 1.295 ;
        RECT 2.150 1.125 2.360 2.215 ;
        RECT 2.055 2.045 2.360 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.645 2.595 0.945 3.990 ;
        RECT 1.810 2.650 1.980 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 2.195 0.340 2.830 ;
        RECT 0.635 2.045 0.805 2.365 ;
        RECT 0.170 2.195 0.805 2.365 ;
        RECT 0.155 1.125 1.500 1.295 ;
        RECT 0.635 2.045 1.500 2.215 ;
        RECT 1.330 1.120 1.500 2.215 ;
        RECT 1.330 1.520 1.970 1.820 ;
  END 
END AND3HDLXHT

MACRO AND3HD2XHT
  CLASS  CORE ;
  FOREIGN AND3HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.280 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.170 1.605 1.605 1.950 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.855 2.785 1.230 3.180 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.605 0.310 2.015 ;
        RECT 0.100 1.605 0.610 1.775 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.630 -0.300 1.930 1.055 ;
        RECT 2.720 -0.300 3.020 1.055 ;
        RECT 0.000 -0.300 3.280 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.265 0.720 2.435 2.960 ;
        RECT 2.265 1.330 2.835 1.540 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.505 2.900 0.675 3.990 ;
        RECT 1.660 2.635 1.960 3.990 ;
        RECT 2.720 2.295 3.020 3.990 ;
        RECT 0.000 3.390 3.280 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.130 0.785 0.430 1.405 ;
        RECT 0.130 1.235 2.080 1.405 ;
        RECT 1.910 1.235 2.080 2.365 ;
        RECT 0.130 2.195 2.080 2.365 ;
  END 
END AND3HD2XHT

MACRO AND3HD1XHT
  CLASS  CORE ;
  FOREIGN AND3HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.460 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 1.320 1.520 1.490 1.950 ;
        RECT 0.855 1.740 1.490 1.950 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.445 0.510 1.120 0.720 ;
        RECT 0.820 0.510 1.120 0.885 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.310 2.015 ;
        RECT 0.100 1.585 0.640 1.755 ;
    END
  END C
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.505 -0.300 1.805 0.705 ;
        RECT 0.000 -0.300 2.460 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 2.120 0.720 2.290 1.360 ;
        RECT 2.120 1.190 2.360 1.360 ;
        RECT 2.150 0.720 2.290 2.960 ;
        RECT 2.120 1.980 2.290 2.960 ;
        RECT 2.150 1.190 2.360 2.150 ;
        RECT 2.120 1.980 2.360 2.150 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.645 2.680 0.945 3.990 ;
        RECT 1.505 2.725 1.805 3.990 ;
        RECT 0.000 3.390 2.460 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.170 2.250 0.340 2.910 ;
        RECT 0.710 2.130 0.880 2.420 ;
        RECT 0.170 2.250 0.880 2.420 ;
        RECT 0.160 1.125 1.940 1.295 ;
        RECT 0.710 2.130 1.940 2.300 ;
        RECT 1.770 1.125 1.940 2.300 ;
        RECT 1.770 1.520 1.970 1.820 ;
  END 
END AND3HD1XHT

MACRO AND2HDUXHT
  CLASS  CORE ;
  FOREIGN AND2HDUXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.775 2.465 1.130 2.850 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.310 2.100 ;
        RECT 0.100 1.585 0.495 1.755 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.060 -0.300 1.360 1.295 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.640 1.120 1.950 1.295 ;
        RECT 1.740 1.120 1.950 2.215 ;
        RECT 1.605 2.045 1.950 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.535 0.405 3.990 ;
        RECT 1.325 2.575 1.625 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.105 1.125 0.865 1.295 ;
        RECT 0.695 1.125 0.865 2.215 ;
        RECT 0.565 2.045 0.865 2.215 ;
        RECT 0.695 1.520 1.550 1.820 ;
  END 
END AND2HDUXHT

MACRO AND2HDMXHT
  CLASS  CORE ;
  FOREIGN AND2HDMXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.765 2.490 1.130 2.870 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.310 2.020 ;
        RECT 0.100 1.520 0.540 1.820 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.115 -0.300 1.415 1.145 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.635 1.125 1.950 1.295 ;
        RECT 1.740 1.125 1.950 2.215 ;
        RECT 1.635 2.045 1.950 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.200 0.405 3.990 ;
        RECT 1.335 2.860 1.505 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.135 1.125 0.890 1.295 ;
        RECT 0.720 1.125 0.890 2.280 ;
        RECT 0.720 1.520 1.550 1.820 ;
  END 
END AND2HDMXHT

MACRO AND2HD2XSPGHT
  CLASS  CORE ;
  FOREIGN AND2HD2XSPGHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 2.785 0.425 3.365 3.360 ;
      LAYER V7 ;
        RECT 2.895 2.895 3.255 3.255 ;
      LAYER M7 ;
        RECT 1.590 2.885 3.345 3.265 ;
      LAYER V6 ;
        RECT 2.980 2.980 3.170 3.170 ;
      LAYER M4 ;
        RECT 1.745 2.425 1.945 3.285 ;
      LAYER V3 ;
        RECT 1.750 2.570 1.940 2.760 ;
      LAYER M3 ;
        RECT 1.180 2.565 2.055 2.765 ;
      LAYER V2 ;
        RECT 1.340 2.570 1.530 2.760 ;
      LAYER M2 ;
        RECT 1.335 2.480 1.535 3.285 ;
      LAYER V1 ;
        RECT 1.340 2.980 1.530 3.170 ;
      LAYER M1 ;
        RECT 1.195 2.765 1.630 3.180 ;
      LAYER M6 ;
        RECT 2.975 1.875 3.175 3.360 ;
      LAYER V5 ;
        RECT 2.980 2.980 3.170 3.170 ;
      LAYER M5 ;
        RECT 1.590 2.975 3.345 3.175 ;
      LAYER V4 ;
        RECT 1.750 2.980 1.940 3.170 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 0.325 0.425 0.905 3.285 ;
      LAYER V7 ;
        RECT 0.435 0.845 0.795 1.205 ;
      LAYER M7 ;
        RECT 0.155 0.835 0.885 1.215 ;
      LAYER V6 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M4 ;
        RECT 0.515 0.410 0.715 1.645 ;
      LAYER V3 ;
        RECT 0.520 1.340 0.710 1.530 ;
      LAYER M3 ;
        RECT 0.105 1.250 0.905 1.620 ;
      LAYER V2 ;
        RECT 0.110 1.340 0.300 1.530 ;
      LAYER M2 ;
        RECT 0.105 0.885 0.305 2.230 ;
      LAYER V1 ;
        RECT 0.110 1.750 0.300 1.940 ;
      LAYER M1 ;
        RECT 0.100 1.520 0.310 2.015 ;
        RECT 0.100 1.520 0.990 1.820 ;
      LAYER M6 ;
        RECT 0.515 0.425 0.715 1.730 ;
      LAYER V5 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M5 ;
        RECT 0.155 0.925 0.885 1.125 ;
      LAYER V4 ;
        RECT 0.520 0.930 0.710 1.120 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.745 -0.300 2.045 1.055 ;
        RECT 2.785 -0.300 3.085 1.055 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 1.555 0.425 2.135 3.310 ;
      LAYER V7 ;
        RECT 1.665 1.255 2.025 1.615 ;
      LAYER M7 ;
        RECT 1.440 1.245 2.405 1.625 ;
      LAYER V6 ;
        RECT 1.750 1.340 1.940 1.530 ;
      LAYER M4 ;
        RECT 1.745 0.810 1.945 1.640 ;
      LAYER V3 ;
        RECT 1.750 0.930 1.940 1.120 ;
      LAYER M3 ;
        RECT 1.535 0.925 2.840 1.125 ;
      LAYER V2 ;
        RECT 2.570 0.930 2.760 1.120 ;
      LAYER M2 ;
        RECT 2.565 0.800 2.765 1.710 ;
      LAYER V1 ;
        RECT 2.570 1.340 2.760 1.530 ;
      LAYER M1 ;
        RECT 2.330 0.720 2.500 2.960 ;
        RECT 2.330 1.330 2.840 1.540 ;
      LAYER M6 ;
        RECT 1.745 0.425 1.945 1.730 ;
      LAYER V5 ;
        RECT 1.750 1.340 1.940 1.530 ;
      LAYER M5 ;
        RECT 1.440 1.335 2.405 1.535 ;
      LAYER V4 ;
        RECT 1.750 1.340 1.940 1.530 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.630 2.395 0.930 3.990 ;
        RECT 1.810 2.230 1.980 3.990 ;
        RECT 2.785 2.295 3.085 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.630 1.125 1.450 1.295 ;
        RECT 1.280 1.125 1.450 2.555 ;
        RECT 1.150 1.980 1.450 2.555 ;
        RECT 1.280 1.585 2.110 1.755 ;
  END 
END AND2HD2XSPGHT

MACRO AND2HDLXHT
  CLASS  CORE ;
  FOREIGN AND2HDLXHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.685 2.460 1.130 2.835 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.540 2.015 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.115 -0.300 1.415 1.295 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.635 1.125 1.950 1.295 ;
        RECT 1.740 1.125 1.950 2.215 ;
        RECT 1.635 2.045 1.950 2.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.195 0.405 3.990 ;
        RECT 1.310 2.660 1.480 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.135 1.125 0.890 1.295 ;
        RECT 0.720 1.125 0.890 2.280 ;
        RECT 0.720 1.520 1.550 1.820 ;
  END 
END AND2HDLXHT

MACRO AND2HD1XSPGHT
  CLASS  CORE ;
  FOREIGN AND2HD1XSPGHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.690 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 2.785 0.425 3.365 3.165 ;
      LAYER V7 ;
        RECT 2.895 2.485 3.255 2.845 ;
      LAYER M7 ;
        RECT 1.995 2.475 3.355 2.855 ;
      LAYER V6 ;
        RECT 2.980 2.570 3.170 2.760 ;
      LAYER M4 ;
        RECT 2.155 2.050 2.355 3.110 ;
      LAYER V3 ;
        RECT 2.160 2.160 2.350 2.350 ;
      LAYER M3 ;
        RECT 1.640 2.155 2.485 2.355 ;
      LAYER V2 ;
        RECT 1.750 2.160 1.940 2.350 ;
      LAYER M2 ;
        RECT 1.745 2.025 1.945 2.975 ;
      LAYER V1 ;
        RECT 1.750 2.570 1.940 2.760 ;
      LAYER M1 ;
        RECT 1.625 2.510 2.245 2.770 ;
      LAYER M6 ;
        RECT 2.975 0.425 3.175 2.915 ;
      LAYER V5 ;
        RECT 2.980 2.570 3.170 2.760 ;
      LAYER M5 ;
        RECT 1.995 2.565 3.355 2.765 ;
      LAYER V4 ;
        RECT 2.160 2.570 2.350 2.760 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M8 ;
        RECT 0.325 0.425 0.905 3.085 ;
      LAYER V7 ;
        RECT 0.435 0.845 0.795 1.205 ;
      LAYER M7 ;
        RECT 0.205 0.835 1.025 1.215 ;
      LAYER V6 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M4 ;
        RECT 0.515 0.720 0.715 1.675 ;
      LAYER V3 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M3 ;
        RECT 0.105 0.855 0.820 1.195 ;
      LAYER V2 ;
        RECT 0.110 0.930 0.300 1.120 ;
      LAYER M2 ;
        RECT 0.105 0.815 0.305 2.050 ;
      LAYER V1 ;
        RECT 0.110 1.750 0.300 1.940 ;
      LAYER M1 ;
        RECT 0.100 1.585 0.310 2.015 ;
        RECT 0.100 1.585 1.365 1.755 ;
      LAYER M6 ;
        RECT 0.515 0.425 0.715 1.750 ;
      LAYER V5 ;
        RECT 0.520 0.930 0.710 1.120 ;
      LAYER M5 ;
        RECT 0.205 0.925 1.025 1.125 ;
      LAYER V4 ;
        RECT 0.520 0.930 0.710 1.120 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.900 -0.300 2.200 1.055 ;
        RECT 0.000 -0.300 3.690 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M8 ;
        RECT 1.555 0.425 2.135 3.130 ;
      LAYER V7 ;
        RECT 1.665 1.255 2.025 1.615 ;
      LAYER M7 ;
        RECT 1.335 1.245 2.125 1.625 ;
      LAYER V6 ;
        RECT 1.750 1.340 1.940 1.530 ;
      LAYER M4 ;
        RECT 1.335 0.785 1.535 1.715 ;
      LAYER V3 ;
        RECT 1.340 0.930 1.530 1.120 ;
      LAYER M3 ;
        RECT 1.195 0.925 2.835 1.125 ;
      LAYER V2 ;
        RECT 2.570 0.930 2.760 1.120 ;
      LAYER M2 ;
        RECT 2.565 0.825 2.765 1.675 ;
      LAYER V1 ;
        RECT 2.570 1.340 2.760 1.530 ;
      LAYER M1 ;
        RECT 2.485 1.140 2.770 1.360 ;
        RECT 2.560 0.720 2.655 2.960 ;
        RECT 2.485 0.720 2.655 1.360 ;
        RECT 2.560 1.140 2.665 2.960 ;
        RECT 2.495 1.980 2.665 2.960 ;
        RECT 2.560 1.140 2.770 2.195 ;
        RECT 2.495 1.980 2.770 2.195 ;
      LAYER M6 ;
        RECT 1.745 0.425 1.945 1.750 ;
      LAYER V5 ;
        RECT 1.750 1.340 1.940 1.530 ;
      LAYER M5 ;
        RECT 1.235 1.335 2.125 1.535 ;
      LAYER V4 ;
        RECT 1.340 1.340 1.530 1.530 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.900 2.175 1.200 3.990 ;
        RECT 1.890 2.975 2.190 3.990 ;
        RECT 0.000 3.390 3.690 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.940 1.125 1.715 1.295 ;
        RECT 1.545 1.125 1.715 2.285 ;
        RECT 1.450 2.115 1.750 2.285 ;
        RECT 1.545 1.520 2.345 1.820 ;
  END 
END AND2HD1XSPGHT

MACRO AND2HD2XHT
  CLASS  CORE ;
  FOREIGN AND2HD2XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.870 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.800 2.765 1.235 3.180 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.520 0.310 2.020 ;
        RECT 0.100 1.520 0.650 1.820 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.350 -0.300 1.650 1.055 ;
        RECT 2.390 -0.300 2.690 1.055 ;
        RECT 0.000 -0.300 2.870 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.935 0.720 2.105 2.960 ;
        RECT 1.935 1.330 2.425 1.540 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.235 2.395 0.535 3.990 ;
        RECT 1.415 2.230 1.585 3.990 ;
        RECT 2.390 2.295 2.690 3.990 ;
        RECT 0.000 3.390 2.870 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.235 1.125 1.055 1.295 ;
        RECT 0.885 1.125 1.055 2.555 ;
        RECT 0.755 1.980 1.055 2.555 ;
        RECT 0.885 1.520 1.755 1.820 ;
  END 
END AND2HD2XHT

MACRO AND2HD1XHT
  CLASS  CORE ;
  FOREIGN AND2HD1XHT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.050 BY 3.690 ;
  SYMMETRY X Y  ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.710 2.485 1.330 2.770 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.100 1.585 0.330 2.015 ;
        RECT 0.100 1.585 0.570 1.755 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.105 -0.300 1.405 1.055 ;
        RECT 0.000 -0.300 2.050 0.300 ;
    END
  END GND
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.690 1.140 1.950 1.360 ;
        RECT 1.740 0.720 1.860 2.960 ;
        RECT 1.690 0.720 1.860 1.360 ;
        RECT 1.740 1.140 1.870 2.960 ;
        RECT 1.700 1.980 1.870 2.960 ;
        RECT 1.740 1.140 1.950 2.195 ;
        RECT 1.700 1.980 1.950 2.195 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.105 2.195 0.405 3.990 ;
        RECT 1.095 2.975 1.395 3.990 ;
        RECT 0.000 3.390 2.050 3.990 ;
    END
  END VDD
  OBS 
      LAYER M1 ;
        RECT 0.145 1.125 0.920 1.295 ;
        RECT 0.750 1.125 0.920 2.215 ;
        RECT 0.750 1.520 0.955 2.215 ;
        RECT 0.655 2.045 0.955 2.215 ;
        RECT 0.750 1.520 1.550 1.820 ;
  END 
END AND2HD1XHT

END LIBRARY
